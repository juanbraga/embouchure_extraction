BZh91AY&SY�[,�p�_�`p���2� ����az�>                                    @P  
                       7` t (      _ 3XLCT6��04 ��4���>�S� �  �v- Ţt �  h� ���V`y��;�n�� &A#UӠ 7)�w+��         � �UN�Xj�Uu�R��S�� 1�i�Ӧ�r«�� �  ;�ã��N���RX�P��uu*ܹճnwR��swm
q:�C� 뺤��Rqwb9ې������         �)��S�aUw;�q��bga����u�v�W�K:1hV@ݤ��ʧ\M����3w0: n����;s�uJ�w
� �hunp�Jܰ*���[�5J�   t      P�&�
�T���,�]M\t -ƳN#�B�tv��åu9�D0 �q�B��u�n6;[M�	� u��c�d+��s #�ڱ��
s����Gu�M��ᠳF   h      �)��[����wAV1�.g@� 4��U��7t�]r�����  ��KN;vm�.�Uw7v�K���.�t����������sqT` t�B�q��T�n���]�ێg`�  ��ЛUJ�� 0   A�~6�*�4 h4 �H)�44Д�M�jz�'�4��L�B���T�'��4     ���HmUI@ ɠ   	SHeUM�42h�4�7{���p�����ٖ훴��4ٷ�T2�o�"4�"%�P��W2����,d�
��B��ۯ2���e�׌��Ɍ.�FV1�a��#+��tJP�
P�1!�UTU#M)Hb��@�M*PEC��UPIJ5�LCR�P���&�)����HP% ��1	d���!A��B�)CBbD�)*�����*�
F i"T���iJ�&*&(�ƒ!���%(ZhH����J:���)�9�*��"���b�)�S1B8��0�!��"���"��@��e*J�&�	h�h�(J�j�!� ��:���fD�"b�bk%	C����A�)�
F$��&!���Ab��D��*i���������Lb-�l�u�ء4%b�
"�	��)��m��]&*����( �: ��� �B�������4�	&���B��Z��p%"PM�@U	BhJM f�P�u@�@�!�ѡE�IZsUY	BP�T`�
jj&h����F�B�"E��*���(Ջ	̲D	�h���ӫ:)&���b�	"f�!���"�&B�(�	�	��0� ���*)Z���ht6�4L�c9U�(J�f��(J���*bh��������)J�(i�X���R�4ii�(i�&�ƍ���A������b(b4Ѩ�� ����F���"�(J����(q[	BPE@��RДM��SD�BPU%0E$�RIL�DP54�P��Q4�T�Q)T�%	BP�%���"�thJ�"Ji�	���f$)��K:�QZ���UTPU%ETБ!Eh��R%�$A1IgU:��`���	��-�TIEPUQLE2�EEMZ�E����lD�QADS5P�
hU4����������6���4j���"e�qI,�CV�
�)EV�D�3s,����%	Hmb��%h��	ѨH'a)�֓QPTV�Ƥ�+JhJa(��������M���P�BhM	BP��m��T�E-*4�T�f���(J��(J��J��	�4%	BP�$BP�%	BP�%�BP豄�ӡ(J��(J��ƗBP�%	BP�5��4�hJ��(J!(J5I�(KӶ�D��H�Ʋk�lv��ͤ�hJ4�!(J�Z�hJ��)2bt:�D��m��BP�:t8�h�Rb�hJL�9�BP�h�$�Chb�YMBP�Б4%q�m���ɬRZ��(�fƜK�@ca-��m�Λb�Y������6�M�Dk�4���h�i�V��T�1U[j���M b�HPD�ITE+�JPi4h)��Z�hh�$Ԓ�!�lTh��E1��Śt:4BP�	BP�%	BP�%	BD%!-0	BP�%	BP�%&�BD%	BP�%	BP�%,0P�%	BP�	BP�%	BP�%	BD%	BP�Q�hJ��(t�J3&��Ɉ1N�KjA�3��)44�8��+�t�J��(J!(J�� �!(J��(J��)	����
R��2L�TU"�*�-	E4�S.�MִL�	h�D�QD��LL�QC���A4SU@jj�#�A� �:J�.! �H4�����Q �
hM �QtĪ�+BP�%	�4%	&*0К��	BhM	BP�BP�&�J�К��.�"�l13U�"�M�%"P� P�a(J�4%	BP�&�J��(J��)��(`�P � �t*�eJAMascXӣ0XƔC�V�*�P���B1(h]+LH��MP4�J4�!%KF(H���i]���"��dȕ���
�H��Ε��6)�(H���:
J��)5��A�1����N���N��I&�֍6J1!E���*i(�j1�(J"(��:G@��-�a"$�(�f��j�t�J���
]!�.,I���*��b���f	J6X�D����l���6ME�P&�lجZ(���Eit��Z-�X�M	BhM	BP�&��%	BP�%�BV�"[	�(J�l�iqA�R�
�P��T�D��H���$�L��K�+T4&�mPV��F$�PИ�UTi���5�����I�EX�A�I�gBT��ZB����К��(H��)1��C1�X�D��c. ��ɤ0�t�:�	BP�%h�Y��N�1�"�Bm���Дit%	BD%�a�C�N�Y���bְ%[DF�LUCHM)��!�%@�H[)�P*�*����B
)(
()F� ��&Jb���L��uULALmh���؉b�)u�(��&�D�]j������i���Ц�������_o�>|?���_��_� EP8@ �u �  �P U @�@*� �  *� 
��@
�Umm� T�P   �� b� U��u �����A� J� E���ȶ@ )�  �� R� �P*� *�  � U��`*�(         �  � T�  �Rͬ��~߯�*��
ʪ m�M�  U*�@@*�  
��lk�!� � *T���@  *���U�@�궫o&�@�� m�U T �r� Q�U]����*��ۮޕ^�Z�^�*R�إ@^�@'ݫ{^��.ݡP��V�C�ln&0�mܸB�mQ8�]~�
�PG �U��zq�@< eQ��*�' c+:��m���Tz��AT*�f���Վ�w[���uS�M�mQs3��   N  8�e����-�����~�k��m����	��^�ꠜ*�� �z��ʣ6�U @    G�Tm�r��m� < < ���@T8��U�P�R���;���=UK���  ' c �T<��	�®ZUS�Q8�p[i��YE�w:Z�6ݍCp�o!�x����w�          Y@�
Ђr� �i6U�  N ����    
���     S`�K(U Y�   u��T�T ®�װ� U1�p��@^�	�:쇫(yTW��p(c��xn�Ͷ�ӄ�]��5Wv���<;�z��0۹��)ªx%e����^���d� ٵ�H�P��oVm�Gq�qp^̧;g�VW��8��.)f�7n�&K{M�w6ӭ� <��m��������{�����)�=����׫WD.܀�  x �0	�      P  � �;���605*�:N *��<�' c  <�� n N*��8@x wxc	�᳗�  N
��u�x�x�<C�p�1�p��e����[��͝Pp��}U�c �*�l��ft	�����[�U�m�7�UV5[�WV��y�� �8�YB�  ';l �p0w Np08u�z���K�Op��ڝh���Y��y����s9�ѵ*�  &�m�'�{�Cv��=����vdU�c��<   '[heS��B�m�slb�z� ��2 /  /T�]��� <�Tꡝ�;A�q���mˋm����0�xg�����[�ܮ�lw��Uՠ{lk��U�m�9iS��+\��Q���c5z/U�U�Ty�yӊ�O["uP�ˢx���wV-�?w��Wತ�l�P��'< ������xP����ꀿ���?���n��u�R�Z�8@U�+\���l���������3�כs[쪓�V쪧�� ' c�]����fܶޭC1U[���` 󝲛mݏV�Z�Ԫ�fz  Um��շz����mp����dL�V�ȷ��۶�y^���z۷��O\۹���s�Yz�m��U�\���Y;�\�y��ԫ��m�j�튽Uc�\��8�p�����g��+}�͹;�Yۛvm^��;�k�J< wy�R�-�Z��`����Du۽��s�^z�a��l��-�{�)��Mm�UJ{��Leʖ�����u�   �T  wQ� m�n��v�mG��t,���V4�7����kyiT
�*�P�������lۺvֶ�[��h  �yT�  5��VP �[*�3ɲ6ٽ�['�\\Umݢ���Ѳ ?�    *T񸊠PU*�e��*��Pm�<��
��ɹŐF�P��� �U
��  �UU�  ~?l�ޯʫb��6�m��;�ݩUk����` � ��@6����mf��ݚ��6���K��;�c�P�h�e�-#r-�P�Z�y�[]�Y�U����m�.g�{��@�
-����j<�  ��V�@{lNӱTVSmUug�@m�� �김��[b�v�Wum���UT����׳8�;���'yc���t��v�v����z���ٝnB�-�wuwUw m�k6��ض�͵EV�<VL�"}�N�M�J���mon�;�az���wr��e�{vWs{�]]y�*�7���]�U 
��
����={3�x;g�m�v��6ʠR�T��o]��t�9w.�[[�n[�<�l�m=[kݮ�j�  lW��M�j�����t��*�y�ռ��9-��X��V@	$p��*�eݱ�;������c:�۷{3|�,ܪ����[
����fez���u�w�ն���:��g�˷�^��;��U��x�v���y��0��ß�^����tg-��VMmk��{�F�    ��ޭ�   k� �� 
��  �T��� �*���N��ޓ��  ��   p�6�u     =l�  w �    ��5[O;�v;���wV�0�
�I��                                                            �           [��s����l TU       � � PxgsWu ;��    TY� S�w �Qs\�;�~�~ W�  � UY  �2� 
�        [V���߫�              
�                �  VP U         Y@        ;��          ����  z�A�66� ;��z��
� �     vh      뵰��@  *���֬c�T   *T P 
�V�*�6��^�獷��R��p��Ѷ�J��Wt�֠m�Kgt��u���                �          T                                    P     U ��<�m6�ث�    *��P  m�
�             w             �          �     *�                �-��               C�~   B���� ����V�� 75�;YT��wmh               �             �          �   m�       U   U  �YEZ`             *�     �       6� ��                    <                        ��� f�����	�X8@x x p  � ����      �                  < <   lP                                   �?              w            U         p p��@        ܪ         mT?7[*��         ;�<�  �   @�@  
�  
q U  �  P � ʡ���  \��        d 5Ҡ]�@   *T*�   �WsE̫�h�O��  6����{�zՂ�  m��fm��                 
� �P�     ���U6�����T � ��+�����)YJ���  �z�*�*�          ���wu��*��@    U U���;�P  P U @     �C��s�����κ9��p�ET@���D��y�׆�W�PP�z���\s�W����{�����S�T� l�
��TT��7ZTm�� �$    
��*U w�� V�����Ɲ]��{m˷"Uw⩮�� U�Z�ۼ��l���uDnu� �w R� c �]��h
�ᷯl첷t �p��AT U  � 0M���]�z�����eE�DY$���������N. �  v�-; ��'p�=���x7N������xU곶��dp����fn�綛������z�����+��@x��&�0ڜ�� �ujG��ݞ�/TT٦Z�����=�1�Sk�@x]@b�9Yt�-������4�����@�Z��PƑe2I�4��P����ۖ�0�P ��Sq�J��2���7=���mP³.��V��o\�����-��˦�m�wsO=��mfUy��e\��3�������s��]�f3Ԭc;��=��;�;wA[ק�=������dm[����J��4^��7nwn�kS��l��Pn�v�[ٽ�	�m����<�K�<kh��o_]�ݶ           �  \�@ U6�0 *��.`բ�  x      R�     UJ��m@�+%זV�T�ounӭ�ݞsc@            <T�[hUe  �    <    N   U �wUY�  
�      *��P     @   w    �-�N�
��      U      T  6� ` Un  �  w Y� `P�6���  <P�����T�   
�����[j�u=P \ͶS��  ͑o�����}~�� �����
��W�켕���*m��������k��N\������bt����{On�^OWm�]��O^��������*3�WSi��3��o{.�z=�ޭ��s}z�S�Wk���on� Wu��P*� m��n6�Ӹw�r�eUP�UVz��PGpEP�W���mUݖ��6�g6̽ﾫs]W�w��V��Zݽ �L�* 	��$U�u���m[{^����������'�b_�?�t���t�!�8f�)�=8F��NEO�,6�R[�)#n6Yqi�i���:�S�<!Qi�\#�)f��	�%ک���ydA���C$��yHf��QW�}�B�����W	���p�۔<��zk���317#@�Ɛ������
�8�������"Nue�S�t���ĄF@Kp�JE0S�S�����4�M�ɔ�N����N��&��L�Oz��[djF�Y �H��d��kn4�4��͝ѧ �P l��L�$�#�YRF�!f'�p���<�F��A�Z}��t�uU����5U	���p�8�2Q��4S��?S��4�wV��=0���N���o^R!�Sڒ�o��,�K�$�i��:p�]�pS�R�V�F���/d9O��
�X�)�\#{��镣V�ܘIΐ��ߕ?p�s��!���C���3�t�8�*�|s�L��v�\G��-�$&6E#�o�FzB��!�U!h<��4�+����)Ἱ�nI %�{{�=N�OkV{E�ٴ�s��{g�KgtU����@
�.�kkjUl�lnR<�B)ά��
a��w7�NEH�]T�H�v^DsH���5�|�H���܉�b����0M�R��CXG�R)��η>Di���:ꂜ:~������j�*�s:sŤp�:���#�����#?*t�u
bw��>��o�ԟo�"�$�-��2Cj���e�ϙg��
a��͎�ӑi"�U?R)�hb��hH�J7�H�i:x~TcE6�#�%,����{U"���Vgȍ3ο�l�]�w(<��n�]����	f5)`-�al�#`4�@J�ڭˑv�%�$�4LqAN~�j���H��t+��G�7��:zaz�����"�*%1��j8�`��p��q�j���e�ϙg��
a��͎�ӑi5���q�I�1�~�p��i:x~TcE6�#�%,����{U"���)at&�jFT���k>Di�]԰Y8i�Ecr�#�`�T&��,[x�R0��R�8	qD�rH܈RڸC�yf�?CzN:mXE<2�{3�F��mₘi���J�����ʻ{���/um�f:����ꝼ����@��ݫ[]�J|dmH[DƓs��H�����N켈�ç��F1�Sj�0M�R��F���"ܒH��v�ON����#L����`�?u�A�*�8q�
�t��<>��W-�d��,��#����#��B�<٧�ޓ��VO^����qi��$)���a8��~}خ9��+T��"��9!�#�OUCH�Մ,��p��RDdm�Ȋ����v��uR)鷙�3�F����; �?j5b�NU�s���?��J��m��ms���im�][�A�O*���R�r�E�v����A��xr�T퍴��׫�� �+�틺�g�nU�N�뷶��׆��f�BإbP�W,�T^^��'Jw�w�k�q���t�z  �`.`6� b�kwiWt6�m���R�B�UT    ��:�� ���AW�;6�ߴ �� ʹ
��~~���-�xn�O��*)�U��e�k�m����Tm�U[�V��H�@�-��CYf~�a�$ʫ�,��f���G�XB�s�N��6��ʌ"��&Ip�R#��9�㮮u�w&�+V�H�i��3H��·_V�N4�P�ᐤZ�;V���~��ڂ=��ONm�$��#L�}֝�S���5U-X$�(�6�1E����8q�UBi���ŷ�)���P��N��4����'���J�a-:pώw%�ϙa��L:~wb�4��:Ej�~�4����2E%��8�����:��5��ޯmziv�Vˊ��ڧp 
���JfV?�H�l
�m��x|xc��4�t� }�4��Ou�zt�<3�_%��ώ��8e���lp������=#g�T'O�G�o&R!���:B=8D��d-	$nI ��p�E�ӆ���>di�ۊ0��݊�ӇH�ְ�R���%H�j8�f~�0�j|�H�ӄ*�)���D���X=���4�ݹԜ*�fI$��y�#O8�t�b��U,piʴ�d�~�p�m�|�>=/�v�ij�F��L��ɽ�w���z��y�l״�hp@��U ��2RP��K-�0c�1;��hc�i��<����)��ן24�+o�O۷�`�HQC$�6�6��}����#����:��ߑ��|���G�Մ`�D���ޕxPe5!���6IfFڸE=9�w�gȍ<�}֝�S���T���*�8q�V0i����1�,!�,�ۓVs�p����όM��A��8~�����)��ן24�9=�^���llVň��ҝ?Ov+�NE�t�M?R)��C��:xB�aE6�"��썸ٍF��#��۶y�V����sU�vW1w�T� ���ڸ��$2�L�I����Y;�v�"��ڻ�3�F�q>�N�)�OڪX�ӕi#�a5�MĤh�N0i���ŷ��#��^��#��B�<٧�ޜtڸE<;x���$H�nRL���q[x��~{��ӑi4�O�ҷ��#��<0�jȂ*|�L�$�P�pڰ�h���I����"�����3�t���L�ç�R��8Z"\�m���ɔ��Ì걃O��m�yHç�qB4ú�GC٧Ћ���p�E6ܯ.��ޭ��fum��]]ݪ�uV��[[�mS� [7v���νmX� �?��S���>gL��AL4���\��i4�O�Ӯt2iP�%��IF$��#�OT,#M6�#�%,���������6��L�9�u#���RI��aBH�8i�UKӕi8Ϋ4�O��G��:zw#L;��7����%#��䍨�e��i��7NYj���/^|Ι�m⮮�W������d,$䅫^b�Fi��
��iڰ�r���C�mXE=;��$��U�j�+)��k]U���۞@�׊��#�w� ���iu�տ~� ���x;�>��y�y��{e]�[ӹ�k���Hy�����{U�uVfe�N՝*6��]�����x-�]s;���ե�Wgv�۬�3�P  ���*�� 6ª�:�9ʭ�6Ͱ6ʪ� k� P ;�U � �AUR��_�Y� �{mT��]r����W]����7�g{u{l���;���� ����B��Ͷ�V̷�\��m�BV[|�����q�F)�OڪX�ӕi8ɶi���y�ͥ��N(�NIr�o�˱��m�z�zg��
a��pP;�h���H^g�+�:t��yo��w\�<�_#xn��yy��;9�����i��$nI$��ڰ�zso_$ϑs��Kv1N~�R���H�ǩY��Gs[I:� �T��YH��)t��(F�����f�?CgS�ՄS�,�y�#Lⶶ�$m�v��6����촣mv�rk{�^(p.��M�U*�N�6պ�o[n�'#I$��
a��݊�ӑi4�K�y~�˾���y~�F�������w~s�φ$���Q�T��]'v��/y�Wy&|���.��d"�4���n2�#�ެ���3D��NCOԎ7r���:zF�cH�up��y�N��8�p�xs*�>0ڑ6�E�G|��8��PS?=�n9��M4�H�lG����Q-$�1��nA���0=�k:N�o���oI��]ү%�����R���ګ���w�w�o[{:�<ޚ��ܪ�+j���V�������j$�nB����Ƶ+�:�/my�_o�|���9����w'�#7��b�$\j%	.CH�:pݗ�>Y��di���v(:a#�N�?��IH"��m�!�G��ø���t>�<���
�U�W�{î��G��>H������z��v���(JK̚_ɟ���;���d�ld�.S�S���_ӡ(J<����&���/���N�~�w��iN��(JK�M/G�����	{a)�I�_ӡ<��w�).d���=B_,%v�>tm�s��\�4[��>I�_��(J��.��i����	}��y��&��;��]�!(J��&��s�'�����ģ�'ri|�	BQ��w�r_�i{�z��XJ>�i.�m��׆fS�������7�r���^��7�v��}��R��*-օe ;�j�%��{]��ss��ε��K��Jg�t����:�{����{��M/�З�ϛ�P���4���P�v�Ny�Ӱ>I�^�BP�%'Z��xu�i|�=B_,%@i?I���~~ۜ�����W9�s�m��9����)<�K��z���[��\��`4�$��:���y���I�����Q���<���v�_'BP����<�޺���~H��G޻���:��77:�:ۭ�h<��̏0=~/}�>@� ����3�%��Q���n����v|hJO$���z���߽�v%�i;�K��J�<����u�9s]r�9�r�݁�O$����^Y(���{�i|�	BP��I���|��c�����H���\R���M�uԝ�h��Ϟ���d�Δ���������m-�*ee����3ԥ���+�O��������d������;��G�}�W�G�c����m�G�������u�˜��9�^{��Mݽ�>n-۷�����ݹ������l�p 6�T�m6��m�v�n�W1�]u�uκ�_}��|���&��:n��\R�I�?~�R��)G_K�8�p�&��:R��(}�w��}�R��)G��h�����ϔ%���&���z���߻u�uínu��W]Z�s�jQ��ov�����������ԥ唣��ޓ@{:R�r�}�@y�f���ܥ픣��h��#�O�p�W�}���#�ϛ�\��W[�:뮎��p�_dy(��������>���̏���~y�{�+�0������{����Ҕ��{��w������/����13��vM�!��Ԗ��]�8v��Ҕ����=��]|�%픣䆇�4�ҝ�y��Hhz�@y�z���J:�_|�����JR��4>��{���s���t������ ��mUQA��N�����]�%)J9!��n��׾���w�4=ɠ=�)JQ��ox�p�&���z����y!��{�hgJR�{!��y�gκ�����כ}����� mR���N��M���n֛iT�%&�*�������y����P�76������C]]q���.�ݚ��w���c�G����`������ӯ`��UU�������$�f1�`����X  ���l� Vڪ�f{i��ʠm�U@ U    �
��� �*�T O�]��~�z� ȪVZꪺ��u^�V�oq�o7w�v�^ܷ��⫗�;� U�:V,�Ē�0Z�m1����	�s|�3�^(�S�ې�쇂j�/�ߧ���C��^��S�����Ý�H2ѐ��K`�<9!�>S���\9��z7M�l��J<HԵ,R�jD��l�=�
p�ry�*�2Fج��������כ��y�C��d�7�S������y������5�j��;y�d	)$Yd�9$O<4OT����|)���O7۞xj�@�J��܇7d<T�|��=�� �=�{<��[��e$��ae��x��wK��9!�:�����sTP����a��G�i��g66�hĉL��qb�92\-�B�.C��^�| w
��*-օP w]��Z����s�vÍG,3N���t�C�SÖ^����qZo$"�i��ՃND4�5��MDXm�F��v���4�t��B�4�mC�r���Y;�#�B��^sB�$�_G�6\nI�"4��d?S����\�CHӏR�O�ȝ)�&���a|ndj&�S��6�Swt�OUp;�d2&���(ďW���y�C��d�پ��qu@ٝ|CC	aabX-��������5@���9�D�:���s�N�h��x'�y����W����I-�d-�
�Id2ڸ��Ӷ�s����@m� �U*�*<�n�fE�4�KmɃNwd8&���խ�i"x�ڧ�*Xf�H�P�¥1qe��qG���=].��IQDZ��#A��;��)�2YH�[!��=�8u@
��r��잸�S���~��"�F����H���$Ƀ,������G�:'T�I��^]���B8��H�W�6Q��dda�����Yny�� =P���K�(������}�x�����;����(��vs����v��$�dad�.-À��w}�xh�S��i�T�O���w�H�N$}NOf�Ťp�w�m�Lժ^]n��{W.���j��l�;�]�ڧp 
�m���z�E��13��9�7�����G�:'T�H |�����4�:g�I����(�n	�H��!ɶ�(y|E���z��ďV��a�����W��d�ض[m�sM�)��y0�򇃹���xh�S����B�x'����<:�qކ?�V	⬵����I��۾���\�
���䍤I&z)vy,H�S] �.�����&�m�Y�O<4OT��<)�5~S�}�7ny� z�ǽR�J'�x�����<S�şN�d�I-�Y.F�xۻz��6��s���V�M���=�m�*�m��su����VҋS��p�O ��vs���tN���y0��.�w}�xh�S��i�}S�9�tb��V�-�J��P��9�����x��o�xS�}�sf�Á�8��}��8u|�D:'l�icG2KVF���T�{�O$��h�_Tھ4ꚻ�	7&�'J�$�E��H� ��Z}�m/ԫ+am�Œ���Ӟ>��!��?t5)�m#�VS�"LH�LM�d��D<�����`B�ke���]�D��>�O��ޞo9�!膉��y�O<���n�}i��8��vn�m��m�Km�I��P6�gszv����l����^��C�Ъ "�Z���y�������{~u6�.ܓ�w�߿L��Nz֥��{���q��M��.���^;�7k��oY�x��k��7����u
�v��.q�  ��7ҭ� l\�+&gnѶl�T�P�]@   �*��� T*�-��빰J�TEU��E�Z�[ov���s���o����ǝ߽۾��U�gP w�Wul�����x����F��M_9!�	�?�5@�5{u|����:��7
uM]�Y2mY"F�
¨��0�:i7UI]R��!s�����,�]�V���<]P;���G�HtC�O�������>��[m�ܘ����	��x޴��C�'��y�ë��7�yt�vC���y�Nd3μ��{������d�%���0�u(ǹe��qʄB\��SȄ#��p�u�
��G���[u�,�#o����*w���q�:'��>;�|�����>�S8'T�vs���u�:&�lvG��n��w�w_[��v6���ı�2ɐ��b�-�+Ui�������헂[e����j����w�<�\C���x��R'
��ҋ����xj\P8��<�svOCD�{�>?L�e��Il	l��*�G�ɺM��f��A��Yi�Dr��p7)�Bǧ9�M�1,��ж�h�e�|wl���w�o����;ى{�tOW�>{�|�����/��S��x��}w`Z�lR�I-�K<�4|�D>w�yp������d��D<���i�=쇢O�y>�W��_�p��$�m��Y���쇢'����<�
���n�}i��8��}��89!����TP����Y2H�,���N�v�K��Ύ��n�Pp���B� 6��2� ����d�a$��D=��q�T4wd<}�}�����W�fB��螯�w��xP���׹�
Ԭ��W
2�8'��t�9����^�ɇ5@�F���'�!��_���N�A�d=�;�}[)$�X�d%�7�%�l�'*�<p���Dq�^�W��?wZ�iȆ��Z�D1a�$-~�aZL�"��i��8�!dL��0Y�'��=�2=��[a�ȍ��q��rC��+J���U|܌t��t��?R8X��o#�t�^���E��b�{�]���ʽ[vuӳ�;�]��Cn�-��*�wEN[n�i�%k[l����s��}�|��<�}�aEN�/�#��T�Ȅq��V�E��jB�mDR�4�CH�-ս`�^�pњ�=̼�y�；�E��m�H�a�W�?r�݄F�n����Z$�%y��S���H'7ʠuC��y���ڬ�[cV���ǽi�~��I�|g�g�U)�a�N}�D0�����C��w�� HNF�$���DP>�w���!���k�T�t{p�^p�D�t�p�쇂w��4�E�,�䖡b8So]v��};ݲ�(�xU��ݳ� ��*ٵ�Y�Zdlmd�e��U��ݹNwd<��}�[�E��d���i��T�]��t|��	����X��HIa�P5CѺn�g�!���׽i�=쇢O��>�q@�o��Nn�x!�9���
U�!*�,%��� �=�zM��DP>�w���H|!��ArD�Ar�&��r~���&A�4�S�YL��]��7&�'�"��ǣ�O��m��<���U$<�d6Z�H��I!(F�r=�������y'/��-�Z����nG>��}�������_�W�UU �U�  �[&�ewB�T��@U�_� � �!T 
��m�� eP{��J�¨p���� ��uQ��-tU*����^���XL�s S`j�\ <� 
�� �U�����	�C��{�ewj{6  �U � UR�Q����ʣ�ٹ6���������{6���1�<�Sg�-u-n��@�  �����x N �0\8x<�W�V��k�WK����e� ����Now�sr��ޘ ��s���U�B���~���0U]96ރl.S�dk���ե�p����e`�����]ULj������s£�׎�w]UJ��{���Z�+Xm�;�շ�;�Mv���sP�{7my�%EPVU����������m���wP �P�U
��ثҨ ��w^�YJ�X���{v��m���[mfR�{J���^-�.��^��U�کt����Ᵹ��7k������ol�]�wj�6�Fڛ+����m�� �]�nm}�l�SSP�!��U�x��3r��:�`];��w�              �@ ��� Ux' @P �P     T  
�~�< T�U���`;�R�J� �owwm��Z���  <     �     �D�_��B�  �    x    U    ��U�J�D           0         �    �j��
�'      *� ��      P � t@ �  <   `e  ���U 
��P���s��b    ~ú��
���Q�-  �* ڠ���k{��� �R�m�-���gz�ka���]zU�{��U�ݮ�=y-�=�x���z�˾�^��u�����^�����m]pWVR�d�I,Z�ʭB�
�&,�Gk%�d���w^�^��ۥ]�ҠU  vʠ U  m�*Y�ۑ��n�V�UT*��   p  � � j���wT��m��ݭ��V�ږ�ꜵ�v��w:�ufζ�	ν�v�Gp����T {r�ۻw]�F �Q#$0d���?����#��T�S�Џu(��e��<Dk��+���$2&XrI#&��:~��Snڑ<Srk�~�,���1W"x���}ג`DwW:�*>�{$i6J��UT�2ӱЎ��1��'�<FP���S�z<���K����!����t�a�?[��ΒU��V(��S�MN�?B=ԣ喟��OLe,cl�e��6Y��3L�3��o�9��\�M�Ck�x���d�DYtb��t�O��Ѡ�I�ll"G[;:͚ڻ�����n۽d�� w�V�*���ibVB�&+e����_�;1;F#�T�=�8��.�qS"ydq�*���2�SuT
��+�-V��n�pա�a��U�#ܬ�nbv8�<t�K�âاUM��l���E��#��<E�NG�D8n�Sj�k�b쾎���*,(/B�-�#JF�I�<^!H�;x��DtZz/K��a��\�:,�S�M�l����&�)"K-�2yݻ��r��7[.d��_IՈqz9�p�;��o��Je�n3KI,B��Wo>�t˻��{�����*����;� *V�Vθd0��[l����V�:g��ڣ�B9�P��_(�(�!�M��}��9Ǥ����)A�h�ȲՒ!f!����#M����#��������qr���BTzmh���,����sJt�z��dC����E��B��Z��!���Sͼ�qΙ��s��4�I\��^��}iξ�ԧKRJ�%t���I1���d��`[m�\��������if��-�)x�#�6�rL�d_/�������8t�~�͒�)j"�
�k�v�U����y���ml�7YT�U�V@ �ܷw�����ۙTz�X��C�]�.x��c�O"�tݿK�c\kT銽vD6a��%��A��6�.�&��C��&ܫ����71;E�:er�tVj)\d�}�gf�e%�JX�,�w��rn;���.�ꛓ]�!f!�\�-G�q߼��C4�כ�Gp FI�Il��؄a��bS�]�e�.aX�$�!dC����E��Q�R�A�����ce�Y+��4��>K�)�B4��N"�|gjv%���J������l�m�FE-��!)[�P\TIC �F�#BKn]� x
�J�Wvکekd��2Im���+��n�܎�%�e�8c�H~2c��e��lF�KX�,����Hf��Ϸ_�\?Y�BĦ!��B�u�p��\��[���4��o$� J�,��K-�-��WC��!�����܋-F����dz,Ր�k��0�|�Q��15mD��7ٞ���y�z���Mh�5F���}���H���YE��m��M�ȲЄx�OV7p��|��/U\?Y��Lz,���.C?����{��O�����EP�U��{c��tڹ+B-zm�X�����Tsoi�ךl�����NcT�����k��ɽ�tն8@yj�;n�n�=-�u��ͣ�e�mw-�^���;�{wmwR����o]��y��ھl  6ͱn�� �m��m���tw�r�eUP � U C� � wU+mTS���n�< {7H[+2�S��{]���]^��{kv��6�⽮[m�����)�ڮ�,��s����W)g�dB9�:��F5ܙR��#���P!����0����=�5z_�*�Jӑ��h�����W1B)Ma�"j�S8E"��
���V�[��e��R4dm�����S�6_r��E#Ne^��QWu:=�8)D:/����P�E��)f6�,��X�� �%z�e�H뺌��%�3���fz?9EDB.%#���{s�㗋ޙ���܎զ�z�M�-��|��Q�����74ۻ{7v�gn��{�[��n��ݲ�����T \�U����km�0�"�����~>��}�;]��W�ӷ�����w�̒�u�h�ې�`o}���}ƫ�z��������Д�x�����J0 �$�U`�}ʈ�0˚����d7ڬB{�^���L�B�XgH��w���F��&I$e(L�:G�5B�y�3���VH�q�<Lus�#��3q߹�N�z�7���RH�d�I)a���|:��Yi��\�eX��<R)<,��l�R�k�Q�&6�.�j�>�j��׻��y�r�����7m̆���nX ��)Q�m��ڷ���n1����GB���L�#�^0�rήx��`��=�X���6�Ym�'�7@6�Rm]�<FZ�"}�B!�S*�k�m��VH�C�x91�7��s�|so�5)2�1[-��5t��O��E�&:,�-C�1��<C��II�BȄD��Y�m���m����9�j~^O{�G������~��#Mͮ0���d9ڝ�E����6��$���la9�לn�铦�G�|���O"�CP)�p��ܶ�w���f���wy�+mV�T���h�n�yƯw���wZ�7��6]m��[k� ��T�I�����,���g7��8����p�:,��g�>?Ytt��ӈB2�\(��Sj���*m��E^�,�G]��ƻ��TEOm��l�Ĺ���8�76��:+���VKc�Kd��D���3�xV����5�/�G�?.d��(D!��|����<{�|_����+@���B!�891��V���)��;�gЈs�������F�ȡ��&��t[4��!���Ⱦ�y�R�֝hzB}�!��7��}ftGe��$�cP�m�1��wW���g]Iw�S�+��,�ܩ�PguZR�+F6܍��Ǆ_,9��3��v�ON�>t1��=��܈"��0a1�!Q���ˁ��nGf.Z�����6��S"m��P�ۑ�X�nJ�7�u��*�u�n>�����=��Q>-4$i&܅Bd���!���9�sy����6t���]40M((�i8�I$
j�&�����K��P����b�So;�?����� � �UR�m��ŵ�7Yu6�ʺx�N=�
�m�.9OI�����ׯ ��;�a��w ��7�s���(j����[�W�S�-�7nӜ�T�]�wwW��V�Ψ���\h�ꪝ�s�  ;��R�� �6�[H�uN�`�UT�P��   �Rp � �*UR���l�����R�� v(7M����k�m�m�/vvN�OT��Wm̆��-�� m�إ_���6��&J�@�qA�-E]ܚ��]y�w�[ζ����Y�OdƉF7�G�ɞ�:�<�b�wwff��E/wu�fj:��Im�+�.uoGt��{��\�7��j�9nc�4[EA-F�e���;��������oVn��]�jN(ٍ9��U:�rH_���5���[�Ot��|�׽m[*�%��0�ik0`%��܄hAc%V��������v۷k��)B�14�����l��up�{�tl��ܼ�2Y���dIH��!i��q�ܰn�;���������VqӶ ȍ��R$�m�Y����ֵ�g���r���Z���:�$�ƛm�KE9�{�;4�Wz�Zw�'v-���YQl��	I���i%��w8�B��Z�մ��}�����Z~3���b��*Q��H[Tb�sV��w۽��;������\�T ]-�[v��q��m�YEǟi��|�����a���z�i.�0S�#��9ں~�~�<�H�(�I��b��Nԇ&����|l�1i�)��!�}>T�~�:�Ih"��4�uL�A7|Ck�Xf���C�»���XX ��  �s�ʰH�,��쿩�ϷX*���Ie�س.Ic�e�?4&Ax��ú$���[���WM5M�
~d_S�1�
&l�Q��9�]?p��;�1n�of|����꘴������]�o�$��m2D@��*Z5�*��ƶek'y������ ��J��[V����Ӝw��W�A�	w�6���3�~�8Wtu}��_�Tv	��ųŢ�)U�r5M����>�ڹ�O�i�y������O���F���ˈ��h��m���n�q����o|����C�w�bѼ޼����6՘��s�7󉯑q��Rf}�>'�}\��#h.�R-�ya�c���#�wGWܰ������T�t�E7a�ܳ���g�����Z~;��g�C��%<~�o�17��R�oj��w=���l�]�s��ݽ��ZQU��l+���Kl�ۄ�o���服6���]>%�y����e�����#�Sts{3�~�w�24�j3!�I$q����T��>iS��~�<�.��Zl̆��G��E��0�!�6�1��?p����"ՇD��g�Lo,>?R>]�i�z�J�IC$rI$`�3��B��F�xi�w�)���_��������ᱰ䑢���Mc�>g��<�~�0�H�OA�S�#Q���#1t����-�cm�����7V�{��)@�*�b����W)��Z���k�/U�����8tC���y[�z���w{���9+iW�9���
��,*¶H�����9T���^ٴ+w.���z��]�y��,��t�A窀 �j�lT TL���#��w-�m�@ �`   �  � �
���Pws�l��Tٶ��iN�ں���]OlZ[�{[��6�m�����n�'y���r旪n@3���)Z��HK}��g�<3�_���b�����Ȫ\,�q��f��u���޽g�R$�m�6�m��t���H4D"��K�[^:a2{�G��|sO�þ�b6���#h�p�Y|_D��Yk��U�6W-!�3�!Z�*�R=獷��)�c�r,��<ŹO=O&I����F�����:zE�g�cΘBPF�f(�mPk>����^�G��'@�ɑ�T�����j�ɺ�C:pͻͶF��ɋc K��z�޻WuK<��|�+���(�b����2~G�Z�m������<�~e���2��p�����ںC�Xg��=J
%N7�j����`���㑋�p�L�8׈ӛ�'̦�ۇ���L�r4�"Ή�'�ܸ��)��?A�~�f�;�w�{x��~R�I"��d��&O_����71�S|=�}qw����ˮ�TBc�1o�^3�x�zr�	��dU�a95؅�:G�ȫ�����O����Im�k ��b����]f��=N�F۸���6@
�UUV�֌�&����n&�NL���Z9c�g�c�m���J'���E�-�S*�)��<:�0�"RF��d"̊���{�b<p��nK�T#M����8�+�}�E�t��X�UF&�r�ǂ�����醑�p�g+�ZG7G��p�2*�0d�,B�OL����[L-��hY��q�=3��e_#�j���g�qc��6ӨR���0��5�"{1�jFꛪ�CL+�B��̵.fE^\K���8x��ܗ�P\9G�W�l	$�+����$�1��'j�]��t�e};�m�6k"��Z�w�wV�[o]�A��'D�*�v<p��eX��W ��äa]�r��@S���YH�j|m�Ȱh6ĶH�����=3�rc�ZM�"�/�#�����g��F��U�N�6�:�PD�i��@���g��V= O"5�.mw'��+��0��r��rv��w҅*��[I�t[-�8GE������2p�V:+��q����3z%�^��q$��7���BE���y=YMw�,äuɌUȞ 4߰���:-����,��2e6�l�E�um�-��l�וwY���-����v^T m��R�<���7�ym��6PLR��e��R����^��'���ڗ�����X���0�C�Ɂ��Z�,�Z�2��[��t���:,Ղd�V<p��eX��c�˼���=����T���ВK���f� !���1_v��Ր��B�:G�\��M߂�n#��){���6�j7P&&8tX*�ye��G�]_x��c�� !�O�e�-�����UE(�-���7j���0�Ь�����#��V	�UX��'	�c��N �[m��RP�;� T�3�����N�@�<m��ӎ�VQl[:��4���2����pz��ml����ׯ^U��o�wn���إy��<I�7)��;l��mt�8�tNl���r���W#h'Sj�s{j���  nY�*T*���Tm�;�;��� m�U@ �v�
��w   m� �*��EP�R���]X*s<��w"�޳M7}���k[p�$ D0,.Sr��Ned�ֺl�)[eYը�[�ԏ�c�7��<x|Gz��L��N1_v��Ր��B�:C�2��yN :v�N�ې���IN)3��g�p��g��c�喟 -�FS#:�m�@S�\��������Zje#"�MT�=�ϼx|p��+�w螬p����ľ�Q�oIIV�)�m��!M�wR.����ׄYt��51�����Y�&Mr�#ZSE�]6�-��%:lUȞ 4��R��dtY�\7��gØ�ǹe��c�]_x����=�ȶ[J��2�[dd����u��o9۽iU���k �ps��-�UI:e��m�{ᮻR�{��q7bz��,��n�b̇#����MV�l��d!eo3)��ʱ2 R�~8|E�侈l��=ǚD:{ŷ��%���p���N��på�o1�+����	ؒ�z5�+-�X�M"��F��5Q$�x��ݷ���s��G���{�<;��{�P
D�m$�%Ը�t�U�t�T����>�{��-KM��,PJ�ݭ���8��{^�6��n��%�����[����\Ү��כ�zU6S4)�W����r9��]TO�硨$��7sw�s\7�i���������:��Z;���"�ns�e��G^��+┦ɪm�]ؗ~�N��֜~��K�RNT.z������B��%L��A�S�I�&.o����qQ�F�y��^������Ɨ�0�"�������.�n�F��[�;��������|���6�D�Q�$��b(
���ae��U]k��EWq[��q� *l�w+l��06T���W�%�s������h3���@p�YO�Vqe<�S g�N,tNӈ�e�JA*m�i������&�{�t`���׼�+��vg�0�������N :v���|�q�aQ�ldk<~�]����t��`�m\�T#Uǚa�qA��4���$Q�r%$�4#ϲ-�:��=6��?�7�=@ap�>?{��9�S �O��m�D��5#16cp9���8�]K%����o��b.����k�OC�]�0�]D�Q��%&�c��1$/�(��ؤ��mu����䫼���' 7r�jl�v;݀-�j�����=)\?t[���	`Y���X6�E*���0�8�yQl�ς"�X��{�f�w�����7���o�p���.C{�s���^/\�$�Z�F�d�S�`�ι���u,��뵼fʽ�p��b�ܯ�7�]�4�K�%D��~��?WC-U����|eS��E�py�Xt��e�j�R�*�X�$�ZfD�D���0�8���Pxvn>GuoW�bM������r����}�6� 
�@`����
�6�� EQ�  �P,ڕ   �Q�P.JGϛ�m�l�����8o[F��)��m�y� ne*���Q9YUAV�-0��{b�8@xU
�-�;��v�c]@ U6 � P 
�ꁝPpz�;��76��6�vr��P|=ˮ��zV���j��   �k��h ��� ��78F;��g;`�*z�m����{����'S��ome�7n�g
��S�p]�y*��V��SU]m��狻l�T˚�NUw��q�=�P��`�p0!�ohPuJ��+��YG���;��n{���wU�ݳ�͛4���ە��O
�^�Z��s2�&�w�T�bۺ���[ eܹ�d`�Wl� x�l�.� ���ü]�m�=��s��]��Ͷ�ws��Vڱݱ[m��n����/�ۻ)��"��N�W���ڇw�]�x�B�[[kklkhU�:��N��
��vy�l��ŵ�ҷ��ުx&św���]�0{l�l�B�xس ,�%m}�             ��T  Ur��,�JUU@ `     T    �  
���mP  o �Հ�;�y��e=�O<@           �U�@    �        
l  PQ��3�:�    T J�        *�   p    8@��@      U          �  � �4 � 7 � lT@�N*T ^� =u�
�]�,2     NwS��l6��� ��l�  =r�k�� UG�N�m���[J���f]�n�գ�y�mY@\�y��I�w<{y�oS���wV��絝ה�ݶ�u=:x�,�oe�mfɳl�m*�����A+ek�%r.X�XYXQc�&����ݹ�  =�UOT�m�T�ig��p�w*�J�J��] ���J�� <�U*T�U۝
�ٮ�0���oq)2,UrH���IH� ����^�d�� wإG�W�n��N�I�i�?B�>2jv>8zt��R R�~8~ga�*� !��KV��A�i:��
j���-��-�C������f 4�)8~�"�w�,���9*��RIBI-l�i�Mw�4���_u��>�3�{�x��=���<4��/r`h��-RK%�8IN{�	�|~�+�c��U�ώ�2�kx�s���Ǉ�q�����j���,۽�p��b���y<]�n��~���U�'�7JN���dn���PU��}Yvzf'k�v]�z:���^�9l�6M�u���}vu��Z���a10t��e�j�R�1���ӊ�/5���k3�5ݝ�vP&���T�m��ws �)ǳ��ۄ잏�'��ӥ��RE����H�I:.���$���kD��@C���m{��d�B�?W	.����L���[i2�IeƳ����N�`�>6|:\��kN -�������t���á�/��������G>ƴ�-%����?�]Cp� ,�s����)��0zx}랍����)p� �8�k�W)�Jظr	���w�lM���< �X�WmV�ϳxpi������@r�r����h�i� 8�uñ_��KŴ�ݙ��>?}��"i�#n6�Q�N�_�ZCғ��E
�v%�Λ0s�c�f����~x���Q1(R��lP(��8k���X��ZK%�~3����@Yp����r�O݄��q��q$�I��qL�t��_sՅ�Ud���s���Qx�싥��Q�2TRF������_{��V��z����Av%�4���ǵ��wW��j2G$l�R�d�ov�����^��[ݮ�5�x�lJ�7;��Z۷l=�-�gˏ���}톯W��o�����դ��Xx�{�J��_�(��hPT[I$�.����.bw��:t��f����� U,���W��b�%	mI$�Fϱ��v�5�@��*����F:R`g��@�	�
\,��%$馝PAS����������C�&���o���*��/}�(/7#J9e�	�{��M�5e���W��$��v��
RǤx�׮�]U��T1�wZ��N4��ږ��������)�p.`���Sd���w3w����P'T�,�N���f�/�ƻ��4\�`QD�t�W�<_
��I�Fy{WL�I���R#�DL�R;Aw�jέ�3���H}PZK�_<ڝ#�Z�]��4� ٍ�������2;�(�rv�q�F�n)�&�"I.�o�b~@Z��F��B��b�N��"����ܾ̌!�z��Z�C"xwE}3w%/�E�Ȣ�&���6w3���޽+�^n�/%���-';���}����6�6�nU;�wN�XԶ��T��]X9�imT�^޺�]�c��{��8wm�l�G��|�y=U�o�G�J�x*�YF���#��{�@��U�y%�+v�^�Po+�fF�Bԡ�B�Y U�j�� �p����  �*�Z�s�ø�w R���P*�  w�@ m� ��m�* �-ޛm�[ym�ʠ2:���v=gq$B-���ȸ��Z���kl�k��B� ��P6R�G#JE�I	��������w���L�	���\����΁�T	�c16b�͓wW���:*�󷼞������wu��F����	Ѫm�J�U�O����S�Z��%�G}�0�
[��~C�љ|@V���Q_Q1�!�@�|��~�4ϣ��z��?Y��
Gr=r�7&�/��E_ˑIl4S�{�6�ws�E�[Tj����ra�ԕ��x�-*M� �&�v�ʟWc{=���n��WIT���]�UUP+H�r$�-�Ur�t�<;�WJ�EUG=삥�$��5���� �fF�,�������{����U{n?̞��^���g�ߛ?M(��Fd&Ofܔ�b�������n�6l���]�;�qPG����q(�fn��;���{��0�-zkkV�Ҩ�\�Nr�J�D��q��B�T�z,<F��p��^�
�!����G�SN��=�����{=#n2�T[-�u���m^��o:ީ�m�{{�w � �m�
�&����{�y�ݖ�%T�4�
��p�?��#�a�71���5�eX���"��~6|Eڽ�4��i�[m����~g�a�����_L'�i�������~~�74���w�Ɛ���Q���9���l���="�tO�\,��1�+�q�6���i��(6W�II$�E� �������^����"e�����9y0x�㦤�brg���D��4�	j�tj�Iߍ��R[/��!����MiC��H񆟝��S��ӳ���n��ʣ��խn��s�v�g;��w��[g��˚0 *��V�n��vp�&�Q�?Z�U� �����m\?B����~�PZԍ8u�hߑMI!nFۑ,�5�t�t{0�xi���L��H��L���VN^`���}<�AL2�r$���T?t��\�i��1{���>DS���cZF��<a��T;JVT��$��̜���=&�q�?n�fA�0���v�q��^�7��p�H)��#�@�G��i5vw�蹗�z�==����wc�rI!���;��m�l�g�e�ה�w_-�T�	��Pm�� 7-�[��}O-�1&�1˯x��e�^���$����<�E�4�Ϟ��@�m�H`HKt�:�}un�z��p��;���m�b�ζY
(�%$mARO7�Z%���<]S�SG�/(�
zyn�����2S2$J$�v�A./l�?{ٵ�վ\�����|�w����*���d����Z�C�OJ�_F����6���2����_���N*� ��G�)��G�܃�S�j�(w�ڨ�k�]=H�<̇��6'�z���(�{�����nuf�׷7s�U�μ��v�ޮ�u�H��wUs�ɰ����U�8�P�L�$a���F�"�s6���@ ��l6��
�;��6�m�u�m���U[ ��   p  )� �PT��@
�{l�ն��U����*yf3ڻݲj��%v4ݺ��e�إS�s�U6�M�uk[L�n�rͩJ������\����U������S�O�;��H�V�hI%��m�����i����r�`�!��/��T,����%����u�Т�I�]�����p�E�ϲ-,��a#�~z/�����t�p�?wW�G)�Kb��B5c�Y��X�,4C!ȕӆ�&;�Dx����Zh�yi��U#1���6��2O?x���,�#�9f���/"=2���K4�vw}�IKmŀۉr*�a���gS���m9��kg���]ڝ�PPW����4���6���?3���#��|y�#��_L$x�O�i�<��:u�/Ѱ��bjG.S�8V�81�Y�g|;X�g�d>��8a��H�i�ܲF��(�rHI9�:a��1���񐫧��,�&������,D:z|��H�J|Lp��EH�
Y�t�=���r+����3�M��0���[m�IY�ｻ�G��=A���t{�qY/���<��_I���Z��=k�o]�}��wkw�u�^]%��+�P�@�㛱��h�l�n%DEt�E<:(_q��w�Ӽ�E<4�}��4�4�+��~���|����m��FW����,{�4F�9�?]�&��Qp��w^~�~ ��4��ĶIQm�H��O�i�'��4���V9��=�¼�cH����Mcܰ����*� �F�uTH�]����<p��_q���kG�2���	�w'�~jG�-��R1p.��e���}�����I|o��r�Ӳ6܍8�m���9�
"܆8[,+)XAc*��R��*�w@Uw 
�&�Uݱm�����j�]�#kU��/e[O�un�z��p��;��o��4�0��2I 0'���K��/h����x��:�{�/.�_�6�m2Tn%NM[��O��z	qz�����Z��N{rON���M��ԍ(�H�s���T{�-^׾~>�]�ջ��{���Q��M�ڍĔ-����m��g����7�,�yը�o��۪�Y+���ň9 ������UqbT�e20�l�&]ڝ��T6��im#E��m��G�n�8HS�һ��g=v���^���{;���u���j �N8�qH�v7�5sӞ�z��m�����{�;]���m�n$���[��W����.wr=�{�g���Y���G~E���mH�V�����3F��~��(s��e������BT��nIm��ǽ�N�䞣W=9�^EE�׾�'���$I$�6ܒI$� �U�yC��Vf��v�Ү�*��� ]��׭��{��cx�k�y����ܪݸ��룺�W���wn��cz�;��w<�5���wC& �m�B̈�S1�I"�Ǎw]�y��v�@  ��U[ � �Sj�*�/���*��sT�T� \�� P 6�
�mT�*�R��|�Z��@VkԠ63�m�;�u�添|ƸWw�������T��( �P nwy���6�p��q����yF�o*�s���^m�aEȕӆ�-鴑*��Sm��Tt�E<;�cS�j�]m�������W*�#��虒���W���U/�N�#d����W��S���w�g�o�3�=���8r��H�8�]g���]��ŢG$)$��NL$x�O�E�7�T"��S<�?v����#�;E�W1B0����B&|�iH�PF�y����v�8D#OmƧ�j�
�R���㇏��U�&G��^�UT���Ooq'�۶���ݷ�]C[V�������U� *l��mm�ү���2$J$�2�����{�=/��k����ߡ���gd�t��Ă�A��t܅FQ�������E�n�n�/���0[��SSl*cLF��&ۊ܎�{�c�x����B4��[�}�V�~�f�xgO�����nKb�m�����L�#
`̗��r�+�&��x�~�,{����=����;�$Q��%:��!�n�#�\:+��꡾�ra#�~z/���B)pY�)��_z��=�II+de��$��t�;��뾽���L��m�V쭪w  �[m�ڎL�`�A�[tФP����A5�r�L�"�J������G��W���Zv��ፙ)$Y[+!y/)�����\w�FD̗��~WMV!���&+�x�E�Y��4�h%M��wFb��;�0�8W��mH��s�!g����b��2!|��C#��`��n6aq�,����;:�E�6w��=�120���0�/U���p�늙l2��Ȥ��3$����;��0Er�T��=�W�;��^����~0��j(Kp�v���Y{���޻���<���m��w� 7|Fjݷ7;��؋��}�r�p���gcG�E=v�L̹����H�6�&mM��m��ګ�2!6#��7�����qx���ژ�,���.�p��\�#^m����d��[�=2�����������1��8E����DȄxX�y��~y���"����m�Q6��"�"�%���24��p�Eڮ�;�0��UB�K�6�L�_F��������e�ҙ����%ș���#<����rqx����(G�}�6܍���c�����U=rn�+���e�r�%S�T�
����?�Ȗ�Y$��fy��|LI��8v�L�Fb�3d�;#��:B�;��7r�*�� �T��I�];F�^����b�"�%��x�D�j\"�|�J�>�=$��V
#6M��}ϼ�;|~���S��\�����PɑrPTn�d�)ƔrH7�f;{�L�׌ohY�.�)d���Ec��e#ӎ!_GJ����q� )ŗ�uӌ��`dmY�D5;�0����{��|���^˄C�ߵ��_��  *�� ����֮Os�@�T ��kU� �^L[j��m��Ǫ��jw�����筼�va��seS�i�)��n��ț���z�9��v�B���λ�m>�n���kuq]��^��@ ٶ�ɻ� �U*�m��;��p U*T �P  U m�j � �
����*T[���9� m���e�UW�q��˖�XEp�K%�z�ˋV]ږ� +n�Wc����l���p��?��#������.ԉ�ɓj��0����D�G��a���KP��*	����ꛤ��H;�0���Lz+��#(���C��{�y�Yt��k�D��}{}񙱩le�ڗ����4�D�+#��mF��{e�#y^�ɮ�B,�+�Z����<GS�Q!F�M�M&���A*w�]�c#�#㇨�6�ԋK�VH���s��UȸG��/���ae6rF��"�έb)b���Ǣ�\F�tNp|G8�ݡJD"���݅����'�$� ,l�[lT������5ސ��
��
� �n���^�z��E�黄+R-0�O���D�咮E�B4��,Q��HMv!�;�U]钓l��t�5c�^.#�J;����\9dw�8��0M�E�"Ò�U��S<3��|�5YR�$����όe�G�����Џ%�;Vqi#<��R'w9Tf$�)�#tPW�3����"�tZh�[2���dv�)*�-"��,Q�M�# (�%&�qFK90x���ذ]Y��<D��.�U�VJ�F�Q�m霮����l����l��e6^��졼��/;�7���R�ܪ��� *T�*�[`R���K�,��o�q�K�ֹ@��V�%I2t]z]�m��T~4�ۤ���
%P���Iy�Yt�2c�FR�?.%��#�dO�UȞ�����U�B��$ i�G�^�)�V!a�%��x�|����˄B.�p���G7�""���ɒ(2KF�%������}�#���UȞ!�Ί��土�3fo3L����s�Dac
���UՎ�18����|a�^���">̘��1�����=�S&r鎪��W{j��z���[ݺ�{�Z��Wwsխ���mS� �fһO�#s���l�i7]+$�`��]/n}����u��qx���\6a�>�B��-�L��@����ZD:n�U�.ԉ�ɓhX��t���Ur'��8�4G�س�)!R�)�T[t�A�A�#8xA51�f'���p��V;�O"�!��ɍ\#�?){���i2D�)mdr�<1�5�g;���i�]��g�{ 718�~s��M�I-�f�%e�e�8��]~��t����p���=Y2m����W5�:g�g��d�F��%��$%w,�ѝ�f��k�k�.��>਷Z� �	����{wŚJ�K���{�����|,m	p�0���c��N-#(��E��y�����i�K����%Sn�ԉ�WJU�����w�<P�6+�\,��<�Lċ�!�L���G$ʒ��j5��w_8�~3��K��#1Wq[*�-"7F	��jF��o�9�SOL��������H�M�\�ڄx�e�dz)��<øFp�51�f'���E��ړ��jܩd�U��n<�^��y���mH��r*{U�pÄ/�U�O��t�w��E����ﵥm�$�@  T
�6�0U ���P�  
�  P �P 
�U�wEQWOTm���nm��/*�:�� x�T���]��7�� ,Ȝ��UUGp 8�W� U��`��P�UO��[�7�Ӹ  *�P� �
�.���U��sǎ�»�A7U���v�m�n��������l6��  Ze� '<NyT�b�'��޺����n�����.�0ƀ���v wp�[.����2��U<  U��B�j�.�ݬ��2�p�ٸ�UOm;l����Q0��V�]�iX/l��[U=fP)�춼�=�m�ٍ�FԫL��,(u���7�۞{u3/rY��n�@�-��r[ʠ
�� ���;�[mn� \� �
�Fɶ�=l�U@ٷvMt���,�Yۻgf\�l[{F��n:+��͹*�կn�/t�mwk�����NX��׺�77��\���޴�=V]ʎ;'ok�ec[s�W�{m�Z��]��f�v������u y�b���ݹt��@             {-� B����nj�@*�*� U�  
�  
�� @� 
�ئʨ 
����E]� �Uۑ���j�;u�  �         x *���    `  �      6�   
�l�b�h        *�  *� 
� �    m�   �
����   8          l  �  w  \� �  ����*�� U�}�` l��T�����   C�n�@ *z� =�u )�  �٦����� ��WuR����櫸y�1�*��=fGp��G���j���o/<;���鷱9�v׭ժ�\�y�[�uj���6owg�_T��q\��Kmx;��ǚ�U��+`�,!SG!��5�ַ\��{T� {��K(  �sݶ�Wu�m���eUP���   �� ;� �*���S��o�۹�*����R���O)����{�o����\����o��w̀�*�m�w�k�[�wZ�a��e�UH�#�/îX���u���Uܖ�{����p���_[|��%����Y	e��Қz�\�����ӆ��[�=B��=�LtY�ŤzybF�Qt�uUI!@�E��y��\�up�jD���*�݈pÄ)�dw�=P�O6���KIV�bܬ�ҙ�|��s)�C��,tYi��:��pلf*�{c���L��--�d$�iUU4�"ڸEڑ=Y2m���K�W"v�9��=���OPW�w}�I$_!�ܠ��V���$q��r
##��B6�� �����۹���Y%�����x�}1��za�^��'�Y����W��OʺF}�9�xi᝝&��b�RK%[����z�lWl�YyM0��C���,tW���8S�p�f/u�H�k�l��m��uW�i�0MW�R'�&M�ba�C2�E��8#����{|渫Ib�%�IKr���=S]�]���K�����s}f��ݿ]ҮI��m��������-o�v0�����ZG�t��bjE�+�>F�H��-S%�[{����v[�[���]�wy�y����]��*-օP w{��:)�n���6���7pلY\�~��M�Sh\!��ɓhX��t���Uȳ#��_��I�$*��H�n"��3�w��ڱڑiD�aX�>�ȇ��(/��Z�B܍�J���|�T�U{n�8a�����j�i�]��dC�YO�є��}���Ӑ�$�SN�6ԋ�W2�\6aWP�r�C�A�m\!�ꛓX�0���2+-�!2��u��L��6�t�=��� ��=P)�c��N-#(��"�>�m�I�J�`�M��;���ol�u���y������u�ˢ�:@lJ@�r�"[l�%X��%ŋ����b�-}[|��=�þY������η�%؀JO�q$�-L�[����{��l�A�y��M��o&���Q&"�Ƒ)'[���nܖ
���y����N٪�q�sʝl�\pI20���͜��(|���c��_Vҽ�����>��{�7�*E!�"P.J����s
���ݘ��8���A�sw����(���d�$�\��I��Ny�׻�[�J�⮲��� ���κͻ}��G&6�BËd�e���Ǵ�Nל�i�w�C�:Û�=g�/"qղKam������!7/M:g=YM�c��}��s��#"�MO���`���j�o��b�m��6�}������.GE�Y	�)�3îX�^3_�`y��æy���mDIeI,� AUW�}P)�|C�ܫVL�V!f!�3\���M��'-�:� ���}#�d	�a��B�x=嘪/�*�񇈽V=2
���|y��WH�jz�����$�I$�6KrI -���mE�ۻE�\�����k�+^�[ � e3�_�>8A�'w����@VX4Rel�0�.KA���k͝�6�u��m��9��f�e�ym���V��w��9��u�pwc��ۛ   {l*��m�U� mLq�w�v�R�@ � @ �_���� �UP�[7�̀�Z���h�i��wN��m�m�ω��vۓ={ ;��x6G��m�XH��a�R�������?!_˟�|�W�`�ﲘE9�c����<:�.�r�u:U
a�n�T�i����a^dw�}�
|ʾ"�r�W2mX��:C�&UȪ��zn�E�#l��Xڤ#Ξ��_�ss��g��8p�V8ݪ��
�|a�,��g��U�:g��p�	�Fd�Bӑ�?Z���4��<pӄ-���u}�^�)���~úK�N����E�IIe������ǽ���K<��}Of�qe?Z�Ş��x�OH��6�P����'7�vow���]^��M���vj�*wAs� p*�m��m���Ά�{��I#A9�˘���=>?^.��ϰӇ�P��|�}����Ɵ���|)��m��$D�9�}N�Os��?Z����[�Cg���?yM_Y�;e�g�}:O�P��m�� S5Y�xu���j�S�S�O�G�?e���,>��~�_�e�v�-��¥��f���J=�e��/�e>OO��V�>�ϰӇX�_<�Ej�o���2
�6�`�3ǆ���O3�W��~��E���wS��}�8i����^������q��P���K2؟���,r���1.�wl��*�+m�� �ګ��[w��3�[<��a����|T�ƞQs��j�[�S�O�|Vy缾��������$䍶M�f��ܷƯV!g���L����2�'����ܵ�0��i����BK��A�Km�X�8�����%>4���3j�ҋ�/r,��V��>�=8c�u�0�2-�%��YϺ�����_G�|�O�x�:��\����Ξ3���EXL6в[m+�'����1�3�)mO�=����="p�*�+k�,t5�ض*��ꩤɧ#�K�0R�I �@�K����7����sB�
��.����6�:�iSuI���w��6}C��V:,���¨x��c�%ؾ�ƺ�Ư�ƻ��g^"M��T�@�V��8a�E��w}W���y�Dz-Ń�aO�"�{ǘ�LV/����Ed�DR�F[)	.<Fb�(�/��ѓ�"�w'�%ͫ���dʫ�/�߻chRuT)�#&,��/��<��&}��=t�|�tW����P>0���tګؾ��S	�a[Km�m�:g��[�N����^�%\嶾�bv˅�轫&xK�N�O��5-�E�ZH���2.2Id������.H�"�rwE��� �R����m�NmLZ8z?�_��1?��3����3H�Kؾ��&!|E��'�&M���(E� c(4�6�.4�.'��q}�)�t������\ÿ��8.�c��N/�*�񇈽R��d��I�ۀ���}��.rL�dV��_4��x���<��Z�W�9��g�"�oT��K�	�#mƙ,�ʿ���8u��qʆK㇈�U趥�@C�тb�"�w'���(�uL��4)S��a�C1U�O_C\a�y>���v!a����E�[�㽿�����QSb�;�T�t�n�ֹ�m/^���+m�`�c=s6��nc�����3kɷ�u�g�s	��d���;v\e�Ovoi��hwn{��;����ek{z�=o.�ar�c�ֻj�[6͵@ ���*8
� `lc[6[m���l�T�P \��  �l
� a�l p*��PT�ۺ� �Ng �ES�g���3�{]�;���]�;�y廔m��]�ڧp 	͵Vuؑ��ϴ��ֽ�g�������^�0�|_���ԋ֟JU�vfL��JΛґ�W�
*���F�����eN�kÜ��9��6G.���Y�f�V%>4�%�H�����ڎ����ʆ9��H������q�z-��,�b�>�C�Y��E�ꩺ4MՎ�18�����0��bI��b~�^=���-��})W����N�]#����m��w[���d�Y�Y��c��p֏_X�+�*B�vS#1>�lmē�H�F)�z������U웕�Շzt�w�VE[hU U��mݼ�T=�z�m�G{�i����ԉ�ɓj���#�d��D�~�F��7��ɘI
$��a$�$]4�~��P�L��1W!�e8���Wǲ{����쎮u�o���1�,�X�y�rp�\r;螡�u�.GE�X �)�"t�r�Ex�C�g;�P���%M��n���U�^�4�t�&��]�Փ&Ւ!f!�	��g��sI��Y%�ʲ�%m�4���|�	�b�B0Ç�@�Վ�18����|a�^�����a���m�hyڶ�7�w[�뙶V3{kb�յ��B��<� ��U����nܞ&4�m�@�wx�OʺR�m���^�%_D�C����p�:,��aLq�鳛��$
����Ɍ��������l�l�3x䗱i�7P,�:]��nп����e�-��m��n�.<�g?i����7�t^v���8}B6�-����?a�-i�n�J�YV��ۓ�����������5W��MvD8a��WO����iʛ/O�__��&�$���mȃG��xSӣ.AK�j��l�N��������	�Q�Y��&�I�i&�
��wu��Wf�:����=�����&�r������ fl�ٵ�j�y�gJƮd�w|~j��e�b��7�:~�*�O;�?a㇨@�؅�"GCgē�T˪�]��h{�
��a��3q���r�^�tfՑ~3���SP�4�u�fҋZKb[Yy��=�{��K��=4e�)ȭC�k��)��i��Y�zwo��2�U�Y,� �l���,�&M�$B�?W
��r�C���j��NUv�v	���O�y�O�1�R�UT��§bԈaN�����}�!�|�֯�{����L�dC���ͱ�dI
�)-�� R8Z[�k���'AuU�r�l@��-�vY��X�[+�$����3ӓ}�i�G��&�>���܆��cz�����"���[l���n�n�!�C��#5_�׹V).mY"a��H��O�t�����5m�Tz��.G%�t�#=P%6�j�"S����4=�_jG�u���*��1T��M��m�*ݫ"<~3���U�qn���������!㧅��[[9���$�[����"H9q�t罗��qu;T����Ҫ=�;zo�@���� �U�[�)�y���ץQp���m(*Yzۦw�Z��q�瓖�N�r�g�ۺ��KיS�� ��{�nΑ^��{Y���mhڽC�i��;��Z����Wz�����_w����t�UC  v�QT
� �k�Z�C��;���*�� �  @ �T �߿? �UP��*�Su��[]b�������v��*U�@�@�dL��-�� � ��T�Ul�I%1ƣiܒD?{�o��A77:�F�T���<焧��X��3���S���e���Hd��ZRE�a�>�����p���+�9V�#T�|~㶟�.R<i����+��e�$!��������e8~��9fU�4��Я^}���;�9�S��n���ꬴ�TlF��֑��\2���]��G�P�����Ȕ�|a���MI��$�6�t6/9Y|\�1��ϊžJ	�b<~3��~*׈�*l�?qg��)W�m���SS���;��z{K��緝ӣl�+���� M�պm�R�o;�*Fۍ��,�p���ːt��ap[�x~��9fU�4��Я^}�w=�&H�1��L$�<a��G��)�#�gY|~�Ǳ�~#�8p�cŕɑ#�M�BM��h�H�t�Ç�h{��^�"�9�/r,��5�w ��O����iX��6�{��A��i��)��]y��x��^�J:�#�r���NY�p�<9��0]ԅ%R4�
�_����ݑ���p�>*���9p�~Ӆtx�i:xV�5�M��孧���n��4�z�k���e��Uw��y[j ���nY���dӑ�R`�T#�xJ|~���9VN��/r,�������<Y���&�I�4�J9$�6T��b�0����~�A�.i:zT�A���]�ܧ�}/��5_'UTKI�4�"�8����>åEn_1��~t{�R��8}ˆS��/��)�&Z-�#���,�8|p��)�c���Ȕ�|a����VgO������ϧvi��Q$�X�^��r�P��gg���kAt����޳�<}�I>�fE$�����"V�+J�W���Kgt_T ;�lR�s�ګk�*Bԉ�ܑ���zٹ܈�o�{�k��jһ�U./���W�D�Q�ڐ݇�ۍw;�CQ��8UP�9�)��.��9V�g���n&�l�$�4�Y�<k�Z~�g�t�m��+�����0������sj���bnF�O�V�!鯦��6f���hW�>�J�ܾc>gO���2$�i$2I#P���֟�y��NA��f�ç��ݬ���6�CۗѶ�@�ځKu����{]�W�4̷<���޵gu����*��~�m���ܝ�v��s��x���ج�|_�/�j���o��m؇?P�٥b�0�?w�O�÷y2�*ےI(VR8t��.A���}6�8~�e\#O=
����Q?z���0!X�[%e��ҝ?N�u�F���3��?x�Z;��~#�P���Zg�8h̔��H�9���L�϶��mAg�b��U6�C���pW�ұis��?E�\�Ne?S��4�=>��i�j�>�f�!�DV^.��oq��ц6�nHL�H�u[�y���-�����P;�g�V�EՂ� �nK��n ��0{y�<wt@���̺�K��z����x䮼�����k꾅�h�n�Tn��m�ed�����2e)ʫ(e�.�����v�  �` U��l��"��Q����*�T*��  
� m�T< ���� 
�����R۽�[g�K&����uˋh� �0��X�,%`����w{f����Eꅲ 6��V�K\�[F�]�)���T���B�,��;�_׈�3��4��Os�F^2Y��4�A�n�	�aZ�r�H���g5at��G�{mO�˜�V0�QQ�E��J"��+������4�i3�?���h�VEq�~ 2��H��+h[m����|3�Ð��y��.�}*�,���P�)��gY`igx�p� L��.FIL9�#�H�(^�0�P�9D�WN��XF�2�w��������J���J�Y$�-*\��A�T�L�����k� ��*7yeUT����m��v����	9\�k�ੳ˸������h�VF�T�n$E��e����}��2�����h�ϡҚ�e���m�J�H�t��Y��rB�8�W|da߈��<�2ǋ+ɑ)�|@��wk�j�4����@RadeI(���|U��Sn�8@����V�E���;K6�<T�<t��/�i�r$��0iej��}�~�.�xGO3E�}�չ|�@�g�i&	� i����L���?R�Yr��
&�����u�� �SjH���E
��dml�Y3���3:�K9Z�s��|G�<&^|t�Z��8�m�:��$����u3���O�Ak٥W��C�	9\�Z�!���<��A�i8�1Em��1!YH����\�H:���m���L{;�<����?S"���"d�&5�m�bx��-#L���~����w�aӇ�8)�8�ʈ�.�6��4�6�Q�\���.�}��OL���&}�]�5]-�p��u�ZC*yI%bXŗ�ڣ�@�r��zۭ���׵�j��W��ȷZ@�ݪ������"R)ɔ�HT�������ua��:p���8�#�l梊L�ґ��a�T,8��Akt[��~��bR��4����8z�^A3H�����4�5Y
�$�m�t�֙��^��zm��U�S�{˼�>�J���߻�x��ͤ����#J9$5&iX��>{^S�0��S)t��.A���}٧�w�HD���=��q(\�yr���OK�7�W�kcK�e�}�3߭���+��$D	�ҥ�z�u]�gַ��;n�M��� wإWw�컵��%�$.#��Ӂw;΢t^w��Z�ݳ6o]��9Ӟ�|ׂ� di(�N7#h�y�4�}V{4�ZF�3�򟩅�e��D:z}� ��8E�ƙm�*1���i��i�)�4��:/V}�m��񆟯��äi�͂��K$-cll���O�8}��&i:p�wҿ)�k�v�{��8SI�"r%$�$Ò>���?s=�z����\�ֺK���_v)dm�$�I ��PlUeSb�m�wB������T n�  
��**UUTW�@U����ih ;��om�UP[� �S¨A+��T z㕽۳����
���TuQնӖ�n ��U�*��ogw� '�`��Ӻ�ss�   VZ` U +(
�����r��f�z���c�^�;v6�s�Coon{(�ZV��޷{�oL� �V� x< ��c ��[ʽz�v
�l�)UlT���d����׍�4����8�ݯWwR] �*��*���*C�����{��z��k��
<�x��4���M�=��Հ��j�T�β�V�Wu���RHJ�)%���%Ƶ)W\�wc�������w{?~�����ܪ�@�����{��ܺ�t/l�Ps�n� J��~o߿eJ�EUU66l�:�AYn�=�l�rv���YB�wS���wz�m)q����6���mz��1�]Ez�v��n��]��s�6.e޾�ݙ�yV�;����w���N�+��7۳o��`]p]�w*T�7uhb�ջW;j��             �Ѷ   ]��@m�w] *�      ��      �  `u� 6�`ī� .:��m�S|a�A     @      ~x~ Ͳ@   w  P  *�  m�    U/ww8�           �+(   *�     w    �
���     �~           m� ;� �   <  S�T�   U�Jl *�-� n�n�uX   �l��� �J��y� ��� T@ w*�����~�_��U*T�TU����6���]�y�@�捰 ۭ݃��-��)�m;.�y�wp�uj�;��5P
������l��r�'q���=��K�T+ּ 5�#��'�b�
4���+�����  v�U[*��
�lBv�����l�T�T�   lST� �j���
���ՠγ�ڕ�-���r�@�`�!DJ��/���T�;��ۅwV� 
�mU�Ժ{���Ӥ7$�+4A�7��c�ǣx�^�{Z�査��Sp$�RC$��K:~��)��5�xsO�a�*>�:a�>?Cw��F�K�m�Fᕗ9ҟ�&��3�{�T˱?N�r�l��2�)�2���n,�e%h�$�N<�C���r
YӄN�lӇ�>�9e8F�=gE�ϡ�
��|�!�$n6���2,8i��y�K:F�e8�?i­���C>6P��m�YGI�Q*�T�j�.����ܲ8���j���+yU@�<T� \�Wns�g�;l�ܽ�?3^=�آ<p��1��ψ��T��ǇO�x�H�!~��?9j%#�")ǚ~�K�28w�`҈d>�?C�Xdp����DL�J6ɢP���~���V!?yIA��a�|~�]O0p�C/��^2�HF#m�h�)؄GH(C���_ȏ�)rg���w��i�|�h��1��R����;��R_��!����龂�!�݂��﬌��&�0�Y�ҥ�C�(#c��oYwP]� 0[���V��o+l�@̂��#�j>��?-��!:G�4��<����:F��-��M��m�-�v4�Ep���\$v	:��H�o^�$(D�-�6�hj��#��%��3�`]/��+�.�<E���b�A�䪚��5M*��v�,�W�Fh��+�~Z;��<F������=���#�#��aߍ���*X�}Â�V>Dp��<?Qm���=�������a$�Y��{���n����ֽ�-Z's��m�wM���kkl�׹��u�N®�?��{�
q�#M����B>��{�M���x�FN	a0F�%M��n��D�g0���20�-G�_�B�t��t(l*5�����>�_c�꣗c�&�qN��.�����[rI"8��ڽ$ݾ�O2f��N�����~��ƀT9E���2Y1�W�z_��m}��i�[�f���I�$,F�PZ��	/ꔑ,Y0�m{�s��x.h`�r ��w7u��ۨ��( ������ ���t��s�釯W�pi�{I��
p�{���*�Jq��RtAlX��0�p_��*E-����{���=p��훹��lH�p��%��r�ءr�_y[�A������v�'i�[m�B�E�5��}��n�
�����W�v�[�~H�"I5m��A5绔zxn�}q��_��&���������i&�IF�2-��T����2�Ǫ8�p8G�Q� ����u������ǃ�ά�wI˛o�����y�lZ`[Ν����r7ӞĜ^n��n�n�[�ע����wu���u��ٶ   6u���
� ����J�p`m��UT*�Հ   p@ � �W��?U@�*m�w:Ǫ��l*��.�j�n��s{��{^+mR�T��V���;�,� ��J��]jۻm}vw�iG$�Ƥ�-�������rl�wֻy���r�Ї�)2��i8�J罗7��v�d�w�vr����kT=���E����� i��t��6��@��1}x�"����s)⧦���9���i�$mLO2a��"w,���F
mX�;���b� ���Z��:D��Lߙ��ܑ�[�H�OA�)F�;b��D��8� �GFވG��q�]mUQ�m�U1ssf���ٮ[�wZ﷍�nu;�����6@
�Vګb�z�����w��#�"�¶T��R0ӇY4p�ܰ�C��#�X�6�ȇOt��!k!m��,��L�=7���]p�ܲ;�qeڸY,9���s:e:zw��!��TiY-�v$VaE�96x��Zs�,�6|�yH�T���0�����j6R�$����"��6�R�"�ҶT��R0ӇX�qAj�H�=�R�9�]�ԟ%Ŷ�-���[�2���&:�"��t�^�dC�!w,���FF6�D�\�JSt]�-�ʱ�$0�a+e,2�x�]�T�*٬�«]@[�k�[��w�vP�%N��!�:e�bD�#����g���<���S�E��)�O
��KZ�#%e��d�嗔�)��ok�t�)�S�S�Z�Vʟ^
Fp�&�4��0��t�
5
Jc)f�����:_����x�)V�)ᧄ+Wӄie��!4�7n�m�:�,�6X�&X�(��/�,��,���t��#�t�*DlD�q(�l���D4�]��G����G�m��b��<ڟ-�[�$��#A����շu��s{��z�l�=��۶����� )Q���m�i]�˷��T�K� {F��6�=��i���߻�緝�ף�����-�Y,�<���]v1|n/Y{�}U����zYY@�QQ*�L6�m��/�(��W:�H�g���Z���i����8u��I���q��r4Ӆǂ���;D��Ǎ�d1[��h��,zvU��:}p�j��<p��p�2[uM���s&O<!Z��#H�Y�^��N(���R!���},�0�����m��l\�{zmw����fz�e>;��ut��w��[`�Cm�ٵ���u��!j)�6X*s���0�NzR!p����D4�_�	�OH����8E#�ݾ.�[jL��T�4�<�}��Gw���U��������~��W����쫑"V2DN�e�ۥT�6�5{��<�p�d)�)��C��(����dCe��*��"�>�%��&�:J�l�U�h�C\G�"·�mC�SÌ�Ք�i�_<$x�OL�ξ�F��Ʉcy�3�zM�ӄi�]ڟf
Fp�&�4��0�.�)f���(<�6ܒ6ˑ���N�S�uJ-˹�3�ǀw�T��ZEP<��w�Z�*><�A�]�=����^*��m���r���S׺�{�O\+ks����M����V�W��*��/w*���ַ��'^�  m��*�T l�ĥ^\�p`w7�m��P@ � �  �� �T�ߏʠ{��:�`��gU�[�d��S�]���v���w��\�f��v�w�lJ�s2�u ],��n�n�����a����|�)������a�S�G|q��a�`S�p�=�9���,�[c-����:zm�c�3Q#���<Fb�s�jG5ཙH�T�-��4�Ri�cH \�H��t�_]	p�C��~�i�7��IZ�)4��&�;W�p����Y ��6�"(2�i��}���dC�}�cW�c\u�ҕ{]�p�5�o:O����`R�ij�2˅��a���Uc���L��tL�C���g��Z�s�B�ㆀ�έ-��{��vg�ն�%��w=W�;���v�B��*UڥJ�wn�ݭ��"F��9I��Fb��d��R�<#sr�_����׋#|��~��؄a�r�\��%UeY"Dq�3���|*��/��������%n���'���{�_�(6��n4��HbjIq��#৪W���U:�c�Ҕ�^$}w�49�2*�����K��7�f��w��/�|�}=�,c�R����y'�Cl�M�HʒH��/uF�܁��y�=��#�L���H�Aq~�|�6�lylq��d����^ךfǶ���:�n廷��0Seܪۻ�3���k{��
(�
q<Ʉ~<#��˟��O�|�ҬQ� ��Uc���#��r���4�dB8�m���Fb�q���f���~!�O���D,�"����w�>� "p�m�ۉ����!��l�`3�p^��=����F����6� 8��vq�T�'M�䑤ܙ�1��]�>�}N���hdJ�D{��	���|G�p��[1B�F�S���s��i�3|�6S�|E��V��EB��;{�b�$��U�#j�!�H0p/���t�w�02m�-�� �u�Wku��Q4�e�TSt�V�÷�ɆF�aO�m���CB�Յ�l�i��ݞ�0���d-�$1��o����Eq߈t�hΔ�q��,�\d����9ҙ�χv�����mȂ����N�o�4@:�p����?kӾyH�ZY^�mu��r$ܑ��S�V#d���Z}��3V�g���OY:)��p�v�GXbN�%��RΑެ�u�OÇ�VzL�׍ȩ�`Y�d/E#�?	ϣl�]/:׮�m�m�.�ޝ��v�ݩ����d�A�@�-������Vݽhۢ[d��� �����,6 ���8eN�7ɚ �K8Eڭ�lF�k�F�Q��)R9�K2�}�#�����h��D���J�W+�x������.V��Z�	��{���[�K:Gz�o�ם?i���Hȴ�)����x�64�D�,6���'T�-Sw�X�
m\,�r�|mL����?_`ڡu �8���3�RIv�R4�nE�ھ�{�)�K�˗� ���ք�j��}c��7�O���l�UzVSb�zwnor��ծ�@�+Ԫ]ۭ
�sו׻��8G����U�4y�ӽ�m�󕹽�W�ػ�8���:)��-ehZշ)m�k`��U���,�өr[���s^���[�[҅wu�l�0  �e��T l M��l��`�*�T�P��  U l
��6� wl
��~�
�������0{�P6%AT��^�S�W�����ռoX5��;��]�Nw 
���G�aU�"@�j,[��~Δ����y ��>4|F��2�_/M�G�FE��f��R�RI$@�T��B�)��/�H��W#ܰ�S*��ㇼ��Xy�%R��0��e��j8�`��#1zY�_l���9����-w�������M�Jb'$i(������΢tSۋv�Rψ�V$�/b�i�PS'A��m�Qq�&i�K���O{ ��B���_á�M����Xo�������.:������=ۛ[wj�W3}�s�;ݺ�ť��MYsC�	�UM���d��t��G$�6�6 �zFb�sf�|!��摘��,�|�i��W�D�8�r4�e��<^/��#��U���3��tSup�@@��Y��W}�A
q'$�Fq�|:^ҳ�>x�^)�eM�,�������_	6����݌������N~�O���f��^�K?6�&y�����*����}�7j [��+Bb�9�����{)x��i�~�.3�&��Y4X6�P˒I#p�܌D�d�X�#dqBĘ�9h~��	`Wu�(�
� ����Rrͽ��]�{����11:A{��E����i�SҕMCf��qޚ��x͕�t2�I �
�\?tVX��*�Ӆw���rh9e8~�^�<��N��X�F�R(Kl9
����Kŷ/�}���؄�5h2��>?{��>V1�`Y�fW#�&��I$�eYA���\ˏt>4~�Ll�W��9���t��)�J���N~�H�,��*�[m+o�2%\?tB�]U��=�ڂ���:p�����~ID��6�m�T�v�^��4�M��:��ݻ��]�7nTU *l�[Z�y�ͻt-��̘5{��Ɋ�mK}K�0�^懰(���o������M��d�$���Q��h�v����M|���=}��̑�=��P�1��M��m�']�pNN6��<�=&���9����}p�PHL�'$,��d�����n�F^��պХ�9�e���,��q��q�����l�=���B�M�/p�Cd��OK�U2ۤ�%_<X��rK��˖.��r�/u�[<�sU U�����[�8wP��߷��yT�\�����|�:mB_]T{����/�d�&�m���{ʃ��'�N\��F�&�����/v�1�DmE���hMSw���5<~�/�|��S��D��{�5��W@���q{��Tb4�)�ٍ��!Gw��:o��I�F��*���u�,��;�#
��U���i��h��\0�$��N7�?a�Ӷ1ڰة�h<�N��O,�C����)��Ey�~�I$mF�I$< SJ��]cgq�ob�9�]@��%���L-�OIqm������V�w;�˝޽��1�x��]��
2yY���,����{d���;iٻ����0G޵�nr[m�ٶ}h  :�0   e�.��Gp`m��UT *�   p p6� w*
��_�����mb��T��`5�]ٻRı�R����KL-L2!׻e���*8\��x
�P�6���R���ZBdi0B|d~0�<"_b���R:}|�8l��P���qx� ���40���i�`��$�T/�#uX���:}�1��c\h�tt���6x�
�s�)dR0�=��D#M�܉H�l�9L#jӃ�=Ń�COO���M?-,ӇHºlӇ�8{���R�(�%��YH��E�>�<#�r��L����P>6G������0�}݇��%\�I-R��s:sǧ��d�4a\2�'?q���E���'VNp��=#n9"m�#QIOY���o5��v��{��=�[;�����*�M�mmki�fm��8���̥Ur-0��1Zo�#��������=3"��YNF٥$�i��i&ܑ�$�x~��3o�x�}��pKtD,���R�L����P>6Gu���,�$�J���4��Ѓ7?X���#�]��:}�q��Q�{W]�T%&j�m�j��}�l�9e>�5C��`��"��L�����t��bk�����TA������d&4��G�9����MWfE�Y�G�<l���.G�:fo�b�2Ia$\�IY"�[\V�(��գ21[��l���U��m��Z�j6�m�Q���:��'�g�8k`ӞZx~��Җi2��)�S����sR[?@��lk�2����{t>,��.��Za ��7#Nu`���Ǧ�$��0��rIv<i�?Nk�<C+���=���Su������������Y��g���}�f�|�%����g�7�Urܹ,�ܒI*0�/;쾋����E��sa�U���H����aώz���ڶ�%BV�@UR�~r�c�Z�wkͯi�[;��r�p-���,�?�����e��Y�34��=��N��A�D+��Oo��4�n��rz �-��1�^`��dt�r,0�ќ������j�5�0i�-<?^{	!��ʑmFCN���2�~0��둸�E�Z����L#v
嫆�6�k���.D�Hp�0�9՚}���Ǧ��4�Zt��]0�ߎ�ynt������[&KF���2�sv�O���RK������3<�!f>��USiq�<�M�S����޸���n��^��:�����T��6M��Օ�g-�n8��4��8����픳H��aM4��پjR�t�,3� �L#�|((�n�t�l�Z��@1�+�dx�c�e\ q�+�4||~�W�>2���8Q'�!%Z�	9ӆh��R����"��l��k�n�zB-�d�I#0�$����}�#�練t�-Ħ�~�ﲳ)�÷�h����*7#��'�>�L!i�}4���ժ����{%?i�7g�v����x�}q�;%AC/�PP��<�^��
.yYJ��1�V$E�qJ�4��Ri�QS��.x�1�*B�1T�����|��~�_�o��2���o^�W����N���Ȩ(}?~:?�̨(xy�cѮ���������T;�p���6�W���Ɏ,w��RXQ��,*$Ĉ	UX�U2�d���EAC�m�v:<�fד��PP��˷�~�]^���<�gIPPͻ��ǧ��
����(xqa��
���_{nƪ����Y�ty3�j��&���ɣ�ɦ7d�u�����?��Ҡ���6]����{=3��kL�AC^�yPP�׏Zc�q�u:t��cN�ݟg�&{xt�1����?,�5�ۿ����Od�(roٖz�hT2�?�է�Ƿ?�1AY&SY��W ߀`P��  � 7'�`a�>���  �J�;m(�  ������n �f�Jd��
$v+U��C���۳�q�wCwsm�j�t6�b�J�z1�C��B� *�(� d�P ����M*�YR�
m��Ѧ�Q@ �     y��E �!�V�Xn�5�f�r�i��bi�ۛ����K�wn��ng���l�.�C[wq�;`�Vtv��!@��iŐi�y�����9� ���8�h�=��ƋcW\#�Y��g�1���j.3�{یٹ�s=g��z=�Z�wt䖠t
��ds�]�{��M��{^�y�����7^z�Wom��u�N�)�6{��޽�gy�<����Kx����E�s'����F��p�נu�/;ݫjmj�Ey�q��`�n�-�($Qx�l�ex]o=�h�d����ƺۦ���x�7��v�v�O.�X��Xn�p��{P���a��e���Ề
+��4ҝ��N9a�� W� (�Ӯ�z�x��^��N��]�o1Ҟ7�Ṟ�8�v�K�WG���k*�g��Iy:[�w�w��EO+��4���QH��m�����\n��՞3\MR�#����f�G^�h�W��ܝ�`��ޞx��
�2���H�avt2�2���+�x�M����4mwS��:�{y�ۧ��Av�a�x��M�$4nu�qu����\���^6�,�ɧ���]��{ڀ/��nWJ �s����������:��=�zx����w������;tz�g��<��cu��9����l�p�h(Q $�n=�Wx��wwmu�E�c5��i#pS�89۝�=��q��v�l齽�w<`���뫬��������p��(	X�j
��Sh��۞<e�N��K�vq���]{7cw���=�{ٛ��m�]��ٷn���vUu���� ��)U M  �~�R���� �i�d� d��24��"��@��Q�  )�H���   I�@��$ڍ4 M���{�O�����hikk�zm]�(בM<߫]��I$�}��� I$�$$!$���I'�� I$���B�I�z@�I-! I$��@�$�Կ�[��_���ַwX��n�� )���GS��&�F�hc-�m݄�j�J�3*�����̘�P���,Q[��ڟ`��<��TQ(���T���{4R��V�%IIxB�U����Ke��]�Mf#bBu7m��c�����ӡ/i��0Vd�Ye�k�c�5��`�(�����r�1B��Q(��̽����<f�Vt$D4�j�$*��A,eQH)��D)�Ė-QLPQ`�J-U"�Q
ʪ��P���8�dQHެ,d�����X[ڠ)�Rq�l
l�.�T�M2Ri��!�Kv��T�ʺ0�g9ab���!i)�`)�3���.�nP���suz3�p��ܡPĆ0�Xu!IR��
`5Q�$��e0Ƙҋ9wj�*�ƚJB��5"�J`,��.��JR��u���d2@�TR!UJ��InT
t�q����bCL���&�D�R��
B�mf�Qf�P��j �C���4��CM�
N2`m���T6��@�!�4���'B�/@�Sc!��H,2I`hd4�RC�
d-!�"�L���1z���e�-.��U
�m 7T�heLi(uV�����`����u�RRS!Ia�4��
E;�-&��4��!�����d��Hm��G�L}�l��Q�QV���w@`�m�o鱄oZ4i�T���x��7iѱ ��.�`;��c���m��8mтhCxX�Cf�
[t����jX�*��e6�{�MPr˦�}�� ��Q�[E��Ud)X����CD:uJ�$J'n(��+�wBU���E������	�������]<A�7�C�@��4Ч֫Z�©���ju�9K\\��eZ���.��QC�<xq��w@�F���B��=[��'r�6��^�k�N�#cM�6V�,5j�r��Lm��G1���«��Z.d����5�h�V�l3u=�h�i��]?�,�%I�Q���3���/Qn�F�^d���{Z�ٗ�hwv��"�P�T��k`T�r��+f9�t�lz҉BF��JK已a�e\��wjaD+�\���ǀ�.�:�p�U$;�Y$9
�y8X���3.��������<��{K_��
��*��q�n�K���c�O�"Ă HYH�q�Kx1�͢�ث&c�%؊��C!�
CvV��t���Z�2��&��ɥL��k2R�:vܺ�����!iۆȤ�I0Խ���{h*�͉�����a�u`��V �LM��K8��Z�����*�y�:K&J-]�4+)����J��t��,
Cn�R�vV�ټ���7�WA1�K�=��v�N*�ܥy��#�i˓e�Mڧe�B�33�f�eU�`1����2�V[̧ͨge��TOc��T��-�Q�2c����*��L5�Z����B�0�{F�0�܌'����2�G6;ř[�)m�X2Y�Z��)IW�V��Az�KT�݄��XѶ�Y�nA1S��,)Х��T�Kbv� ࿩A䭀�Y���6h�������Jx$��j)d��כ����}sv�+� �S��˨�\�`=�sSۿ��7%�5�����ɩ���(m01�=�����Ze6��@�-w�R4�j�9�CO����l(ŷ�@
:�ʏX�У+W##
�/0B(�2�$�8b��)��ʧ��p�cve��#�]m�X��m
P&ͥX���C7V�)d�T�᫥�u��N���=f*�nŊ�Sp�	:�iuy��U�$��6�ͻ�t�3]���)����*��ز�%���j�J���ڱ%B9�.:������d�w-����6��ֲHǐ/���Q�N۽���խʽ&��If��2�$1n���N�W�`&q;�94�;�D0HW`�
��0r�Y�93E�3)-R�����1����iڽVjG���{V�;��
h/��kB��+����,6�R��bKh��@��V��4�`�J�[�*�̦�͗VAO%��[J�M��j�N:q)^�C�q�8�p	1���vCW	)؏V���R�R"Qgq<��8���+$�;�9yV>�Y{J�j��*�N��ZY���u���Kmn�*cӋ"��0dݴ�Jze�G�E�lɹX�d����w�5�ջ��V-hӹ$���˥d�D���B���Vf[sK.غ�X�F�.Z�{N��Z�[��!fګ�#u̌QQ:FԭsA�˫����`����pBp��s��fb(&�JP��oj^�^�S�ًe�]�e26Z��f�?e�����x$�Mc���� �L����Yk�'N`El��!���6�����B�Q��D�6�:�
ݨc1	d">Y4�j����S���[S*�(�E�H�����1TT\k��i��Xi���i��R���B�Jvo^�1��A����Wn���RMQ@����hQTP��Z�Y�Q�-Y������w���8��'H&μHm�@�^�.��J�̸>�(
b9E��tB��6���,d^3}��> ��X� �@��LB�)���p�ّD�pq�  �
�o,@���f�Bf���b����eīhF�ە�$`?̄��!RBD��e�#RJU�	6�n�wL�2�a�Nƻp���gh(c�ݘ`eԺ�a}ޯ5�.���ފtA5T�#ġ�{EDL��A�Ս��Q�5���x�!S$<yL@���@��D@P �#�Ѝ�U*@��-�M�~�(�a�͌�8)fԩ�a��Ifԗx������i{��u���^7`+[b��ɝ���u�Rj2R��� u��¬aWcr�\�F ��\n�j�,��59����F"��W��72�`��(X�;�&�(6����F��t� ��rS�l1�������j���)kU�cτ�Q�Ʃh�[W3fr�E�(�I)�N��H���`��j�0ؙ2�-[�l�t4�Q5��t�pQB��y"�_!Nɭ���� w��9�7wV�8��(4�V�6.e�]m�B�QP�ʗr�2$��M�7W����V^�F;�^UWu@u ���
Z�Rm%#UH��aJ�H(�Wζي��B�M����n����a�ʎ����[�ی���&���x�o;YNn�=�H4���BZ[O-Pb���("+�ed�8Q�4Ja�\�M4�LiXZg5z�E83�UZ��]�W6���6�*��[N�����[�B��2эo7��B�t���@�
QE�)v�S�IL�7�4�2c��H�H�w}�iب�wT�CI)�m�0��q�eShi�S�F�eJ�|�tK�y!�P	4��)d�D����GE;��)C�wԤ�����yE��h�0����Ŵ�MCw��&)=�Ib'i�Kߞ�Ǘ�@hn�L�̔FE���S4�,s2�t�Q�DL;�2=7H�ݣ+�,�;����7.��t�kש���h�������+�֠>��N6aYJJn��.���N��jś�B�m�z5e����/C[-e؈f���ͧbah�����'
�:5�Y�&���Q"����M�ψ��B�%��TT�5͌%l<��R�P��DV�stRxQ؋�R��u>U�B�]J<��]^���-��w���f+�*��[�n�W�4��7��7h�����m\�0�������Ƶd�P�k�jU�a�r�qJ.[!a�P�F����-�wa+r6�1�Cu��J1�B�?� Z��h�ykv2)� ьS[6�ͥP�=)�����BWgQ-<б�mӫE^���F�լ^����ɚ�o$�`�vH�KA�����pd͹uy��31N��9�K!c���`f��5{P���&T�r��ha�f��F\���䛑���kLf���vѶ��yx�E������y�.�S-V^�pɵ�bX)F�x�W.a�&�8'De�ڦĝ��27 Ɔ�5���2�d泖���p�S�%̶m��z�˭,�^��f���FTܲ��8�]fjB�6wpSy�ػ�Ȧ*�y�U�� ܸ]�:��;𩖦9��a����������
7z,e��Ȉ�J�Olje����6lV1Y��T��Q�ttMq��yJ����-�M�dQf��1:f�AM(� �C���S�E;T��w�K���&�,����B�#B��b�d��Ʋ�B���m�W�M@�[�%�r=�(�{R�[�X7x��������X|cyz3e��N�dǆ)��e^q˙W-ҡBe�H
����>Q*(��e�fM��.P$[3i�ʺ�4�˙�9{�`���-�vF�DN[�A��)�q����Hn]ŪC� ��"��L�]L�"�z�U[��P�V���p�k;�i�E�ʴi�QV�E衾j���n���:.��kQ�%*`D�fn�8�B�+s6^#t�XN�Ȉ����O ��ZWIc��z�u�:����s4B�[��h4�l�YMJ��^���˺ �3*
R&U����`´������BMB¬}1\X��Kd�ܻ�5(U52������ދU̗��#�
���o9n�7f�l��X��b�5WeӐe�G�8&�ȉ1ER�w��Q�`۱oU��B��{V���*�� �������F�3k!L^k{Z�5�@�;�]�B�Xͪ���*��G�B����9ZVn�j"�qX�ԩ���#0N2)�k.���]E��.�j�����VM�*���Y0ս��#H�ŧЪ�ԑ*�Q�j�"=z�L{,̨�PZ���Z\pX_@9��GCz�n�o�m��uÔ헶��H���ͷ�e�,7C�u�E�w2�)աSNE�B+)�s��x�@�^ٽ��r� m��q���AlM�1��(;�����0^*A3x`m�r��L�;����*�M^ �e��x$s�v�9w�*`8gʰ�$��)�y�Xh H	��7���,+�Ժ�����/$�&b�ʰʌ�jo�f6�8�57q2d�	��D�EE	?2>�UP�3�K��R�0-���N~ɡV�Ɉ��3j��[[%��:u�U���9�!�D���1���T��b�eB��E<T3o��/Z�h��&7`*m��E��,;t%�w�N����EX�t�xf�͘�=�YJ���6��N⫇(ަ�G�s���Ơ�� 1�Z���%ܪd��C�9���P�n�s��o(�N�Ԫ�(�J��S
�Ji�R))!ı�HC#���b]�Yn�fm!9��!� E�y���Р�ڨ7F��a�T��&�'��"jD���mt鴛ʕ�2�#,��X��[���Yv��܅�����,Qu��34 �EK:�w�/7s�eƄLwz�fV˗�4gW����ɜ��ɣUC��
ә�J��l�mb�^`��R� ��څ8f�Y׋7ihM"�r����Ų��5sV��Pu1����W�V6��;�!4K�i�U�Tdf�^e$������}���H�8�H�q	�5S��F��m歱��q��TA�X���Z��2��#E��ʲ�؂Ԕَ��<��M��Q����ԩ�[$,ߐ��R.�.CG(�n���������5ڥ
�Ouk��z�h9��0��"������@,T*��'E����"[wpKc��QX�Ŋ�vC�%�T�)w�vӫ���6���fhR��	D@V9�(���	9T(�ʣY�k���J{t�Yz���B�Z�l<�(o҃e'����$!����m^�io�ji���,o+��w[0Qs,V^n��C�0��v�"U�� �MgX�Q����[���bӧ`�R@��E���Q�r)$TXhJ��j��hn�:��߲��իݡQR�	c�Ѩ�8I����̭�St����Q5&��25�S�r����� �l��,1�w9QŮ=qG��$?Y�l�x%Y�mP�%��	<���v�ܘ�8pe��
ҳ�3QoT�6�T2��ݦ#P�+)fK�t�Ѕ�7�R��PP�D�.q�P8Kw1�T]Nmd�t�^�Ub�Rt�IN������F,�ͬ6��k.��-w-�^V2�4�	�LZ��Y2ŽM����r�Ɩf$�NhyX�G>�R-8�� M���M�0�yf��4Ж�$o�ݨ�S��omV0�I�X1aY!kv�PE;;,���E�Q˄��R�m+"f\����+����-]ݼy&'r*�wawI�/7�T`�2�S6E3�Q�"Hu���<��b���{�:���Ϊ�$f��ٜ��Gm��E�+��nX5��q�X��ǈ'@9�G|��wwt$���t�dկ�|/�l�'V��B}T��7YD�!ۓ1�3�-K��'H��\��s��>J�.[đ:�/r���1+���I����m�P�n5\���(��I;�NKP�O5�I%$�\�G_|�/�}$JS��u��m��K_,��]�R! ���܈V�y:�یU�Me ��֡����X>�3�2���}�S�9N�Q@緺9��b�h]�r��v�WyUǺ�sԕ8��אr���pOt��K�n��j��D�1vN��Vw�T�]��q�3��֝��;U;4��8QЈs
��{��f�*��M�8*/5�
�;�+��Gq���X*�3�}�,	ݓ�# �r�x1�آ����2����%Z�S9��m�dmsm�&a݈�Λ��4�<�D�&N��LK��I.�6�1.nI'$��|�Hy�ʖV�%�ηt]��}\�޾�-�%�T��)L�I�����Df�m@�YJ��{���fB�����gP:o9|s�F�Y&m�o�C^�5.v�^ˠ˖�s���H�*�<Df�u�wFg"�f��4���%aYv�A1��*��m^�GF���Z�7���"huq���]�O���藒��n]��O f_k"����>�F`�u�)	㯉�¤���i��fSr�]�0{t)h���N��M�cI��oYT�Ep�;�5B�Zz���{��'��j��-�d���(�n�R[��c��N���;S��.��'@ju�/z���uYO7e��x�PV�vj�P VY�;swf����>����-ͤ�\�8ȑY�ݢ��.������[]3t�ջ���h���2�:b�!`�i���P����!ڍ�j�7tڍc5 ���5v�uF�}zc]�ݹ�9!���sV8�,��6�)��ԕ�v�g+DwkkR����S��IK�v>|hw=���d.���ū��X��X�7���RL;�WJ��{d���dAw8��-f ����U����2Y�[&��/;u�"��t\hI�4T���V�f��$_b��Qa�BD��qW��Vr�Vt^N��_P��1���}s+����{�v�����+t�a'a�oD�����bv�W�n�����Qв��uy�w��z�e޺"c�J�)�/PN�7��{l�N����H�Y.e��{����0\��U���n�	 �N�����)cM��{���wB���Z���
�����1�b�sQP�/��0)���c,�����nSv����Y�R5�+��p���e_s�]�yj����:��Vze��l�nY9&K
�<�<�k�4Gs�B�M:
���.��VBI�ܕ�}�"WtgfE�v
Ցͽ"�U]E�
4�W*j�w��@����W���(O�G��|nh�|寀*�p&t��&��}�֡��󝓅 S��y��F�r����5�z}���[����evP�{����N1u;d�t�e�g����ұ�3n&2�P�8�
oO!i��룙A�*��G�"f�A�n���Tɽ���=������֕���w��
7��,&���5�Q�ߕqn�{+H����ϡ�3��-(�=�|�ʼZ�Q]�wt�Ǻ�]o���E#��IR;t�vY�N4��yWt��MS��(��WD�OZ�ܺ�ڍon`-ؽԘ'(��t�t;(=*�U��E�Nu��κ9Nws�r�MS��D�4���D:g)*2���ZR�ArE�(�;睻�-��Q�����9f�M\��=Ηt+�2�t�Ύ:�J��ʌ��q�M7d����AN�9Եi�+���ݚi�\bEKmZ���d��1�y��4yNޔ7�r�Fc��҃�:ڷ3�(�n�nq�1%Z ���0bJ�[G NN�{ٌ�d��:&�=Y�N�סiM�b���h���˘V1��kJ�jIEdPw�;B���Oc����`vYO�N�B�X�fӫޔ��#�n�0_r3�2`:G2N����Wo/��!ju���	A���meu�z�����4UfM�R��V�>\͹w�pt��'J=]�V�$W��\��2̣{@���٢��}�/�y�Ò�Ჴsg�֋��f~����)�=Bү4)l����՝��Kb��`��-���9����h+��2,F�;,#2�� |��f���,����^`�K�����6�#���N��t	�����޲����z�
󹓝y\���z1�.t�x���Fg���W�F�R�'.#)V��2��2>��+�q��q#"��X۝���S]1T������fJ����q����\y�	��aXIvq�iI��n�M�4��q�[��
���ӡBQU}��6Q$�ҸB�7�wN�4	��umۚnޒ˙Mow:��K9B�X7�ٱ�Z`F�/s�2��pt��uы8��><D�5&B�w풮��K������fn�2�[�[9�R�ܑ��W2�YzTqw�qEGo]ޛ�DU`�"X���.�q�nY@�n�t
�]V:�ܱ�#n�]����0�:G6U�}@��ܾ��:0���j��73_=�ҝ���P-Ƚ;22I�Ӷ���oLr��\]���2�sG�W�n=U�n>��=�ה���NZM�Jy�f6�䑝�{�'G�ۢ	@���Ϥ���.h����=<�T�$��s��2V���t�7&�c;�5��˸�����'f��dڷaw<{���}3}�ÑƩb��܄9�ˆ�����T}�kg)��M�lq=z�#kz��ff�cxr�9i=9�ѥ���m��;�r���z��,)�l�#�����f򫙷H�&�ɂm�ks��mۮ�*6q���#����WY|�/P�J�B�k�˵�#���r���pl|���Զ;T�{�V d�W'���v�4��t[[!v�.��X�i�����(V��ٴ9m��N���ڬ�z��A���M9�\��i���T4M�F��.�_]�#�$�;n��6l�;�Y�6(�7$\���ȡ���&n0:��h��u㷠t���!��)���9f��ݘ
ѕݫ [��a֣�ɖ�Xԁ�� ��Xt��7��K��etq,ڥ��Ql�
'"�Vۦ74a3V!�l����Z)6��|�|Ԧӥq��˙�wړRY�:��mq�쭌���|�3��of�n��'�v�4R��mN��f��zt`2�ۏsV�n��'&���_i}[�V���m�ya���m�둪�tQ�P�����Zo�2ν�p̼����0����]
�W{��P����A��e�0�k�b��ؽb鯰�d�=�S�x��.�t� �pm���Wk4|OC��3a:Q��ٚ.N�O��naMf�}�Nv7��y=H�A����3��NK��޼@�j��΍����aXpͺ��\��������H&򠡽�����2�.�+��R7��0�Y����R`�wؕ3��Y���[��
���Pt�h]w���S�k
:m�8��81;�RΜ��n#:
Vjf�M�1-���hQ����,.7F�_�4c�;o��x�C�]:;��B�*9�u�
�zN�ɍo:2������2/0/�&&9I�-�½�/�&Uj�)pgk-^���	���s�l�sFr��̋rJ���ɇz����Xyדz!���������I���'s�E8[��]u�rDۡ��Wt�c��F�D�Cz�u��%�=B��Ycol-��v��O�(��2���2)�I����d�J����%m;�N��ϵwJ��n�B���̈6�N�����F����\���s��L�f7z
��|[��z�ŕ��iLmS�Db���4�TO=�k9���Wa�U�X���/m7C��1�ّ�������ٛ�Vr���w��ީ1v�u�	,[#ur3�w3�Zku�u����$�[1	��p�Լ��Vd�ۘ�Vǵ�7I�F��Ծ[w)-�����ɘ9藶�\������7��%�_n�f��,:�"bր�Wv��݌��%��1�oV̫��WY�=ݭӬ��\���CU�]��E�Gn]�ghc��:6�P��N��I��ŋ���RJ2j^2�1N;�tEo<1����b�a��R�f.��}Iګ۬0�'L�38mX�u�:*:R�:�z'P�E���Co���S<�fۛ9(�����4��*��y���B��w;��R�"_d+8:�dN^&�r���Ǵ��+�P²�Y(lDjw`SU�YR�E�
�1>���S=c�n�W̦k+��9�U�I�R�y�����JC��s�k�тr�Yh��Q_t?�J�{t�t��əʦ��r�h陚�S'�Se�(o
���T}�[bS[�k��h��֮jճ�v^ŗ�&�[*�=���j[����T�N�ٜB�jJ�us"DH@ʄ����.à>tc~	Q�:46|rfGO)u�z��w�����j�^8
��/2�s\tռ�X��(�7p;��Ir�Z��G��g'B�J+#wY/x;-}n����y�_G;<��+��ѓ�c����6c�6�wn��Je���t˲�fw
�d�љ6���ק�ꒉK�{�\8)mjx�DQgYd�� �`Ҏo�`-=�Ŝb�X3Cc�pnU�L�=MT�d��u�2�n>��N[y�.^Z��.��h�Y]f��H���uW�\��q:6fV�Y�];̒����u�rʔ�BZ�1���.�5k�yoY��LG^um���X��K��$'�ݿ�4S�6�N�'��`��ga�'tIī;�:��q��`L�/��gR�v����Tx�,3�$^���<>���
U�ڕ|(�Ǻ$��N{ݛ��Y�F�LD���c_5{\'2�;�{��ۭ4�b���7�-��J9%뮏U��k�����N]�PX-t�ͅT-�����=�6NYA\!:��MFLJ��\��P��wm�\ʗA�I�X�^|�nox��a	F�"ER�]��!��V�2�_FB]]�5w:a�z���lG"v���1skc�Ԫ�}݊��8�G��F����^ೲ���[�Qܓn���s��C���y�<�˜r�;�'2�53:���QwgnSIy�s�42��I��2�J�[�7[�nۙ���&��F���Dd�;����G��5홖��y]3�gTc�.5u8�0�Z^��k2G�f���SZ�MlCԓ1J*M�kh6� �:�ּ樃��[�&:����_�}��hg$109�9��yLg �S��+Fa;{y�Le���Ӂ�vc�ɪ�������J��V����s�!�l���ንfc��7u.�;9�l�c�Ncqd"5[�V��ͺnKɛ�5�+����S���D1��KYV E�Vg<�.j�%��!�uIp9�T�ɔ {(�El;�.fa$AWv��]s��k����p_���F$.���+�R.͕دG#�%�Ѫ��up�ҩ�G�ŝ��{��	����r��#ȇAL�G[����J��uD��
��������;(��,�*[Y�U�m��]Ԝ@��v <Vw���3����Ι>�y��¬A��T�Ѽ+T��R�^��
)g��h���꺴�յ�K��R>h�tܬ�G9l2
���Z�����:��� �JC{��x�j�d����sk��[h��f�vp��D΅��WP}���5Ӷ�9�b����d�����qOx6�Օ&�ǿt����T��6wj]缯�y�!lV�Z�#����.(kJ��
c�q�Me���K\��_'-�_J�{"�ع]<r�ČNƍ�*b�S�\/��^27(݂y���Ðf]>��6S��OwjqI��Qf�] Ьޅw)���g?���..]��#�+Z�t-�R6(iU�glod4�k��M���v����]�t�p�&F=�v�+x���1&�]����r��ކ$����G}�tv��.�I;���vb"��2���G.g�7ٔ`������nV�v�o5���2��Z�[&���Ǔ�S�$�m�uk
麺��cfݸS��9V�V��y�oWR�p2oh��c��;�Hy��+��툰�{�և�p"Lj�}�AiXhe)K�5��(��č��=^8/�&���AԤ�ӝe����_.�����V^�}VOa�f��jc;�Vrշ`���P�5�WS�޶��,Re�S�Q�޹%�ӒRZ�yc$ɴ��1`��m� R�m�e  � r      R&��6��c�J ��`  �l  ��  � m�m��        R)m� m�   ���� $ ̶�m���l    l�      m����411��a 4�r�I�          m�                     �BIX0��@    4!�         �!�� 6�    �I�*E.d�  �(      m� m�             ��`   m�  �    $�C` �`                                            �   6�  6��      �1�� m$�m�4�6��`�`    6�    H      &D�    �u@               �m�                  ��                       IS(I@�dcm&H��C��̀ "��2�
��pᤡ��@ L�$ m� m%26�ll �Ls"I!$l� J��HCԒ0�%��)�Id�L��S.XKs$9��C�h��     @ LH4�      �  � �   @        6�ffff7FP��B�I��	I$��$I	��$�L�+���՟���i���׮[���{ĭ��mp�dO�'[ݼ�;ԑś�_��n.�[RFVd�ȸ�zh���ւ;.i��Jj�,��軡�7c3sA�+2i�V��yJ�|G,ᙢ�c�њsPȂ��	ıt=�(]*v�`�S]1C_���̊u(�gd܀�To�[�vR�%f<=ϩ�UAS�UUUE�o]�u�U��:�%�;	�K.�y��}zs;��ޚ��M��ͥ�p��� �pm��]:ފ�Y�je?��|�׮�W�^Z,��VX�3]E�E\�\���V���r�Vy��}n�m�v7���ΎӐ��j�K��Y�VL��X���<r�Os��c��չ�z��um�eDݑ7q���@��vu+u�S
V����v�o�?�V�o�Y8Pl�u��cH��,}�{��_KK#�aM��W^{u�w�ںe'ua'�wEKZ+�W7� ���踊'r�#U�����E�D����5��c��"F�ce�\7^�"�ྊ�ʜn�Do��7�M�\��v��g5{�����GE�ujU�+�o��DgP]��p����
ʖsJ}�!w�sK(ғz�oG����72�=�|3�=��S$��"K4�����i;��/�v�oW7Pɥs4:�:�;�vw^���W�L� 4�4!� 6�m�2m� D  HJ�         �0 e��     �              dC lm���           1�E*m)�5,�D�	!���*D���l ����̪���@$��ȯ�5�k/����ϴ�UAFXحlLa9�t�0����R�iunRٱ`V���%䕨GVJI�Ǖ��t������L� �6�$��� lm� 0
I��"0ؾm;��U	*m���{�2�4̳Csm΂U�E�#,�rü�{t�V��)�L(��P�x����mh�5�j��N��ێ�p�R�8Uȹ֧�Y������Z�#{s���*���T�Y�h���{�'+^���kB�[ �U�(�@FAH����̮�^2oe�kN��dj�ɽʍu�Y�ak(jy�h�����ܕis� �]�-7F��t��ٝx^�F���U����7�ݫ�ά�jN�K�[}Kj��m�gYD`�v�ޚ��:�!�ѯn�v�LA@TPQX �(}@B�;0��t�����͊��"A$A�PQ#,GG���V�|[� ���"�b G�(d�i���U�����)���뵗ݶ��n|�Py����7k�r�˥-¾�݇����#��M�v�H���Ϟ��2�ͫ��f�H�DtZ�w��h��u��N\1MڻT��ȡ����-k��b�w�.����^�$�μ�C�QM��6w*�s��Һ���$�}��Fwd��u�\ǔ�w#z�YZ<a���N�
,o���^/��P�97��l$n8�Xۦ�=�ۺ����v�-΅��ݡZ��J�]Q�[s�u�MW]�J�m����ݭ�L��^���z��	��hU�9f�v���9Ք��s:��JEyeR���y�p5���u.igE>x������N�{�O9�oyu�7�8\������,E�, #�6�:�sޛ[�x�p�]I1���s�l���9��}���)$X ���P���xG^c�:��*�S\\;O�Wt�yev1�1.����G�Q=�O=��ۅdT:�g:��K�bh>�����)�sd��ٵY׷u��ʋ��x_p��{G��\��m���vY�F�칳\���5��}�g�|O��|u�Yi��-�1�D��}�}��f�g��9R��j��36��pХ������η�F�fJ��L*��N8�)��r���i)�	�ٷ%L�$qz祉dǼ=�<;c��nj��������"���z��P��Bq�>��:�:'rl� �ΚYk��{]߼""��#Q`��b�H�Ċ*0�,b�"0�#I"0��y^��t���J���G:�p�OL�T۾�f�ݍz�����k�+�y��������
���+ꪨ�8ƹ�_b�]!(�# K��(oO��K!�8�%yq7Վ�Y����u���c��啇h��U{x9�<_L'�H��R`/{xõޒ�_t�����3v)��Ah*z*��L�{y�l}<WK����Zl�s9�[��qY�� �FAcV �"_���k��;�^�j���:�m-L7�A�͸k!ѧ�A�I�Z�Wu���m�+B������@͍RNL����'���0��q�8�ɺ�7]/簪�z��M;����:�$;��Ⱥ&ST�]�ذF
�Ȩ��C~��C㷽�֝���H�Ec?Da�ˏteS���~������s��x��x��V�N��ޖ�s��5L]b����+a��{��"SA�]�2�>�I�^�Q���0$Ru�jߵUʳ��:fe���*�tͨV��n�Y�<ȫgU�[� �y�7UN�l��k�J��t<�CI�@L̃m�hlm�     ���d9%Ȗ�}��bى���8Rڹ�9��\Ѣ�Z���+2��h�n��_��u�� ��ܬ��%)Ȱ�����^��^���wٿ� o=���-�!ҷ�J�I�Ƶuڼ�5��.��D�*��b>U����NN�c�CN�½�������|>��0wn�1�CE�i#ȭ�em�$��Y��l�d�K:�s���Ꝡ�6v�ܙ.�.Ƙ�x&���BNT�l�� }��� 7�v��+ף�
��E����)���`�"�"���Wy-�G�Mw^6xhs[�m�&(���e#'r��C��#��'Nd���˲M/�igm��t(��]��
E%���}�3.\��Gdd�c�f�yW�{��榘`�Hּ�R�W�}�d���}�����,D�WH判���p�^�
��e"��k��k5i]}ǺJ�.e]E)�2��1��� �%Mٛ5�.^�:���5�k��>��j�1E�`�Da� +~Ѯ��^���/]�}�Rs���p�,}�')�΂E�4������爽W�\��ؽ��.��Eo}��}�y�p�t�w3������]q7�o!ڐG�Ұ.ي@�s���u��g<1/x�R��U}5�=~BR���1X�X2A�$@Td���@#�X�E_j{������o��3.�3*��5^�~�&��H0~�
�Ó�;O���mk�h�K���mn}V˦<�������b�6G�5�,�3D,K���jVE���F�J�U}��{��+aήoG�Y�e雎��Y�4��S�>6�j��:�9�GS�}� ��\�B�.��ɝ��at6��SPȮ��>�{�n�y2��-V[�/L��{-	3�J��0l��Y
b������R`m_��ۭ�^�PݩPo����� md�����}�t���r�Q[l�ک�Wì6{a�s�ʨ�-y]���1�F�A�}�;>��}wm��	N��`79��T����>�׀O�?��N�K�$�C�M1��,ɉԇ@(�LD����>�j�r�ӎ���ƪ��w���0PET���E"EH�PE����1=M���s3z}�~��a�n{~��^��s�?�@�%�F��iy�b��E�7��C|F���l�ݝs̆.�Q���S/"O`�\��y6�B�Z#V���| ��Zo_L�W�T�;o��Hh�D�xmb���2��̈[{6�Ä�5˯��t,;'{�����ʆ�Q[Q�.U"�DyU��c)(AX�UT�lk �<�� |�k��w)48�H]Bi-*���=]g1��Jk��M%��/1_)Ϣ��X��	H��d�ʙ�#�������ξ	Z|%�����Zb����8��,�ڤ�;�E���:ހqX׃�-&5��ء����R\�u
.��#b�^��ﴚ���^W�ef�4��؛�7[}�1�JR+�,�Kg�'՞}��ɫΧs�K6Vf���W��<׭k/Z��N�PdA�
���$P�a1AQb+�,A��9�`�H�@Y�F�#2��G���]^���]>��v����U�a��<Tjpכ����ǵ7,f��B8Tú^^�]P�v�\�3vT�}�U}S��g̚��k��-�'&ۥks�\e�W}ϙ ���aR�P�8N�Ӟ��i���=u��TP`��X��|�{��w3~���|���H���*r�n�
����Y"��n��ԶV�hM���rIY��C���O��x�K�)�mp8on<����f�ɻ@�T�̠ �m� �� m)��)%ugdi��]d  WU�l�e>Q��ԣ3T��hf�������-^O��s��v72�Tj7Y�ٖ�}�h�}ܪ滦5��+fcR�m��\��J�p�n^�a�.�����G5�Fey�;�D��m�DE#"1�	 1U�,�"Ő���9~N޽��f�$�Q���ky}��7y�}��	e�D1湴�_^�����h۔M�=�M��Z�=κ� �\�Ӂ��F�9�~�������`\��a�f���'���;6�[U,���0,v����Lh���3Lb�*�`Kw3F^�ڱ�c�q.�2�n�G��X�B��Wl}�J淍?]}wX�r%n�M�Җu;w��,��p^����퟾����B&��V��^�k�GXt�����;�r���g7hR�4�����r�uLe<��!�/�f��v���4�ƼZ� gW5�q���.5عމ�;�ƨ�yN��6下u�����]�^���Owk���Wl3�����u�7���z�ml��	dG��׷i��ֻ�N�`Ċ�"(�T�R �)��p�f��\�u�׻��	�@���@�����h�_�f�V����|w%_A�_c��KҲ��x��kK�	�����ƴL�J��UUS��J��.d,t7$��m�2�?��	;1'wGHUD��$Kڊc���m����vH�k:ؼ|9r�0�9|�_V!ӳ�r���X뜥�h����X 2 � �=Z��>6s��^kM�]�u�Y�Ki�ɀ�Dޅo�h���чS�|+��2�wR����U
�cMnTw[Ȫ����;�/;�tL$���
d��I1���c$��<���0$4�%0b�	l�'R@8��d�y�i	��]�3~�N��w��9��ʱ�ER������
t�F��-ܺ�P�w�U���Ped���7�R��W��f�Y����U�����UB\7ފ[�Dzna%�7!�7[X8`�w�V��z��6�1�["W}�f�eшe�ק^�ON@M^�vͲ٘��v��\�Y��	R)�V�gIy���1�#+g%#�*1�M��0`4RU-��"fQ��z���:�0�o��A@�6���(BĪe'��s"���6�>�d�U)�U�h�;�w����V�њH��:ݙU.i���`i�3�i�m�zn����.�I��ru<�h�RH�D��s��5x5��2޾�E�]�R����հ��W7ۛP�����5�_�0��:�!(ҷ����%�m>�g�p�D%�2\�LN}4`m��8�O�F"2�����$���г31���f��笥�j�[w�n�J�-�*���)���o�aY�K@tGƟ0�{q�ܪ����o�{Eq9�)5ea�K���R��Yl
.��;��o~ki[�Bڮ��V�ʻ�]B���M�^��Q��]�%
�R D�M1�S~:./+E�U���V���Ve�C�ۯ��I,ov�����a��o�'�ow���]
�h���葰"��},���Fwwt8��pe�@i��k+�l����Y�љ;.�|�g�պ�yp_3����J��΍��8���yq���䤗�Rwlu�AV�s/��J�͊���� �3���z�N�j},
���H<yG
�͕�Nԣ����o�ǔ܈S��9|����n��tc��;�¢fr��gWC��w�%�Z�a�:ذ设��ѭq�;�:��!`�¾�n�3V�)�Q���|��5Ʈ�A�e7�B��<n�5�5�F�y�O�M��/����RN��ɝ�6��,��F�b��,���Ի�C��E_^���޷/��WY��.��ƶ��{��ECmـ��P���oPٕ�=e�����Y�N�ڒ��]�1p�Jm.��E���d�6��P�l��/��{��v�4-+���o���Yƻqo,,���N[��N��C�u�$�ZI�݄��a̵���ʸZ��kmM���Ȩ����(],t����ӻOL��csW\��=Y;!�Qj��n��!���.��=��1��DL�dɐ��Oq���ψ��5��Ji����$��t�}h]s`������^�ѦK��%��h�LB�q�oi��-Y<fw_0i��6���d���'�$ֲ��҄0c���z�賹��Nlї[�j�jl�w��o����;�5]���.�Z��_�sF+����+/�;�Ru^�B�<[�v��P����P9R[l��v�px��(��4�h�֎��(š6�A<뭍^V�~(� �QP�@R�Q(�RJ)�E`S%$"�?f���e{�
"��F((�� �7~�q�Nh��4��S�D��0إ�;�"�v�9}��}�ʘ����*��)]U]�9J�'�G4�s-�O�M	A�燨k�[	�N��+X���׾�<�n���r��� ��:�\>V��Y���-�<���7��*$c�3�h�¿
�џs��G��j߄*��X�r��r� �Zˮq�8RJ�Z����n�5^���A#�o�����x�)��w%I�����O�l�eN8/F�p5�+2;QHa�$f��y���zYM�_JW/�G���d#���B�FG7�Q�.L�jd�|>��>��	� ���������{yΛJ������H��:�J�|Io5_�6ƨ>���f���r�ڒ%��Oׁ�[$�lت�.o9�6%A�2j:f�K��2���{;�*n�
<�7
G�ЦI�b�qYf��t�Jd� �*A��"�� �#D9�dq�u�V���B)g?*��11"�
�� �XoX_��o�7��f��¢�z)���C
��<ڎ����xo�JΨ��Igyr�*�8�7����PG@H̅���qŚG.�>��nj�OH��Oq�E�=�}��;��E����U^���YO����kva�k�B���x�#��\2T��g�č�g�ّ�d��֣Btͱ�J�����뤶���΃P4�� ����}��Ǘ3W��;�z#v�(�g$�=�$[ʈ�U�˽h�])r����^���]w@�-�3B�2�JJ�.�hKJ��`���*�6Ju�x����\lnϾ�]TQ�+
mJ���Ew�˻X��$?UI�R� �� ���Y��Jz',��Q]�N�T}�p�c	�t��nAYV����H��-�m�m�x���:�fnd&%&jD�
dm m��`  H  ��2ۄ�$���.�y3��Yy���o��z?!����|�ik�����R��d�N'��H�S�m'X|�d7ʇ�-��Pm-"��m�7<0QX(($b�1Q@H(�E�QA�#"��� (���;��o���ߡHO6�z���'��N�z��wg�	�+�O���E�J�SAUUQQB��Z�AJ%P�T��U)
�%�Q�O�{�N3��_�$۶O3�L��%�HN06�ɬ���U}�/^!��RM�ɍ2Nꍡ�LY-'��rC��'>�\&j��=�
a�6��S&�i�
����K�I\�r+��H��&��>�H��z�s��nH3���������}5c���U��i��
��e-hz�*��uev�C���H�hf{w��!>M�{�����~��׋���2�
O����&�i<��4�`u���ćM�9�'���m��@�(��d�
ʚC��ﺜ�/���}���w�}�7�DE��1&�[�ÿ�uV��~�Ԁ[}�d�JHtf�T�d���LĜAƃl�$�k;K�{}��B|�����
d�GTN�b�߾�u��q����<�5t)��m&&"�d4ΡL&������*8   �S��1�DT��S=S�:�H^��A��'�I�$�	���)'{��~�C��0��q	�4�I����
�s���g���<HuT�2|�*������v�+�КO�B�����s�����G��<�>~JI1�NeN!J�JgX�$Z���Z��N�- ���Ϯ�e�m��':ECR��ԥ��V�Ӄ�#o�V�롯�U�9�$����vw�3�٦�`y�ԓ���;�H<���y����ѓ�9G>`|����LKa�,1 ����А�ho����C�<�N��EEUUR#0�Y�b'�s;_eg}Z���>@�چ�I�O'ܩ'�e�1&�ağ!��-��g���`�tC���m��M2_5�UWs^�w����Bq�@)?!�	_�x����� ~a�PM"����q�j�u�����B`��޻�*zU�=X�2~�|  |;f^�w\D)��-�'
�oP������;��Ю��?Ct}4�����+K�����$��A�w"]��:j�s��m���Y�����Ts���@�u�{������a�#Z�S�����VU�@�!���J�3�a�YE[Z�Ψ�=��{u�r!�0�lɭ���˔�h��c[~�CYN��j��9�_Tb�e�%=��|>|׽P|�d��Q���"ld�VF�4�UKx��*�)"^#N0���XI�|�bn���������w�LA�����g;[w�Mv���\Ϯ��Db �1�A��
A"
*$QQ��""�^�߽�j�b�*7g���<�d+�[��[GNO��{iv���+��9��v��̌�]\_U�]]��<��;}� ��5�����+���@��CH~��~j�+ҹ�t���V[��}BcM97#+:a#:��{oJpX�ɏ�cӻ�xۅs-�[c��0O�Q��Y$E��,*i<%�E�M��yz����ﾭ=�bz1�\��[�JQ55�;�vc\J��&��"Fn�d��J=�����.�j�o��;�˔����(2LB��g׶�����F�B|��Dq����>���""���� ���՘���+a��b��f��V��`q�A3t��	��)h������&av�O����������33���̎�n��][��#�l?&s�]n�L�}��'7{�`�O�g��+Ln4
����&b���T+޶yj�n�I�S$%
��u/Ѻ�l�Z�X�}�7>�,7{��N�(�.�����]���)cgw�� W�Wι����w�}�՛�X
�PUX�AF(H"EA@�	E|��^e_?g>�ۭ��x��/{@��L���\8�۟*��ݚ&���1�b���{�B�T{��}��ؕ����wĩ���Z=X0��N�I�Q�"`jo�)���ph[6�t;�dgݤ��=A�ࣺ�QW{:Dbm�Y/�U3���}�G�����_�b�q@ �a2�7���喔�yh�b;.l�H᫭1��<m'�N7���'�M[�#l�7ǋ��78=���Yg0	�Z��z���3W_�}˿�e�N���B�z����������I�*���9�6�h�kc�ݩU��Xk�]0�ٮ=co`N'#�b�=O�W��ٚ;�R�ƞE�>@��Ky��õ�)�>��c*���T�wWL�W���9���Tg�s㇎3�:S��f)q�p62��F
��,i{��yd��[��si�e��`��<����t~�!�B{���ႌF*���@c0�Ϩ��zz�N�u�����U+�S���y{�e滯��
5w���� R	����gt��a�L�/cJp,<�W�ܗ&C�rrVVi�D*t��n	un����Frn���o�=D��z� �@)��!�  �   ���0�K��d�#��U�`6�������r#�� �]��#��1�F(�A\�7���z�ʛ�N�������>��J>��^�f�����6���ڼ͍=\�ͫ\nU���KҰ����<&����������6\�n�ٮ$�ˢ��b�����9�O�0 ���p��e>���m�6n�]�v��<��1�v�-t��>�9���w�q��\CH(H�"�Է)l�s���;	��D8��8�-��R���ٚ�������ht\z2#��2wa@8��k}LʚA��Z��5��A��U���Yq��i=��F��[�\.���h�x~ݍ��M��~S�2q�0DX� �T`A$��l��ڙ(�J�D���I�~�\}�A�2�DE�P����eW�VQvk��kѯ�s�n62*��.8G.F�r�7b��CƩf��dOdօ6��pmd=[�:r3VZ}�?�!H�{����zu���s�8}{�O��S�s=J�N9aԺ̕u�^��30��״b�W��;�l�;�=�㬜�"�N搾Y�龳u��%����,(9u� �����jõ��B��ś��g1���^v�	Iv!j�nl&����f�8&x�]�W��l�C��`idC�z�1��:[����/���3UU��r}��5\C�"
�0P�4��P�)"�����*+U$d�PIQ
�I�z��ֹ��ۿaQ�D��;$�VR벝aG�ՠ���I�c�O:���OLK���]v���*9�s���O&�8\A��*��e��v
�F�u�_L�u\���lq?b��}� �/J�)>��"Ԗ �_GJ�+��"�h�3�k�73clm�=������K�}�8���p�/gu஗��`9��\VV�
�Z�v9��f�B�������g��u�ݽv�I o�A�� '�_�w���{�{.����ڭ��DUb�A*�(|��n��{޼�W������ߕ�É��][����7T��Y�>�V@�Sݝ2A*�#F�����U��/�5;�<=��o_� ϵ^�y	?$�$$�$!$�}����U]��t����[�x�yᔧNY׻4`-1��"����+m�ğB������L�@��ֶp>n�&9��څ}Z�9�*�_x�(�L�t��;()�8�m�}1j�k�Z�'����*.f��y���|��ଳ�\xvչus��˵ݟ�k�v�w�QU�ಓS#�l{�> ���<�ծt��GR���͒l�tp�l��n�W91�����W���v����gj7�O��隸�,g��J� $�V>t�㨝W�'����D�_�~�|>��tF)�}2�!���f�gdu�3�f�v�c�)r��\��Nnq9��3�gbrE�|�a3��<n�����I��n�O\�W������'ߤ e8`,� �UU�0Y�XŌH(#�}���Ս>�>���`��
fX��^1[�{{s�b��^ٳ����.�F��Os��*��C�����+w!=dj��X�W�ʎ��i`S�nV.�Q�����Mn;1����O��f�I�ɘnz	�RHO?W9��U��o[����<�\ۣ5���++c�����b�3e�u��U!}u�﹮��쏞�N����k/%�H�aB�,���2�F?RQ��p3n^w��s4E���).�F��.��}~�y�}�ʭ�s{����	�DFF10Y@�_zں�k��{��|�:M��	����+��
�՜�4���K+\��cW�.�Ҍ�wQ����s�g��'���h:*���ӎ�	[�������^�F��z�UUh�-n��f�ṗ'+��?q�C�ŷҏL��oGna[2�,�����ֺ!NZ�+X�c�r���5^{�[��h+,��b� �!7_����z�}�Mz�׭��I�L �~ͷ�^:/�=i͘�b�D'�1��kb�)5������ի�~������vR�A����"2_�O�ۻ����S���0�*(msQV")&��bU �� � �>�>�4iR�-y{��x=S=�e@������j)�D��$وk�=S*�H�G��Ɍ^y:'�o;�\X����>����n�+D^�Һ�7���3��|KHS)��� q��$'0��Mr�FXbB[$��@��s�z}�9���sY�/��c�o鞔���rs�BQ}�s�ohHp/d^#*rt1J35QHȉA��l��w�*(��ої���jT+W�_(:.46r����Db5�M�a\�5������/GG��w���	�tvv��0��:-��ZF1+g+QP���U�A��rȺ�ZYꃪ�3e�O5��s��7Гb~��/\��v�`KQ�ې�QEY�$m6�H ph�2���e�����ΩU�͇U�����9T���WnUЋ�M*��I|5*�Q���;��3���3��׫D�)�C����ahKp�]i[�����j������w5i;Mқ�͢�Nm����;w1���Z�9
�>�C�I
���n�c�5��
�W�һ5��r瓳�<x]�;�z�p�{�W)��%	H��48@2I5r(�ʛ����w��b�6�n	X�	܌/ `�����F3xգe�QA|s��s��B�ۇ9Z.`p�������+�	��D��"�HŇk��5��r��);��T��s�Vs��>X*��Z$�k@}\,r��-O*]ED�I�M�k�e��fR�V��]��R9p:��ܩn�D�8�h�	��r��(��� 2Ctl�����X�}5������c�]o{0��F�qN�nh�s��n8�8��̮����e���H���3��g,Qm1�3vU���&���5������h����3@�-In�!${�޺�nM��1sk�^���cZW%Ynަ�3Pb��<��(�$��5��{���(h���Qe�\ٔ[�%Pste��цe�hu����(���]������)L
�Yնq-��Y�94��&��:�%N����U��e2�Jy�G
����VM*���Iw�;��jnT�������wy���V�61jl��9��r�w� &��fŢ�˕���qV7/�S�,Us���q�s��Y4��y��uZ��&������x���-��ے�>��@ތe�i�T{Vd�7�)gx�z�W���-�32���5�AII���w%`�J2��7�Y.��}[f�"��gL��Ww��|�>�޹}��t���fL���vut�8����E��f�1؛�D�m���DR"���;6���'g��U��f:ݮy�м��5wv��6B^�֚��z'+7��Y� �%�IT��l B@      �cl`       lH m�" �m��  �m���6        �`  �`�   Cm�           (�K ��')��`BR�i�rL�c� 6�  �ǿL�U��~$��۫�ڥV� �e�S��V�Kى�����T�������%+�R��.� RrL����       b�(M!7�F�3�2�cr�&S��$����@�m�үUr��-xDQ��` q �몿�| ���p%Do��Q��Z��Ť=8��qe@)����"��7d�hS]���0�z���b�t\�
%�|�<�l[��k�8�.��Ǖb�K��dYw7U�K@��d�L�MK3�=�}.y��1�(��̩(�޷a(�nbi$�P���n}}Gl���q�ƝJO�T�/�2�m�ݐ�ׯ�������fd|_N������A�a�ݫV}t�YU�=�����D�q����	���Q�O�N[�-�s�� AO�A����AV�}ﵲ��WT��%�AR�q*�S,�������=���k̓ୣ2f|������&������U�t�9�v<+Ԟ��Kv�(8bIM"^��o�#��C���엿�9m0��z�m>E?IC���z�fn֒�����N���q��ƴ8��*�r��3^>�E��7����a�d��
:\��7w֧��̶�(���h�O���D`�ETU��b*�1QDTb��G�B��EX���bE�
����TD��Q�����Q@�DX� b"�UP�$B��DH��#UEbk�e��y�~������iE�:�F���v,��9�*w��G�x:� �6vAo�c*#QP4�dVM�F���a��uC�΄C.�~�� _��J�
�1�ldE%奔%\�)�s��	��Zk�#���p�S���M����s�����8ߘ�3$QnZ����n]�\���|9��]��б�!���T�p�b�C����}U|��Ж�=+�U�Q��%DƧ݌�������t����<,xAio`K�5���woA�I`��*qk�yF�U9���u��`Ҿ'Kz�񮲯Y��LǱ�Mb[m�>+��m?�@W���#FbH��0T�dX(�,I��x�$N�F��%��^�yF"U~��
҉;B���l'V�G�̪ѝ��|��qؒl ��K&:xN��IrW���;�ibN$z�\/K������vsUC<{��G���"�%6�x��GR��a��z`m�<��9Q3�wˢ-cZ�\��tv�E�>�#��H&8̄�w�3f+�,����z�L��j�W�T��WUۇыg`k��2{9��Д�*�#���s���֯��Q^, �A"��B��=|ϯ/{ˮ}�}�u��?AHb (B�s>�y�c+W�WVv�}q[Zp��2D:�� 8W8���:Z��+���U���r��ٲj��V0�b�p���� -̘Z��^�o3Ƶ�L*�]\B��B^{�u�sn}"&y�~�כU�-e|�"��](�o�"'_t򆭸P��PH�mCi*��9� ����|3�N��ǁG�ܴ�C`�d@�MűT�X�9ڭ�쾾�Y��5���겋f��0.�| +2!���0��9��^�ٕUݾ֖��g���TU �b
Ĉ�D�D@ �]���'�M[��hr��]�U��7IR�줾Z�,EDA��S)V
�RG�HA|�;wFR{�Qͩ��~܈���%a��[���9j�k!C�0�mwDj��7�ޥ�]t��p�a�^�LIɓl%):��W����Jw3oYD�ѷi��r�	�C��/:eϾ�|#��{0�#
��r�u��V���6�����|��ի�^ј�`x�f�R]϶�B�]��j="b3���9t�L��r��YF*\W=[�?e��:�_Z�%�E�Mt����D/*�j L�ڠ�G�s��VEr�;p�S�ݎ!B   �>��f�SY����3���I�F�����\�/�I���K��uf��hqza�e�Im�Ȋ���L�F�E�I��J�c��`UL.��!�U��]��9N���fU	���c	/���=8�h�f�RW��b�C��"}�V���!�xF��iz�zɐ` 7R���JL��
�֩Uu��9;˭�ʑ=���i����%7���Ӏ����*C����'�$����?+ ����e꽻����S�c"*�X��`�1�t�3�+w����ϭ��fk�E���A��=q���4�3��څȶ4�&�Y���i�:�O�U����͗���*.wf���쁶��n�2|=)��3��ԕ(7�K�}�|���1$Y�&�z���j�s�mU+���[Cx�H����R:��ȓm��A��nFEr9����EF2+�+\�����܍�/��#�ő�\p^�*i�fI��,<46�A+;Y.n�A��Ǖ>}mcz�}�YMg;z��BC�V�!���U�ü���ܗ�n˰ð���*!F�zw.��R��p��z9�9�[A��4Yq��n�S[5|kv�  s,m���� icl)�Hs ���[x)�̞(�J�	EZ�}>��ƥ�Q9�QO�
ڹ�Li���]�<�d��ʭ]?#��P�/��fg����]�Ț��U��w|� n���rw]������Н��8"�oiY,�i|�.J���?f��T@c"��""�)U��1�� R�]w߽��5��_�l�77��S/�����k
fV��0�f���q����0�GF��_*�U4vB�en�ΚDh�[]ROCz�O2�v���;�K[n�����;O=ÏA�.-ϖ��(Rn�n7{C�q/�����>�Y7f�e��4�wm]U���~w���.q�m�����<*P�f��3c�Gd*`�L�
���/������o�����ߍr}es#ҧ����]���M��)$ 2e4�L�{w�5-�
P�n'8;����:���A2;�q�8��N���aU����O����Q��S7�HL�Mn�Mk�#QT,Q#�8�xsʿL�'(�*�`��PX4#�"ŀ�X����)"g~2��'����3���M���ܨf�˓*+�wh�Z�E׏s	/���7�h�ޘ`������b��@7���h����>��h�Ԧ1E��,b���n�d�I$�� O^���pi�~cWL�[��V��4m�i�~v:�j7�(��K���'Q�\|��U�DT��D" Y ��"���QC�W޷��Շze7i���[uC�!�~��*HB]��d�e.o���r"E�3$����Z禍�[<Fj)IL�}�.��k�.P�R� �73�Ҍ�uQ�s7T�����ћ�<�>Λ�`Q�ڴE��Ӕ �IU�Mx}�_P��i��zb������G�)�ز���D�<�|硺�d�e�����nvܻnj偞��S��_��Ӟ�=n�0  �W��$������g;����L��2�q#����}�jaY	}��\o�7����	 ��o�}3�{�3��Mհ�2������H(%��̉ݪ�O�F���q��A��OXOɻ�3�M��JV(x(����)�f�
���[���B�|�]��k��3ʨ���ԏ\�� ��!n��l�Zb�'��$u�;O[f7Q�G�~�F���:*��'�Y\��\Uӆ�sfS�t�N+����g�ۛ\y,�sz	9AF�����q�\�w��J=Ѭ�^od�1�$H��$i**mr��Zo/$sY��;��suN]������?1!\�8�n��տ�w}�s�z����b��H�BEH��$��9������V*E�dQ@UB,R	?or�^���U��[�vF��"&�|�(��ԆR� ���I��؍"����t�펾vD�DL$h���,�[��n�2�t���S��Ñ��o@�n�T&<>=�w��ZĦV��k}�-k�zc�-��5���bUeh��kp�l�����v/���[ݹ]Ͳ(t���l��[���c�b���ڇ��μ9���IF�W^��r,�@E(�H? {�L��>)���글�����5Z�Y8�+�0�26�-[Yl�z��N5���Þc͐�Ζ�"�@��N��+!�c2�f	�󕴶)�cR9��$	�{Kn�!I��"����{*b@�S�ZG��!��n��Q��OV��α5!$��C�%Һ	�u=���r��}��.���,RH������=�EF�&bֵ���um��D�Xp�'d�ئ+�X��:D��	�/�����^묻Vu�LSLõc[�G%1*w&/^D��Z#�SPj��s���:U|��Vq�acG9A�(��X�"0`��$ �A���
{\^V��>��Z6���`�LF L�e{n��u3p�
݊�_DI���z���;�L��CQ&lΤ����z�9�� ����#�!E��WU��H���I"���4���^9�� ��r/aԱ���P<�I|��6j�U��>WLB<Z��S�u���a>PQ�(J1�jWN�11IL�LoP
�Nr�W�=��]�ʵma�D���g��:��k�"�m���#Epב���AY,DYb~������~-�J��C7��n\�E5{/Dl��o�:����%����'��F�3�d-�;!��w��[�ݰ�~�ݛH;��;ѱ]����|�Ra�\�yZԮ|��*ڢ	�5-8����X/��|�a�QE-����G��]�u��T��b	-��.�.�����'���g�5 �vH
V5OT��G%1���Uj���]V�/���9^�(DU���VEPT@U R
AI�U�� ,�H,ϯ��Zb��l��U�<��J��3$�:�܏��7���X�eh����o�wz��=Oe�ݑl"�d��cs-�        6�2K�H$��T��� m��늪s1��q[�-k���zhEJ� �7� ��z%�%"xYwh��oD�L��ۺ1;�q!��[m�d)�L�uL5_�f����z�󎊉x�>e�Y��]�Y�&&s�ļ�5-ע�L�X�~H�����Ϋk�+e���[�i��L��BI���눅er\"d=� ގ��P�䈥�Z�qY#�j�"a���]r��;��v�E��dǢgL���LچU��1H� ����T��0H(`��}�>ֺR���|�v"}��k^��V���p��|��h�[P�+�ȼ��2wtK�R[cʞ�pl���oމ�f<�AU�qq��N��2��]�jn�B��m�RB�%�K��� �ķ�#�oDA �v6���{�Fw�y���C��rD������V�My4��q
���a�=��|�4d�8�[���Fs�ŷ[S � ]�ķn��{&%Sj2К��~�	�|�>$&��M�[]��ʮ�E$�"�Y��HA`BE��  OЮ��x��u�=X�E���5�^�ʚL�q�]b���(�/uXl�m���;j΄w;.��W%��P	z��hٚ��<��jg��6:�S�
�&J�lb�^���X"�>6h�\�V�=�YU�q㉊�k��&R*�MS��lJz"tD�h���iE�K.�t�^�B�}� ,.����o����xHD�!3�Ѭ��&1�]&�]a3���;��[ޚUUA������A��[�/Jܵ���H<{�y/Tq�<T~��(B^s7�� >c@�H �[+�/�CF�B�x�?%���6q�k����Fsy�D�-�v��;�lEJ\%����w֦�Q5��;{�y�l| T���p;��d*	ϒv�L&}r�"gt�#?����L$�����%����b��09��S;*a�W�S�SJ�zd�UYJr�ˉ�6���hY�>DTcwr��J�y+Iq��`��C���cg��7�#c�m��D�d�ATUc�E"��mΞި���\.��|� ����#��y�koq�~���[#V���FGJ9��
G��a':L���3	ɒ�$�,���'�S��I�ې�����P>�+H���i��C*$�+vb��ʁ��%${YVۮ�Z�c�&�נm�.�-��Q��k>��x*�
E,�`�KwY���87�+�
����*���E�EK@�֫�:��Wue]����b����:�J�A�w׷�4b�j���'�S�lͣ�;vtv���ݷ�<�0�y�V��1�]�i�[��A�N�M�
���h����.	UA@�9O[��ׂ>וww�#x�.��͊����o��U�����,���/+'�f�DR) h� �Af��ї5�c��������/:�b��k,crS�	{i����lh�M�OYh��kI;�f��<j%[xv�S�����K�[	:�s�Hr�w��y���n���k�faHl���hoUU�o��bJ15�,0HJ���蜻n) ��WMoTfz�H:Lw�������A���U��6��g�

M�Ġ�m�=��ڣj��D�R�4Ym�~I2I�9j�ps%�u��8�*�M�9Us���^�u5Z�zn�ɖٙe�/2�*�j�j��T!CCIwW-�)� !Le�n��C��.�6-��
*h�ʎ���#�����OQm�qC.��>�0�'Rx��K��q��/��I�59�U:�Ȥ\�A���A�K����s�nu@w���[�S�d��vգ}��#�=�W�����p��%���N�v��)	Q���F���{#+tԧ?-fT�HFO+�YR��H`��)���&%۬�H9�t�QׯVVjv�&�K��L���%F����-��Q�wO�+���WGB��'5ay��]�sCw՛�d]6���j��[¢BZ��r���kw��an:VX�TmVܸ�=2�e�ѕ��) 9���\֤�nGx6\��6�.�q�0%ݧE&�]��yi�-e��y�.�̓&ɋ��v��ҹ��P��:�1����=�{��ם���{�l�+th�5�P�Z���Z6z^)uw���>sAj�x*^Q�/Vv�[���:��<�e��XK爤~���qi����14 ������;ݴ��Ζ��_"+/5۰���[�. �J������9��e	dM�5�H�P�g ��|�l��Q�N�J���j�j�-�y3��[�{X�x��)$wVR�"8����7T2s&b���-'HD��s�7�<D�ydO*u�42o��q+k�[�+�]��zF0u���\i^�c��7�`��uuB]�M,���`�HZ�%�ncG{�޾�_8������Æ��1Xҗ[��z���r󹲷?ڤR;{��X�мש�<_dD"�$�g��h����7hT����hd�;��PC�F��*����Q�>���~�^`�&O��HX�q��
�����U�K:NJR��NnT���\���q��e�Z�K����S��rή�n�� ID�p��wPZ�|��IT���>#������m�M��ʥ<�(y�6�Co 7��!k�5��}dr�[���g̨��5�r\�p}��oN��p3���� ��)^�UX���I^���t�.+��S�U�<[�� B�� ���^��鸷q��<b �ɆAģ�3NgǴ��uf#���4�񎬙�kȣ=�A�2q�ak�D�����z����U@Q�b1E����x9[�=�F��Q���7{ƫTF)�$"�$�AFAP��dPRb��`����2����$��G%��(�C1��!,�W�X�z舋l�T^6^�� "�eZȆM�y�:1����q����������g~��k��5��sz��R�Y�p��
���������V��/5����h�!n�Sl=���ܕ��vҊ���Z\f�rO�0��~:���W�\b4*(�z�o|�}��;ϣ�sUv1ֶ;P�y�ìa�/%>�^j�{<)ʗ\�HR�3����\�{��1D6�!?�!���v�����-H�X�Dk��UK��4���Q/j饣y�q�M� �X�IH��~�g������)�σ�"2亜6a���𹣝Wn:��I�m!*_4�y�=S��$f0�зy�6��^��#5�(��k
D��TM��y�:Ҭ�y��8h�a{�f���=�:H=>��A�dA@�Ǔw��ܝ�I�-�V�6jLr���������5��Wl��LQ�`��i��y���F)�-�g���9��v�/:� w��7�|V1�a���C�T}Y����1F+E I!, �G������[0=�-t�9���֏K)�K��Y.��D!�a|�o��{�]o��]w�NS�{W2Xz�9��{t| �o,Ź��س��S7sS$� ��IIچ�z�+����bu�%=��*rhr�.5�j��(����P��u7����i�vh�u�L.B97v��K�$I��nD        8r�0�%$�{Y{wj7w���	��}���PR��\;]�A��C�`����fҙ��5����Zm�����1&>Dp��nD��( �B�؞�m`��ՙ�<��EU����9B�ګ�޾��r樭��c�4�������>^Ls��y�/"R�<J��^pc��I�<���s�y^G �#H������2Ze��R0�����AH{�ʵamGc�ݤ4��B�:6{�sRV2:�
Z��| nv�g�5�"�^��`���Ħ�E��'Uk8\�Վ��L̯��{U�E��jc2��Li��c��_4��#M�ʽ��6$ҟ����|��u�+`�U��@c$�q�0�]��c�TX ��
�*(�P	�O\�cVR�S�����f����|M�����kȠ ˖B�~H�\��)$5�yŚ�x)�F��Æ��Ź��j���8i�R��d�/|>;�ţ��}�����
�^�.D��@�E���W���$�����tf�jY��_M�dv�S@�i����;f4��R�N&����C7�R��{g_^���o��f;U5蝜H��o��f1K��`!g�w+���L}�ol*��Li�P��{��ئ�G��E"$P� �`�D`�كc��~Ζ�rz�7OlE�����Q�o^5��a��1�z��}�w9>��j�x�B�o��ں���V%+�چa�.�F����^��Rh���+V��'O/�m?�
�3�\Q�n�h���N��a�m�T�B�wV�r�v5o��m��1��21�,V1Ru-�0����LD2a�"5��&��뙈,U�,4_�H��{��aUg��v<k�/��*���5A���Q��W��d掅y^սn�j�a*?HY�7�i��;���ndp�59Wp#H�+7���}�=ߣ�&׮�e#����K�4���=,;}�?�;�_>�?]{
���p$�d��e�/�L�Y��^�%"�ޏ/��
co�f$*Z�p�GE��eK�ؙN]\��0�݄;6��rajx:&�NC@�#�1�I�;��a�2\i�\�Ĩ֛[����|8�A�x��}��
����T��y2�<�tB�*�X�5�?s<�ȸ�v��m�Y�V#���VRsہ\��kǑ��{��z��������E���R�O�,�d�m�Ŗ,dCP���`J��Y��j	��u;�u��)4;#O��H�C;�F�e�Y��j �:(j���k�*qr���WF������Q`Ȃ��! -������ڪ�b��DA��u�v�/��$wc'��Ro2��y���q�=���ž�`��DE��_w\7.�I���D��Q�8��ڨ�aɸ���.(��Wk�| <G>��6�yϤ��I�r�9/ �ujg���`<��ڻU�P:�����!��Yoqn�f���q��9�G�}�op�����b町+�Vc�	V^�#p<.���B%���uh�N���<�d��e�"/��vV���H��}r���~Ѻh����ϻ���B}	7@O�g���jHf{Z�y�N{vv:��¸Ո�L��g5e("��;1+�;1��~�b\�y�̌�ɒc`R��PZqڄ|K�O�1����u{� ��NWBx|=W��g#�8؉Y��ڨ�k������0J�!�bwd�+|��q�2���?	j�5��_[�{�w߯^��S�/X4
"(�1,���P@PD`������{T���tF"1$`H�PV,�X�y�~�G��W6K������c,2x݌�v���^=MA�h��k�<|_e��,��}+V�'���)�9m��S{W��%
�K�+�J���AJ��`��<EPB��\��u:�KH����=Q:W)�'嗝9�������A&	�w��ҡ�����ս>��D��omv��ay{z�H�F(�� �}E��'j��R+`�EAb,P�,X(�% �A"*�UDUUb�=5�"�mU��4��s�cvs5�	Y9���A��{�6�\RoA�ME��fb��W����e.S��� %J�@6��  �`  9	 �l���M� �Qw.">P�3K�t�^Z�z_#�w'yI��[��j�
��ރ���;��Fȼ\YHSl��·@oNk��[!��k�E�N������0VN���||��*{�@ЊÊz�g�����M��{1��\zΏtk��x�>�e�kj�2�V���X ��")`��('��-(T.*��nV�|<>�d�����^���~֯Y�gu���q�zx;�"��p���k\:#����|T��M��3����٤r/uzL@�YJ0*imu18jї���}��T�:�7�tOyb�KhJn��pRcܰ�J��m@�n���y��k��o��� �h&%�\��g�W�\N��m��|_��Ōmk�k���]��$���PG�s_}���c�����9j�`A!�b�9��X�}�}��p�v�rZ���e���1ȟe�
��\�'Z�9騇[{u�	H�����m�WKe�����냯.�x.���Py������<�?����2�d=�Dۜūkz�|t��5r�:/7���~��D��$SXf�,�j�o�b�����6�bMA8�����a,�G���s�-��o:�̖���TTl̵�s��^׬�U_,֚��S�C������ �ު���PV0VD`��@PX,���_߷�պ�{o�w�ƨpvCkJ�vOs[,�G��B��1���7z��^8�O��)d��ה%���lcI[�#)��`���3�C_RR5��f}
cx��Pmx����P��B��#X����&D�f�mʜS��t-��![aMGz~�B�o	������P�Gt~���b���[%ℾ�p���(�Ƌ���M�U*�I@H��)���Y����u�<�)�C�^ �aE�}��t�H�y!}WV`�tW��Z�v`�u�:+�_S��� O^������v��v�w|�,Rp�����v��q\ꦬ������o���mt�k�#�R�0�q)}��:��.!�\\�e������f<Cv��=W�5컼s����{?G�}�^�||�uuu�U���RN86f�A�7S�����;�-u�q���'gj&�:yݎ�ƭKȌS���s&�;�y}��U��ޭe9��Pb��E`���$P�"�H�H �H�{�<�V���z��o� e��Q"�$Ac/��P~}y��bw_�l�ǻ/�P�L��Vg����RՀC�<�ܘ�'�������i����0�/Tg,����w��z��z��
�3ǳ� ���x}��~�vx�П�J���F�w"�6Ax	���Y�W�G(J��ݶ����*�3�����.�^N͡:�Us�"�񴺬'�0b�1�Y|8z�i]�G��3��?s]0��8��Is<���U��8��~ى��ǯ^�+Gl��Ȃ�ӣ������*ؤ�P@�t�s���	�����G;��b0a�o6�d�wK��"j�O/QX4GA����%��ܣ��W���J���s�ڐ�Er��"< �@��P���O/E?�T�m�z�h{if���Y��b�G�BҹV���.�Ta��!RwNҼUK��w�`�q���uM5��4	��ʜ��?Zo?n���U�A��A���21�V0d$`��"���"
�#;��~}��|jߨ�/�x�j[X���Ao��`�*x߹�>�$r�X���wbb
�H���b֌Y:����}���D�需�����nb�l���I��P�Ic���3]h�t3�-�-K�Չ�ʶ�=s�g�u(�X��z��.�5rx��ᅩiݹ���i�IATh�R2�T���gO�28��zl/�6U�FP��.�	W���b�:U�� J��x�u��q�-g�]�o`/�u���F%�n�z��#�xc\�5�9i�^ |��W�	)b�@1r�ǐQ
��P}��5���1ٮ�<���I{v��!�[T���%fPg �nM�z	�����5�c�H��*wt�۫da�)�̓�.^�%����5�f˗�,*�`j����r�*�$V����vݻ��Y�k2����5��V��v֎�n��-&�}�lpH
�R黗������3.�&�Y�_,.��EN9��i���q���AA%��
LI�����F�i��X�7@��%$��m9%�Q̺Ț�?X�U�fԥO5�<ͤ�0g(��mq8�i�!����h����w^�o��+��N=ߔ�_!hJ���1]3t@���2�I��d ��W�4�n��g'+�3�z����c�Ź�{R$J�>[��ו�tcE���N����į��5ı�D�$��f`��g&0*͚��t}*���݊W�iK���nH�)�����i�Xuz��m��5|�ї]�Ӯ����6�@�B�%������J��4ܳ���[k��;ܡd��z�׎��z�~��5�� �f�i����i@#1�自�.�Rt��˩�'Ʈ\m���<�Hd��W:�.4��tT�Y*
�}�8CS�S�YǮt��:�eܻ0����!{n�s��/�Uo��Y�q�'�p,�hٴm�x�g:��ł��w�XH�z�J�<�NoXZ����g 7�3<w����s6�io/sn_'��i��m��n�w��Eɶ���%����\#�m��	S)mr�oH��;�w�4cV��;�S$\m+q����Z��خ��<O�Ru��q\��=}i��Qa͎�[wj�Q=7*��k�!I�3��}�uЙ�Av!��[��s�?�;��Y� �eM�z�8�&-��e�۾ԫ��Ӆ���o�tS�\S��9��X��x1��37f��[[ WS��-꫊�H�3�_vТB�VغT�`<#K��-2�MoU?WTN?c�%�P�x��ߨ����ѯe��m]��6��^��l�J�l�@�ϸ�g@��W���q��%��.�^ |���w+)n�X+� �r�ȹ\w
9�
���i3<*c'_X����nu���e�/���X�Ύk�q�v������I��ʿ��Һ���X��o]YZs]�T!�؟b�����u����p�Zčw4�\n����Wn�����*���!�G��ܺ{��I� � 	 C @���  Je�     ��l I  	` �`   m��`           6�H   �   	         RB���K	!��	 P0�I�-L��     S|»;��UҮ�nu���|eA5�1}�$`k�J�ӻ��Y��p��"�lJ��x~��}��]���:�e�|���2��[m��    m�� %˖�p�I(�����کyN  j�u�elӼ^�����dn�#sC����YEkU�|��c1��2#�<9�ى��[�{�0�t���=��Ē^�!�@dRA"H	b(F" ?a�Y��+`��T ��#U����E��7���ۧ�q��g�ܥDa��b�RiV�Fy��2{{q������=~OD�׮��k��;�m�K|�i�kl:'�{0��3�:�����|> �=>8t�k�.����o�6�C�a��`�Q���:a��n¹@m�.�+��+�@�x��{=����nЄ������ �ca\���AdR�?BGC�GO���,�:v��6���f��}�sZ�0�f�v��%{�����tN{�ў̙w@���?6��G��)}/h,�vD��Q�׆w�^x����f=����:�2��	���:���O*��$)H�E�@��V�7����%���%�e�w���3�T��Y5��n��V���uL���*����-j%����u(��.�;����k��}����>\}�D�����`��0�!��g�]j����A��!X�*0"�,��}�{3�i���M�y �
��X�(,������ֳ������"�a@3ł�������:{h����r�Q�W{� �m�m���kT�WK�ݓ�zz��F�.#f��`�}�U������G.�!�,{�jO{����O��n�� ���j���A��f�xB2�BZr��a`�:�+���W��Q݁z^����5��/�|>1����ݡA�s8�2Y?�۰W�K�T�F�����FŸ�t�5�I�p��齒;7�*�X�5M�kR�
���غi13���ʏX�<��K�zCy�y����*��U�͟�[���D���jх�<�E��\��
0^��.V��5�2�۪^���)���X��q�I�E� �
>��L{es|��]�\�pm��en��_\+����9+`�H]�+]Ek�n�>2�����y�u�gv����H��u�IZP�Vb梁�� � �F$ D�g� ��_շ�����n�Wu�mH�H�VDU�)���Y!���뫲�s������˘m[2��n�̴l�7
/o�F>���8�ߡ>���/bφ褍�53U�]��m%�R�|>q�Wf謁�D���3'��;О�Q��s:�:w�
�/�$�5���r��i�G��{���P�������rl�U�:�k7LN^s�^gvz��}ܭ�}�oZ�`(1b,���b`,��P>��H��lx���,��7}4se���뵫쌹���tOM��J��������M�ò��Z������1G��C�L��'�3���	��+� �mc� �k�w��1ʃ]���ƩA�Xn��C�6~f�ڤ�v��q�sаsލ:��:��D��Κ�GDU�'w/W[7��Ub��';�~ ;���т�ȫ"1E (� �E!�O��+��u��e��PB�����N�r0NE�ץ����|S����Վ9�,"����"�Vb/9�}�$%�����j���3s{��G�d�w�f��Y���DPgi��r�O�|WV�҈W����Cr�P��5k��qn��&j�ȮR2�"��,c!)�4�)`ު紡�Z_������-{}�L:���t���e�k�E�T�U���^��Y���<�B�l�?z�5S���6��m4�q$��6B�s��EsX��ͭ�q�}� N���Ґ9�MOj��q��3���e�,cX�ua�2օaw������˄v�T�=z��	��'��ji`&m�(l��\2�s^�������]s��
��x޷��כj^�6��&��MK�h�i�+۪֢
�!�qWE{hE!�[)P����=���0DU�,(�F
��aEFI&V���}�������.��{]�~�� ������^�k���y����e��@0��/����ߚ�#n����]�N`�d������P��o1u���X�}��KlK����+U�W1��m� BHI�m�       73-�T��ΝF��j��pK=�������N��Dk۴u�(ń0�"#���tT�z��iEIo!�̔��|>��u��[�'#�fz�Md]�5&r�!+-n��d�����p�yc<qSPƭ�_��`ǝz��Z�ǱNn��;R�zǭ]�].����O��t�k�~�"B"H�!$XQb�X��f���T%��zw!�u*i5�ͣ
��sj��+5�i�ڳ�-cR�7Z��5��uchC��M�مp�k}�#����kC�G����]uẑ_y�S�,]^L�}�ԋW^q�9�ak�b���;�Y�ԁ������<�ԍ]u��=��m���!m̵��b�ܸ��:�ts�u�TT��$��Je2S*@�*U4��E�����^�{������O�z�Ш�++b#bEI����"��1TX�TQ`�A��7��}���m���C]VJ�Ab��U�g:CGkv��R)i� D���	��Ŝ��`uV�^��w� �{���/��U��]=:������A>ˊ,�:\\ѧB��x��<�s�l�oDu��1�c�
>��������)��!���J���չ-��[�~����,pF�\�����Y]�ܥ{��K�����׷{�^�PcWb��Q��������h�s��$��A"��H�²�R��ɑ
ߍj����׉�^Ô�&��4�q�q�XĒ�9�lr��(7r���1�]�G�����4��Q��W{�gL�Vh.�}��z��G<�`_��!��;Z�m����}2ܭu�6]J�3�fIcy�\�ߎ4 ח�Y;j`z�wb���ն�$�qR�t�F,��X�u�-�`1�A&O_�p�cUQ�@b�(##0 �*��
A`1?~���w�r�W��}�g���g�-aᣞ�T��#*�4X��	S����1]�+�c�P�x�)#�@�B=W����Ϩ�W���6��`,P�]`�n�Ir�v��0B��9S���f[[�:����]��]��\/e�u5�e���U�V�K���t��u|��Q��\��[k��|�r9`�1ɒÊs�d.O�H$n,��"�Fg>s��*��5I�}Ýa������J�Y����=��j����g[gt�}�G�dwP��n����z�a��膭�h[��MX)��0_�N��(Xo���P#�6j�pPrV�_{��dy-�qpʟ��?Cn�m��&���R�]F�17�3��r=�2�(�����
��(�&;Q�<�Q���M�xjJ&F�}m��_S]w�
f-���kb�@��
�U��'�b$��Yy&�e�+��?^�TTU@A"��Ub�����7_g���{<m���F_+�|0�"�dc (H��C�������&��~�c3k�r������3�l�*&̻�U�m<U�I��B;�Dz)�2�����v-�Ѻ��P6kzu��|priB��C�/i_}�����d����|��뻽_���aV�ǦU��L�sxQ���eht���+kJ˰�or�Z�����s���������(�5X������!���;��1m���l'����Y#��3-^3}�D��9ws�l�az��ߍL��NbHW��'Ve��.��?|�o����bA#,���߼��S�T�*�Cn*D53�Gt J�cy\�Q��1f�#t����k��U�tzI�n�z�%sx�I�"Cs�k�I�hfS���f"�w2��NDۢ$��#�ɬ��J<�'X����7�Pt��PxO.[f��v��qq��m���gB�,��6.��������)�5���&��u����o��^?x��(1B"ȃD�Y ��{�O����u����w�h�a�1�`�A"D���?�v�`b�� ��pH#�aێ������^1Yԗs����Z��ע��^����5:+ghtYR�*�����}����6;7�eD�ț��4.5�5q�PˎT���Qf��5��_Up�=��\��l��כ���C(��K-a���cj�;���o'k�)G��c�٘��:.�Ⴆ�\���FܩS-$L�m�  �`  I,r� I���(�]�aLD@p�6��gG���Q��C?z�?�5Y�-��[�3�l�{�hOw��=����Y��"C}��������-N�ǂ�J)}��,a���k�ݝ�Y�d	%�#. A�D�)�ku�j��~�fG��� �)y����\:ʕ3],� � +b���}�c�؇#�5[j�,�m�އ�v�TxԤ���������Q���+K�6���;y�����.QS��퀡F��k-q�]���ϫ�^N��!+G��,��EQY�EFA`���N�܂ק<"�b�K<��r�ܶ�+��Kiw\�-���	����}�l=Vv���v�s�"��֝��˨xf	�Qr�����ם i":�gn�B�"�� '�����,>��r'�Z
�U��b����h��U��{c���S�#�D��T���V��	-���I�z���}���_;^��\�s9�m�s����듩)ݑ��eV�+�l޴�s�v�0�&Q}�ܝC��ͮW	��]ܪ�6&�@Wo;��]ּ3�.Ǖo�ۻ^o��D"��� A���x �4���+o"�Tz��=S���sV��E�_K�I�1σ�y&hD��Q��=��K��ע�����竍^4y'��)��#��+j�Eͦb���|goٯ�f���
С�BW0/5\{F�u���#Pʻ���p��Gma/VO{��X�V՘q���azc�=�7v�}|}�kڽt�TdV"��b��`���~��{�߶w��3�L�D��2E�Ns����GkiE�_��&{=��������ݬ�  �N��R�T�w�1'�l#���u��c�
(�SgU�;�R�<Ϸ�Z�3tveM[Wb�]z�ٴ���x|C'��-�����[N3�*�iqxjӞ�&�1ZaN��A%�h�k%w��K�ԼV��;���k5�(9&{�����7P���@���쁷$<!�j�^�O��E�{�P�m^��W�պ�U���`F�"$�;���Wi�z����i�,�����(��g?��FH�;�R˯����Ʃ��D�뽼�(!�� �4p�r'ݽu�M
P�v�u,p�Un�*��}�Đ��}���֎^�p65)���� ��F2������C�O��r����\
:�kTI�³��>�XЃa�%:���-�\D��!x~���K��n��JP��mc��rɦ�QB�"��R�mu���7v�t��Y�e`���"�>N��ă4�J7A�J�8�oIi�k&0�p�+=P8ضM蠉"�
�V,�i����
_�Q4q�U��u������ɚ�FK�{�Q��2z��b�e�"�xvlO�+���&^����D�2��њ�;�uRKiue]�^����S��	�I)ǁ����f�1�Ң�dhp��WV#q*-�h*s��-,��{��][ʤ�jZI.1m+�~$��S�~�̡ʼJʶRu��"�Z��e�*������A7u��	���pr$@�D}t�2f>����>e���v�Z�a��.�,��ZGYR���OY�S���b�r�ħ�����qR:T�oUfBWѯni(}�:����;c�����@�:��o��ʩ�>p�y��j�$�K�!((��dp��ʷj"��3H@
]_%ҭ�}�n���Ԕ�Q׋%ù�S���R��f�^GG�V��T�zy˵�y'<T����}��TKeW7�����9O��Ga�Ȗ����g7��{S^_���x���Ѣ+�꽻q��Lי�m���&B�Ϊ2�-td��V�ޮ��u+"�8�#��Rn�ʞ�&��qsT�Ŏ�!�F�
����wj��] ڤ��Ѕ=����ʹ�[��Ă�3�wY����r��ƶ�]�G+s�\Y��Z:�t�r�U7������"`�v�ގ��*�Ac3B޹|;\�ڍ��#��F�,��c���tO"�z�h����J'}�dETu;�팶�7F�QM�oFMi*�P��Oe)e�8ﲎP썜ʌם����v"ΗEvR�L��0�'+z��Wc��+6i���A���z;]i=��!�۝k�Ȇ�Ӳ���W�2v=�.��!H�z[��$���[�
�I���Ä�Y����A�JwGˑQ�b��pt%Եf���ӄ�l<�5�,ZMh��S�no+��HҘr�y�;�q��3PL	ڜ��nT;Ƶu�ޝ���܈C�]W�����K#�y��zM��.l%�i�2cu����j�lɚ����SvpBc�s5�f;�p�	5��r�;_�,���h_�;��X��1�8��������Gt��H��-ى7���$�=��p[��i��e�/s��m�W����*�!�8�s�uo����:<I��u�R����c��yo	m���9*'���b��Yoy}O�¦�4��}��s1p��Vz�{?]u�Ub��+��?~ {u�O�v�'�V�Y��/���]�d_�a�,�3�Lh�68���)y�0]Ow���2�N���:f���S4���0��l_���W���^W�欤����5�K=Q
�������=w�Ik&5����q�O��OSq眶�!�F�C���̩��Xi��kJ����>����^lY>n�FE�9�%�s,w���j��oz�{�qٝ��m�F���w͛5omc|���E�/�9��7Iʴ����&��S���R�LZ��z�̈́㤛V-�=�t�}.`�������gl�Nrjx������]%(ryȳ4����$�� K%H=��cҋ�!Q>���E�]��q�M*��Rh^�wk��פֿ"��>T����y�|�[EE�o4�h���ga�2�(��j2V����=��쁰f�h�*1c`�)dTdb�H��H�#�����\�m��&����TT �����L�8R>+�. GE��h˗���Pfj儶X��V�^����ן�c*p΢
C���uaq�%m�{;e�І�H�ĵ���{��V�V/XTx��)�+�l'\(�s����:\{�+�V��4�.��=�����G�^gd���t��m7.��u���g�|*���j����~���IQD�
��5��m��꯹�����w��?��!�M"l����{�w�i�>�������>���,"�d�H�}�=�׍�!w>����3e��p۽Z]��rW{6�9�Cz��et��ʚ�r1c}�/ 3�p����\���.���  �� l �  �� ��R��H�ʹeޥ���n�bӢ+�,�W���&"c"��K%Z����XGH�U0u��l߇�-��ƎV���$j
�W��D�:҅�"�W�j�a5����Z��uǐ��!}�Qg��;�aR�E
ʲѨ����ATF���@��$PY#=��W����;�>��]���ߝ?4}�/��#^�豊H�G��~m�P���y�B�.�7+zgg��d�&�Us���Ⱦi���ly��_��5������xQ|XY��d���}�#��Ğ�TyA���Ǐ����(|J��z��g���[����7M�Gv�oWB��[a[�٢2É"�;�X7�� �5p���j���ifHs�D�!j��~���ܹ���(}!(�� �r�L�)5+��wt��Mn';薖cD<���־
pv�;re�p���^�C��.���1$4-��ocKwP.|> }"��c�O*]��$��u�)#	Ҹ��X�I4&;��3�&�Oqkئ�6s	���C`tBJ�+a+��ٶq�.u9���Ӷ�h��y�]�{m[��^_�Fy�ͨ���M
�Rkh�l���{���Z�5�ׁvC��yn#�CQ��:�̋:j���\���B* ���|>�~s�մ~��Zzn�<�E�Ƞ���d"0c��}��]w^��{wX���[Gy�z���Co]պ�P�~Οl��Md�����}q��nsK���*�V� �	Vڼ����]Ot�u�|�l7�#���FY��|��$�-��$�u�ۓ5D�����/=��?��6T��ɽH8��c��E�T�T�/��O��LP�ǳxgc/R���F�C���>�y ���d���d'��}Ϳj��?\/�zC'���+�]�.��2cd=�����R�'Ã:�'83I��|,��%�=�L��2��)~j��<.��bL��c%��� ;3�kԴ}�d"��&}�w=˽�Z��ι^9ǝ���5���u�{��V.���WF�nC��8����{�	��ilj��r�m����Ē��iG���XV����N=5
��;~<ͅ��}��w�=�M���8]L��L��]g�ӧ�M�2�/�!�������Q��U�
�`��7ߊ�W��� �>Q`�#"0d�2#$b�* 2A~�~ �wc��#m�5�«�֖�[���#^���1���1�Ȯ��89^.�o�R�k)��"E(
g�glt�+�Je��&}��8(٪�9����ﻪ���7�+2~&��}b�Ot<�陨jb[I�!��'<6}xTX�F;���ہ9J�1q��TԞ�1�ZKK�k�D�v	�w�q֣�0�dPTb$�:~����~�`��2��(ŰN79�]qq��UHa��D�)>X���'�o��3���ioû�/�]�Lm��b��I���_s]N�n�L�q=7X7�zk�ᵕ�| z	^�~RW��6��x��)�����M{,��8����) P���x��	6V_��Jd&�wg@�c�;_v���e��N ���͞��`�N�<ޠQ���U�`4�n�.45��_+�!��=k}#���
_�������z���]:��:���X��I"� �UE�@B���#g��X4b��țD9�����B*"�cTb"�#F��� ��I��u3v����{5R�N�y�!�
	mW)'f��ʶ&�f�nn��+�A��f9�__����LaL�b$*1��j�d��ni��{��鱗Y�����v��c��U��s��4Y8����چ�ƯtYr+`Y>�x��z㧭�Aˌ5@�omMk�Q��%�Ձ�����Ŵ�H�Q!���, 1~Ph�{ޜ�o1pĈ�y�L5D���Ԛó�v5D�3�E�h����J|ؕFy)A�[K�c,�Ǖ�i�n�{�����1�Wp�>y��|.�j��~�Tڥݓuz�m�\T����}�x;��t�竭���u���i�8��{����\�^��o�k}V��Z�����7o�5\9�lᛚ�S4^�x�*�(�>�t�Tb�ʀ����_{�wA$"Hm���       ̇ĩi<�-F}�U3bM�l�L��f�2���&1tQʝ�s2���ƣ� ���v�����F""�c#UE�)�,"��������޵�ֻ(�{u1v�F�zר�K���ô s��r;i]�l/8�4�W�~������|&t�c�k�R�G�❷sٵo!Q�v�d�U�y*�A#�a�����N�J[Ւ,���]�`�\�-*�<P�N壝�ܙW��1�N�T���2[���^%���v z^ ��QR, ��Qe~���K]��$��Dx_�.Y��j�c�5rk2v9|������Y��u_�2�Ա���;A9t{��j5:��&��-z�8�y@7��uL�L����6ldE�;l��/��l��t��֙�g��N��Lv2Ww!GHL�tE|V����ؽ^���£
͸�Ff 37Oa~��Y߫\�_Oj�-�mM�YA"�U 0X�(���OX��)g��H8�;�xYM��~��nF(n�G�h�υ�x��͜)jD*���)蹔�����r��^��v�~u���'КcB#	�]�����eοj�S'-FD(����v��6�]啡^Ľ��]3���fO)/U����|V>[���a|�-՝욅/}��O��*3v��\��G��z:r����w'����Z~�&��|��1�:'�ۣ菗�w����KE�b����6�1��3�<c6}��}_�L��=�_���t�D���1+R6ө6�v?��c�޹��wŅ�t�f8�=��n�p!�����k&�#i�nN��>��F����x��{j�l`���p9�| y><�;��Ӗ�����w��U��Aoֲ�4'�p�>C������/AkPX�����&��4n�v�} ��F*�U���r����9����wG��ܣ]ª��v�O�$�AH�P�J� ����_��|}T���~����H
B��߾�������ߟi��V#�CJ}ۧ9�S���l��=�jT�9gT��a�[ĲG)/zp�4ȣ�t���b��Y�e�Ӗ��/X��3�������x������A��J�����N��r�i׵��WK�ϱ=q,�K��ʅ��	:tr����1�1#Ӿ�NkEP�ǫ�4�s�e7|�gR�������'�|w��B��~��S�+�L�/�:ܰɩ�X�5X���s˺����ޏ1���7@���W�(�x��(��� ����E�W�%2��'��8�G���-
/��M��:U�g6���]L��Ʒ֢���y2l�����m�;�8���_�L�W(���Vh�c��k�VlI�O�Q�]�32i=�_[7�@��Q�
�]T��M�҆���Qy�u�^+N:�7��Ur'RS9�Cx2Y�{<KT��c|V����?x ���$V@FB"�PT���&}[��"��R2Ȍ��P?|	����WI�i<��*]�� �6x=¶��.u�;��;�߂���
?|>����,��懳Ţ��Ś3j'K���5�R�Uٗ3x�I������ɥ=�*�"y�+�z�V-�tb�W�yM����Qwo�6�,�2�\��P����c{`J�U�m�[UO�}��PkWj�ق�V
}��n�M.D}�)7=f�ut�]���x�q�*ӊl����U��H�פ�Ɯ��F�3<�U.���M��+�w�n�����W�ns�[��DT��c'ރatSF<��N����w>�躠2��c��p����J��̥��˿;S��P6�'�=�O��f����n@S�k���g}�����}r�'���H{�)�$�#|���sM�Ll@֨ơj:g�+#��Ū�)��~��U�7�V\�� �F10k��	����� P��5]��b(�F"$DUP�����g>�w��I'�_����,[Л3\��J�lI:�X�����95����-ɮS˫�`�TYVI��(Hv�7�S���,���t����L��'��C%c"�IE<�_�q��g\���ٷ�.Ժ���"f�7ct�[�I�h-��UBFg;S�߈�t�u�t�Y�ݒK�w��Ht�R��V��Ԩ37b2�A�zi>t��f�o�^[�9��{��,���se2��r�ڍ#L�ʔ+n_IU�Юp� l<�k4�&y�p�*v��W���Z4m6�"{�kvoMoY�2l�j��5Lr�kN�h�NYH�U��wueS(1�d4�����W�1{�
�β<��Y�Dr��؞�6������͉�c����6n�NA�ê˷
f�\�絫3��J�N(�N��4y׼�m��;#�>[�nu9,�4x
ƲPqPO-�б�Es[H�|���.;(2�9��'���Ɠ驚�+�����q�òE��u���Tu)e�Ζtq��뼭{^�h����|�%a��2�RNPQ��^9X�S���R$� �n՜
�����D��  �/L��wn���l��$R�Ŕ�FR^�7�5r����2�Qb��$A>kፆR��ll�n��	�	��h�m�U`��6�{��Z1�k-�FݢcBLe��?��V�u�(���yݹ�K�v^s�lʾ�\7{d���]m���k/��n��=�QW�1�p����ZG8����vn�wD�'�=��1pK���ۥۺ�omO�P��̒�o�ź�Tt^[ڰ ��)瓡J](��ޱ����F���B���ڭS�J�ɓ���;��eڜwvTK��ه(�e��~��G��~����s8WRM�.����t�N�/2%\�O�������"]D�o�ɲ���[�����y ���x,gw`�p��s�&�᭍����t�2���8�P���5�;x�0"Ŧ��\[n�6��XOB+Wq%�ɸ4)B��8Ete'8����|����lm���D�NTX��鷗���^���`ɏ ��]�����Z48�������V�-f�S2�@p�mvnܧ2ހ��r��V^���E�8IQ���
f�7�jU5a%[-=�Ǹ�N��i��§A��'e�P�q9�����uw¦��M�{������6��d��P!�y+� �j���j�����\p��u�Qfth�p�/sDm=��s�OaBDaWC���*6⒙ٛ���k�S��C���0V�܉�j(��S�������$�gr{P��W܎hCm�6��@�     �lB m��2��       i0@  6$ @         �           m���lI                  H�C��JQ. $�m)�D�P��  7�  ��)V��x*l��".&R@�p�m�[e�r�{���5�D��B��̙�r.I��M��U1t�o+���� 6Ɔ�   I   5.F�8�%535N/2�weQ-P ���S^dh�e�ζޤ�?��}�c�V�>��^z'�<{��={Q�E�,i�r�l�M�R�s���

���g�1������]I�o.���e�k��7U���O��ETA�F0b�����|��3��s�~0�V���5�v4�-��5��y�e.e�1�,�f��5,�26nқ?Q�^7So�:,B9��)J�u�g�,� �<1�2DO;�&4x}�Ј�&}��ӸT����Ҕ0�S(Ei�7�5?
��;����T)��v�&V�Y���ǲ��Y��1Q�m��~��{�[6�^'�M���ʇ��Q@�$�,�$���/>|e[�3屫���k�[�O�M� ��g3����2�#w^��Fl˵���vT�/V~=4�:�1�ٶ5j�z/�,.VV��`Iz\i��6FG� ������>G�}5��&���5�rQ�MU-S,������[����<�8y휜�ҕ��T�ӭ���z�[f3N�qwu%��.s�i_��mC���(?q��&��	e��$2�n$��;�5ֆ<z���tv�+@����D�<	k3�Ebt���}]{ܛ��ٗ��d�`�#� �u��I|k���}��h��]T��c6_R�@�{r�Uڥ	�)�*�ﯪ|��s�%�w�U��	���}�ۧK�c�\�Za=3�H���OE&j�e�Riϫ��Μ;�w�Ҥv�"�QQ%�$��n&:��h�~��ro�T��N<�ފ�a2�D!uUZ(��F#8Ƙ�a���a�`#��,P)�Bk����\�
�ł�b@A����H�6�z�.|��i&�4��X���dV���D��9����4+���r�<��u���p�iA��KM;���,�ڇ@��q�Ff���|}���oBѓ�<��Fiv}��h���9��"�@RI5ts7�V�{����vs�l�
qA�Z�S�B��9&�3��4��v��ft�7l�ؓ}'lU8vKE9�poQ�V�GxV�[�&��mF;i���G=��yZWA��6=�W�_]<ʯ_�@T"�T	��1��W�@�֚hu�s�w+l'k�{bA]�����M����#�B�����O.u#4i�ťep�	�Sr՚��Q���}��������S>�ݽ����r:��`&�S��&۪���3.u#�mW;AQ��S�3g���w��ų�U����it����0���Յ�]ݙZl�TbB�U��F*��("
DH#R#"2,TAs�����5��}���� =��>�\��]j��Ly�鎛���n��O�,ջ������rl�=��q1f�	5�|��w�+z�K��>(j<�"����:�#�Z�_gNLDL�S�gU����T������H� ��NY�1-��Z~:�3�H�� }��ʋ��ؚ�~�S����e��{�z�G�k����'�����|�6%fS�x����C�άדBwt�dr���K0�A��x]���Ǔ��z��sw���o	�%9��`�"�Y$P"���}�l���g�����}�2��O_B���K1"2���	V��e� �\ǳ3wo�Kj��	S�|��W���ƆдǊ\^N��3K&
���iD��{Ve��F̩�~��wlW}=R9����Ǉt�]OV�t��+UN\	p��s#m�S�eL����#��4��ވ¦KU��/���E�tnϠ�VOl��u�wO|Q��~������R"
�A Fc )?BL�����KG7^v~ײV�"���X*���EH����5��{u�ɷ��w�{�#50�H���^̏�pz6γ���n�[r��^?L����kf�?+�6qK�沽���{���}</�F�
Y
c	��[���n;�2b�jb�*��
���]�����A}�f|���:إ-�l�S-����0�a`�wT�4Ң�b��Ȫ��"�b"�DU���2�P��O����A�^>�B�>��U]��Gm�v��:۹��݄���Գm���*rf�՗V�������9qlө/FY�V��D��Je �M�   ���"%J��B��-5�z����	f]Uj�y�k���<�1�DC�K!z��O���K��R�|w��\(��۹��3u�N̼:��kz}JA����>�
���^X����ZN2���VL��o�NS��E&ub���#� ��/%�^��܊4*�Nd�,D����P���0��*�َW�=k���y��PP�>��S�TS����UJ�Q��J�DR�+�}½� {] ���$� ���M��R ��c%{�կ�}�o��W���v���@�"��#j��n�.��]�D1��=�/�"�܊�
�^��$�$ ���w�:b���"�X��)\��������}ˌ�+�h�|qL�'�)dG���{��� &�͝ʕ,"�v��@/��̒5}6��Sq*�in\e��
��E���fۃ�~}���K������A�����~}$I@�$4� ^���b絓�C}k���c,�q��a��C%�[y�"�/D�j%#�s�T��P���,p�;��<��{���'_�[S��>�
�!�׶�l�9օ~�dz~���������|�	�.6�g!L�#��>k���
M]��J�_�|�2P�i{��x�_�d���<��,�ڰ^��^�Yy� ��� �W���4�a��xZ���mn����r�Z����2
�EQI �
H�����ʽw���Z�!���0b�"$@AdbH(|	 ʕ�
m3�Ն�Qj�!�5�.��)>:*]-9;]��W�w���}�=�3�K�)3$b0���ы�ϼ�	\DC;�#kO{�v/��=���=����#���e�}��>������G���>������b�aV^W%���bϷ�|'�������ۇQ��&j��Ĝ��v�g^u���==�"0b����"�lg�����������Q�&dH�E7��h��%E��"�����}�  �Y�#ޯڃ���gL3+��ݢ�D�P=ח�_I}�
F�v.FК�
n�'7~W�K=�nN���$��R�q��[v��K��j������nLb���V��15�2��BWh�ލDf��A�#���|����{ɓ��e����њ��%/����Be���T�}^9�,P�i�w��!����mdX"g\�|_W�� ~�G�iv����l�&�A�Mg4_߾��~�ڬ���W��,QAF  ��H�(0a ]Ne�ݛQa��� L<�;���c��1���ߢ_iq��cy�퍊����/��9
���c�Eu��\����=xig� ��E-j�;M�qXm��|�4>'&%�L��ڍ���Ʌ)ƭ1G����
/�w�T}fj-�}6s��|Ui��F�]E� R��KU�G�U�KQ��D�|	��|5E���n��ά�DRB������(�U�N榀�*�p!	orފCMʎ����%D��ڸH�m��>���G�|Ha�z� �_L�K�R���v�'R.��1L�=�H��wc�=!nmf���:�-eG���v�Cgv.f}f��	Ky
�ek�;�l�!ĶЪi��lO���a��=����srnu��Ƹq����UM��9�4p���M#K�w�u���h��}�@���<�+m���K�i���Jdq�Vt��F�0}�����x'՜���@F" �"�0HF2 ��3�O�AUX��2
*��=�W��k����|����t��%�FR'M}"��Gj}j$�S�m��.����A�i���|��\�5<2.��:���\*���)�r�L�V�MO� �ez���O;c��˵Z�־�C������]�����VF�/�Ƈ׽�d���z6���%�����~��ս6��o��-�զ���� �X$ ّ���َS�HČ`�**�㒛�n��9�f�ٹ�"�t{%v�4��Dσ��V���Z��.rf��j7�!��o����>8f��BOq�ߡ<��EM���q}Y�V;�����D�b��;����`P�]����S42ڍ��ec�u�fή�����nؚL�$  �`  jZ  �ԹM˒ZCW���nBC��EJ�q���-d�z��>/�L��ք$�����\co�u�7��X�ܩ:�x[u~َ�� �!c�uT��tk�B��?~	����T`,R)�W\�w������v&`�VB(EH�B��G��
�sC}3��ϝҸS*:^�[�G$���R�����P&�w����?!� q��w�e�b��dl�5�|1��v�e����L8Pz�<۟1��RK�d�C�Z歗�ϡ��2�]^�$�q�	��=v�^�^X�.��9G���� J^QKݶ��(PS۵�]���D�3�$�}��������� F��؝9�6}q�,�� ��.z'�ֽ/�U�槯�"�l @�S��i��؍�seOy�1� �^���
���3�0�n�U���{�)��}�����PE{��2E|�`�t�[���ςJdY RK�Y+�������w��9A�d�:���fR���n�:Y�-0�\3obv4UG�1�A{0&ޫ�ݠS�ս��O$��𻕖���+����W�F�zTJ��y�]h��<u���*>kf�Z�l]��~޿sRI�(S�w*x�_��m����b�R"��T���Y�E���M��ퟮ����F�����lQ�G1�l�6&�����`/���c�Ө�4�PB��#�F�R��;�- �y@�lk��}�W-ͻr�����P�Ӝ�E�Q+�םz:��(�}EH�]͙��Q.��cuc�ƚ��[*�r�=�����EP�wIY\�Kl�BC|yk�:��������;�b�ܿxUAٷ����]�dmj��vN^����zVX_q��Ě�@��Pl�XH!�WV���y�]�I���:��ˆF�^ }c�ղ���I'ު�a7E��t�I͛TqT��qhLbԒt�����yQ|O�%(���r�BMPz)ӥW�YVV Y�DFr��j��Pr8�n�Y�a3�8\�U���h��T,PjQŖa7�O���M""ʮ����E�̉�*6VIV��a�X�F�P�e^��R���}�j��T�n]L�N��JR�hE�	�%�לi��"���E����p�3�O	�8��]-���SI nS��,J�w���W
:�Sy�_�u:��wk������R��%�44HP��9����\n�xr���;��k��,͚VO��2�uae_*үY8G�n�wu��|$���6r�`DY@ ���Z��&�h�t���X�-y�TR�iE�k��*���
��ְ�x��ק0㗠�h�}��� Yi���y$��\�)������LՆ�D�V���uyy������S�ۦh^�"�3��Ō�~ˣ����9^��kxt��2�o�����s�
UU0����]9�vs�b��XP���+̴�J+���\JJ۫�[��{:1��Q]޿�Ԕ�T���K
6uØ�W��u�1��k��8L���!#��{�6�Zݩ�r����^jU¢�8�ΡljV��w�5��{�}�b�� J��rfP���U�5����2rV�a[ۚͤ�J�յM� �N-��Ժ�.���*�v���G�99����%$2�8Vq���a�Il�@q�-��&��+Գ$T��۫S4N����.˞#b�oA��i��o�,�(�a�ٱ�<�M����������W����4o���i��w��B�7����V��vD����IKj�L����&�DGQ�f�o0L�vs`�
�J�6�S�;�,0�s�,v��[�O6�=ᕊ�hԖ]YDї�[p���5��:���V�Y�Ve����]���u�{.��ȍ���'�*��p�9ۓDP��h�V��Uy�/'dݵ��3�{m1�Ô���I����B{/r���2ͦ�;k8�٫��/��0Z�/A#�N����;Sd�}�P�F�����^���%���un�X۬B��&�^눧���g2P�꽦��0���W��i7���K�h��f�49�4��������M�>�Jp7e��oqm5ҦDn���I�`'0���l� ��i��N5F嬬siD]^k��ٴw[�
���� ���C�\з�Z��+S�R[����{��˻=����ٮ˾t]�AP<�v�Ի�C�c!=�N�ω ��i�.�0�w\D���(a7p�}o ~��
���ױY�X"��)U�	�}|Q��}�]��W&�O'�يrH�^o�6ԝ�}9[v��ҷ�|�<�ձ틷���!���c�]ⷮ�=-!Փ�swޓ���Y�O�������=��{��5u��Z��y)C���k2n�6�8�D�]�`����Z�t�Jvx���g��y���)A��d�ne��湇�������[���R,	"$�F@DX-:��G����wFf�������ft�zSR^yI�.�Jb���L�&�NL���ʃ��o1˦�P�#���LE8t��+I��"A�jVB��摹qx|>r����>��ˊ��!}�%ڿFډ̩��0V�������nv�������^!������L��vgɘ�L1�i�l^�ة�Oď�?1�QUX����`��G��A ���Q*%�	8\�x�[����
H�5�Y��+�;�)oz���خ�4��	�}�d��މ�{�Ik�n@�=y�<��U}�W� (P�# �A`,��~�}\/�0�=Wf[�?�5���[�9��v|f�8c��������U-�����C�?P���K���s���I%I�@{�Ԡ����ѩ��:u�:��|>�x�F��ԅy@�6����R���	�*ٗ�/YZ]Ȯe��zW���A@y��O���R�T��/a���q�[S�9$�rv�zP�'g� � q�߳���X�5\'@���ȗ�qqm�9��'�o2�����_{��u���M�ز-wF���Z�\�!�.������#�I=r�7�x2'q+�o��7-���+�qB1�7$��Y�mA^��uD��tz���ވl��-�=�?{�C�
���~~1:Z;�n�=�}r�,=��Fvr:�=E�U6l<f�����8�ﮍѧo|���
#�����,H�TUb��"(D`� � �Q�#$�1@[�=�~ɣ���ʬ���0��'wհ�m�&G�<�у,�s!�Y�5��X�*RC�D0!G�Jkg5A�˻˙�I�6ē$��  ���儒4K�7D�ɗZ�x2`�7D�d�)�h65�kKe�g��b�]����n�h�$��a�\�m�������K��cu��Zt�����+�z���p�nyY��)Dl��do؆�Df����V��\�T�q��r{����mFA�.��I�7J��V:{���������2���]��E�4T�

���L����O��x����s���*M
�񛅃Y-�#�y���]0y����-1�p>��]�(y7=(*K�ҡ���SZzB�F���r2��c=(ZK!߾ s�6*�^�d�,>ӫջ�#���I��ˋQ�y}�_gw�����u��Nn�Q(�i "b�Vt�#U������+ot������Ӂ�A(�U�*(�@!Q�
��DY$H ���0Y"�]�[�����5�����7�E�~��5���ٽ����}_e�i'�1�?A�qf&tb�oc��ܲa����l��p^G-�N�7���vr���`t����lLޝ֕�p]�7O{��I!�h�����O�^��=�Z����ZQ,�^���|��'#҆���Ø
��nF��2�^#o�䙗�͎�e�Emk]�W�:Q�a������ށq5K�q�D,�T�gH}�q����|f����]�����	�O:�h��[4'/�m�=��z��1㯩DΈ���YѽK*2v읽G��h#�}�6�*��ۈ������ݹ[�6�nr~����|c;d�雜��Ty��Ʃ����j���嗯j�wZ-E�����T`�Q�X1"�,�
�Ӛ�{�P�澱��� {߀?gp��򝏨z�:��Ӊ��7.���Jʨ͵Љ/t��/2��i,�|,��$| �yY;ž[��;{�M[)�P�p���h�3*里:n������Ǳ=����6�:��s&Y���lӎ���)�u�ռw$�UvEN�O� 6Dl��F�~������նivG
گ"�j��A�����>�]����\\<S#��F����^u\���|z�+���>�t���Y3�X2��,�����}ΧL��ם�o9�DDDB��P/��w��{o�&<.��&3ӎ=|�^*F]�ۺ�z�:�vW�^+Ʋ�����V,{���F��r��V�������X�����i�7m����=�ҹ�^co�ϫ�����A��\�w�^����n�XuAD�"#���, "���8w���a�[��ᾙ�H���%d�l�3�S��&u$��˵]�/���k�ɛ��\�]�HW�2>����A`1RP�s�ν�ݯ�3��/��y�Wws�4på�g:�t��v���\�}(���Y�F9��o=:������\�;��_?���W\�SmBH9��e���znB�P�{�ٗ�
�WTOVU�#w{��G�|q=�}{�������9��]sً�ܼ���0��VG7��Z�hX"��"�$21�!_}��z����Y��ߎ���]��[E"�;���d����
��9y��yq�-;��)���3��C��������Wn��}�iֹ��CoaXx�7���}"�=���:�5�هΚP�uw¿H�����j4���w�oY������b��b���B1E`(��#X� �E��ٟeo��s���:�ˣ׵Lkp�F{��Fi�;��g(��t�;c��ｐ�=��5�_>�z��(޻�3��S&V(�i�}����}�}�׫��ߚ7����@QaVu�h�ߎZ���qo%V�ֆw9I)5:�ndܻ��)��NuI��]���cMm�ض��&����$6��X6�6m�H   ��52��%2j��ۥϻ��������X��޾�)�uslm�*�=O��^[�/�v�������ȣK=���Y �Ox!�xH]w�8�Zs�$n�������۠ءY�?u-b�fBz�B���=uo��wY���GQ�E�����^}y�&��vG<��_�]��\`c��U[�w:�:�s���ךǔ:�pM�WoWþ?H�H,���@P��}�=��a�]�N;�w>�� }�o}���{�7֥����m�@ʜ�����;�������>�3��*qU�ԯeø���6��A(9��A��8N�rV��������dyT�uYF��5Egc2�]��IKO���>\�T�d��}U��U}�Z�5g8���&s�;����Z;��vb�
ه�;a�.��}�p�ԫO���}Δ�UM����^������r�F��poC�I���sX.tl9z�0����|ۧ����{?+ @����z֩�k��͛c:sF�{{�Bm��ۆS]}��#\��s�:�-WS�So&.(@��۷�w��=�ޢ<ˑ[[�5G���mhP�x�T��?Gt��y�"R>q�p�Y}���o�߫^��9����c�����$b
�M�$)R��}�S�}��kȢ,X
�� ����Us�:�5|s��D|A/,�!^|i5��Z6�v@����±B�*b]H؞�B�����j����C;������~������[ݜ��g
��i�x�Ԗ��slH�j��w.�����uo�Ϳ����HV>��UV>w�wI�g:8���ű��F����:
��	f��A׸7����cAﳦ��I��A�i��}�r����=���W�@�'�
,@�~�zZ�m%�ivs�����(�U�b��6�5�������f::�,.��1�7;��b2wcWG��tS��������3^����}�v;���vH�������w�B�G�~����5��!� 5ڭ�r�
����^�W���<�" �,�� )�2)$X1�
�`��P$b1 �E ��#AU����y���{�r4S0�d�)~y�F��u���C� c��'��ϲ(zw�S�y'NK�v�f_FY��������6t�
��˧��O�5��F�T���c��u�{'���K��I�V���^�k�W�Ds�=
���T�^����O}]�
埮����	�UA���--AEDTU^U*�*�"#T��}�]�<��[���M��8c�vt���}M�7oP��|t�U]�Y��}W�T"�[�Q7�8NΝ�]�A���)t�础��yQ�7���m�cklsmm��NM:�uc�Q�~�^�fEϥ�܀  �*Ng���V��x�����/�RѶ���u����."/���=�{u����k9�ˣ��޽�y,U��
��2E �+X$H���\���5�����}���dA�,@���n�;G���IG{��v��t�͏$@�Ww��}�������뙽��&���:����5�wY1�7���x|4{�٫X{�_�2��]����ǚ��"��1�a�Fp�}�.�ex��%ca��]���w���q�Z:��q	C�ˮ���O����bEdbU#��2���O��7��R�P��{��>��ڡ���~���e�H꣪Q���;n�Ne,곱_V��s�큏��k���'%�3M�N�B�眦q���7@9a��ЩP��n���	ٽD�R�Q%
#�V�f�՘��gr��S�[h Sޡ�U�`Ӊo�����Ii��g�˼CA�7���FƷHZ�����)���6�L�y/,�yB��{Ֆ:Ш�k9L<�&�� S�:���U�d[���� m�Y ��"��3��:j��Ea|�h˪떝B)�u����x�}��m�:"�ē�J�*�v�M�<��)S�C�B�$3u))�E�	-S  C7P&��^�֗EV�yGp�z�]���QU����c�WC�}h��z
�T�up����M�'l@�x��^����k����C/��@��v�^Rw]b�/�s�2�P5�S%m�cD�P��`��1m@���̃3�&�e�7.�u�IL{Ez�F)��wPr�ɦ_�;��aK�y�k~���B� 	�L�_7���˝�Q�#&(�7�n��{ԭ�0���{��w���Q�-< �`�IZD�LHFd�����m� �;&f��A-��-��؀Vr����]�nSQR�2�h"�:�p��ЬV����Ǻj��G5���Uӥ�uԦa��r�t��s)�U�3��S���{������2��ٌˉ�	�Z�Eʃz�5�ѵN\'Svwz@+-.�,vؤ6nX8!��3�$ ��W�V�,�r�a��Ѹ�6�X�N�ʥa�Vm��;k^�CƷwa�q��%]��FI�ܒ��6_�q���v�"L�3;/rq��Kκr��<ʹ�ao����7�kr�J�wi*���h+nƌٚN�jԀ��lu[X����ڷ�n��]�d�x��$Ӑ�C�6�辛�u�R��b��e�څ�i�ÿ�Ƴ���Ws����f��1F붝d��Rt�b��#��ŷt���(+a�VM&��]�vT����k���ZQ�6�J��2
�A�򤲪�	Jآ��9�?�Lo��>�j`��eƕks!{��J�Jr)�h�oD��j�M`T:��˽㸰5df�%|��c�/�R�2Ѷ���a<��ŷ�������p���t�Nm��B:���ʀ���
ᝦ�u�۵s�_"��8�L�;�u��#�s+���7��97�Y:��m�rwʶhӍ�ݝ�oI���o��ɚ�۫�ݖ����i�e��wۯ��ApqE!m�fgda9�J���[c`6ۑ 4�6� �  M�A�     ���m����i4�    @ m�         6���1�6��`    m�  �     �`6�p��p�72�3�2�sr�	�`  @  	��c�yr_WcQ}
�ɝ5��E]k|�����w��W�&t�6�84���n	2&�F;����y�wwΒCh@��`     !� )�m�d̴�M�N�b��y������EQ��zGVr71�tەxu>�7b7~��B��ܼ'�N�w��H��rh�d~~�;�R=�ky��^|[�w������d�̆��l�r:WX�y�&�����5[=�o���_ݲM �$Y��=�f�~7��:�T`�+��+}ϱ�����mu#���8#l|iծ����4�{!�V�#B���;NT��]�KI�q��v�]�L�0���{�������oҏ��Ǭ2T�ڼ�j	�N�H��K5�O�s���J
M
rro*x�d�����lI ә��=tO�N>�鈘��?{�~��fTV��ל˾"m_���J*��Èܥ�2v�IK�kd�z:V�� 
HG~���u�=������W>�m!:�;��)%:�9����O���t�����wr{r{6f��[���]#��lj�m��7|��w-D�q̆������l�����w�:��붕�wȫ�g��P�	/����c;��}�ltX��g��꙽��V�g̌s�6
�,QF �dA,�^�7�9Ͽ��H�P���X�����>����Y�����7�%�=å��V�1E�{�j��N���Ўu���L�y.�Y�Q)�}�=��'�0ɰwu
���j�J���m3[l%�	��{_����)����~i���]t�^\�>�l��]�W�_Txz�[��쯠~AdR���� ��1葫�:�d�k��d���{�w=��˺��v�׾�f��}��x���sU�3�}��u��$�,�_eb���}�5��;W���ݵ'q�˘n��/j(��4P�J�RΧ���y���m����A���uw��3���E��V�gގ�'�(�X�z��*�Ş[v�>ܼT�]��yD&׋�}��o���"(#PI�1	}�w�y��y|�q����\�$E"0��� ��Ζ}����N\_�y��k[�#^+\]��#��.����J]2b�l</su<P�#IVZMXu�gG,V$�e�"vs=�Q����=΃�)�z�5��^#��U³zQ���s.�e��wb|2��U�c��=���K��='Ց�^{{�7�!��J�ED�y�r��珌�����yIY�k�N���v�̉�<'f�L�o<��wq�4�9N�/���+���T�sm���������<22M�| �B��?f|������_J������dvr�-s��̕7�Ν:niQ_���OY��v\íؗE�ܹn_Z��X��֬q#�>CC`�w��쥼��GC�����{̍�ȣ���T`n�ln�";%��Y�o�|BI.�鏆*�D`���A`
 ��H?	�;̕��d�nbn"
�L�k=3���f�Wm�vy1�+�ֶ)��b���B��;��*��v䨆jݼ���Z�Q�}wں�iC�{6x�ֹX���畹�n�Qs G-7}���/^�yK�Ii���|g:����{���'�ۤ�Dk����Co��{��2���_���,�֝K���.:z|Ȩ��Jo��Z�]�Q�6��V�]N����xmC�)��/���ܳZ�O�?N�8���w�	s+�;���+` �>�����^˯n��`�8��D\Oq�}�BVg"s�r_�ೋ�v�VW
��+z�}�BK�i]1E����%��26�         ���LJI�f�e��1bq@ ��!B�U֗�f7���_|��o��4�� �1TUdATc3���v������ A�	"�����˃x9��$׳v2Gl�]��#F\^Ԅo+���yV�5/Q��������| =��ykփZ�qٗ\O��{���������,Dkv eT��ڭ�������=�îC��2���N uQ�����7[<r��ޚ7�T�"" ����ֻp���yM{Ո���Z�g'۝!\,�8���d��;�v�a�[O�bf��C/ʑH�o���^m��p�ͳ;���a�9�TL��_������~�u��2<*�����b2��M��t+��������E��I�3;�x��PA��Q�
EAb,b
A�D`�c�D��b*������1�*�����E`���"
�R,
T[K�/�����:�*G�*?�ޙ҆j��De��Ny@�����-���q|�f�.��K��ye:�����*�m���[�W��f��}⤅��!���w:n݂�����<��zm���lP;(Nu�x`��������QJŽj��ͭ�/ۺ�{ϼ-��P�����Dw=�Ly�B��j�4�n���3�2����.�C�О�%{��z���GOfЦ���Lw�&�l�sQ}��@�q��;./MunC*
��'KV�j�,�  O)>|{�ƶ��#]������i,�Ql����g�A��Y�z��2-�<�+���{�N|��s�`���0/N֞�v���+-�y���V����۰�/V��������c�3�"$U�" �b�QQD�Q�FE�cE�Q*"��b��,b��#EQ@�~�9~㕟���{�m����E�^=���%Vp�X55]�d
H�f���a����;[�d�������R��4rY�V��N�d�:����3u���xl�t��h�����Ƕ08t��=�d3[Y��˘��g�Մ7]�1�2Z�����;�=��κ��kGM]���l�̍��]c�����?y��%�` 4}N�d�tݙ/�#��> F��w�gJ�_�c��ڝDʐ����-���m�lH�z�����r���&�[�9�.��m�k�1�:bVo�^�Ok��u�}�{~����n���p;`��������S]iΥ����y���=�&��z�W5�x�u�AX�
#�`��UﾭW�w{�o;���09"�AdA	"�Uy�yֻ�?hz]w���Ou.W�}q�}��C$�měZ�׋�wfD^�g�VN��Z]˺ ���w����u�r+��j�C�e4X�f$L���9I۩)�S��/��C�z��C�w2����U�K�6ӡ�~.������Wf���z�}��9V�@BPI�;���ӊ����ݭF�~����2����W<`;F��(�/�{\�T�wǿ�k�暶axzf�m��wuӦ�7�:�I��2����]��3\���1b����xq5�+�Se��w\_d~�}�{yA���U�>e��]�LY�d�+t!����P�QF��=�x�φ�����+�ˡ��[���+�{}D}� $��(Y$I�迓ǵ�̣�՞"�`,X�
����k"1cDvVq�V���Q<��ǻ���>�<�|��}�pT<����o7��w�eT�S��7;��a�w+aP����_h2�;���V�t���p�>���mKTە*e� � i   �@�s$&����j��x  )�g�fN�a{c���7ޅ��k�v��fFJ�EO]43��U��F*ka�م�v�Ms��^�Mm��I�z��_d�b��]ë뺡[ƞֲ�K����� �n�4�2k���C��1�9��s��R��W�ףs�L
���\��{ݔ�GA�H���;F��h������Əc3��I��.���B4\1C_�Ӝ/�L�&��[��^�#y�o(p�u}��+.��97���PC� ����C%��cAF(�XH�����,T�A9���7 �5M�ڀ�#�qF&\�r��T6�\LA�̭)Թq��qd巏���}ʇ{�����ko���;��'�$PO��k����f<櫝�"7~I5
�h���O9[%������6���U�N�����K��s*�X��=8��+c�i��Z�G^�I���6�#���GݒW1��Fn�܊d=�f5�1������{B~�9��'���۹�v�J�b�mBy3;�L����"��C���]��Y{���[߸I���UCj{�N��u����˿d,��&�u�"|���ٖ.�L�7�Ԥ�]aQ]�m��+��X�k{�S�����'�� �����Ѷh���wK&;�o�\����t˪��w��ส �$Q E�"��;���r�U�����`�H�#�=K9�p9��|����{��'|WZ�����;�7����FxI���T8Dq̥dVen�o;n�r� u��;�/�Eh.�t���Ur�	x��Z=&��3֫���o�U�Co��vR�â�
W#q�ER�RgP�DmH����-�F	[�3$�����:W(KX�j)� ��=]r^��ހ5$�;Xؗ��71�e�P`�$��䟐S�ɬX܍����Rh-����w[uغ�L��<M��<<��\/`��k\�`�xe[��j�B�*��WvPW���6oZI)��k�I�!�Eܕu�j�/�n7��]�u;���N��A��̣c���t)*�*C�Ch�T(`)Ungu�^��u7ev��Uv����U]��l�=T�|�Ȏ4�6�|+����et�/`�,Sp�m��3`���ʹ�;�[��˾�Z����ڌB���8�����\��C2��f>�#�"���qs���Z�)�&sWʷ�<�y%oUqCM��R�SCj�  d��L��	��H����� �H!��@�D�ى��;P���Bv�΍���u"�F@�d,��l4�(-��jD\���(NJ�n�K�XZ"�B5��0Ծ,�@  �_aK�Te#�y� t�ì��y���Y���T�p�sh��35�錖!����sڨ�]�7�'��4	��,��]I����[��ӵ����^�Ȏwe@u�JRq�|�U�$+���b��r���T��U{&4��{6�]��f���2��|1n[N��.�1�mfӜ�AlJ�/�c�Vk��ci����Ed�a��wFV�[m�����H���ʙ#�&��]��I����
�6��U��:��(RS���6�}��HN��-8P�}t�� �xgSXf^>�XK� n�O��H2ng!uz�̩�O1�P�[V[:+]�ܔ�̨�C����;!))�؛W��f���O���W1w��3��n�Ǳ�Ή���w
��:���;�*og`�ݛ8�Mu�ǧ�ݬ�P+��-���7è��+f-S�ۑ})�%!�o5�����J�.j2�R��D�=#��2��nd�]��!8sc�'
���Vl��̽���ߣ���:�WR�g)���yٰ��AFRj:Km[b&��KO_n�ko"�Pq��	�������(Q�ꕸ������V�b�qZǝA���˭�̧�qeÆ��iڃ^��U�8�dr+� �T���g���=s�ʮ���}�*�G6�rsB��Qu�s�+���U��h�j�*۔5Q������+�r���z-l��cV\�i���;�wr���Oe�S�pTvmhւ�+1i+A�gt]]���唺�qa_oEՂͯ_�#�	��ɗp��9�y�;�_�y\}k��^_���3�'������~��#����n�ڱ��vl�8���Ĭ���VF�qJ��M��z>������������$㐺���Ȉ���Te�A�{��]˞�]����8Vk�w�R�2"����Y�����Nr��vg�L!����"��1��eN}�䉤 �_�9�s}����s�����pbDF#�1A�oG��w�W7O�z׵.:�1d��R��\����=Yp��h�U'���o]�z���*�v�[w�O>���c����)��k�g^E�*�[�/6���=-Q����]�c� ��^{>3�ⲱ��ݵ�KZ��\�\��6M���p���1��r���[{��@k�k��S���ه�lZ(�~R ��H�����v2��� �����F�UTXeFڑ��w���@�JmLmG�eV_\O��D2�wb3����9��O'/�C�0&7��gݑ�󁏌غ
}�{�\�z9��s��M��L�`�L3yu:'C���z˼�����a�d��U��ytw����ϡ("��Ad̯���UEV"�)"�0`���T}��J�DI�7Qj���
��,(kR�i���Nn��$��(�ɪ�R�|���m� ��9�����3\��24�=e�qp7�Ѳ�7Z5w(e��awX)܍�!Zxޖ������¾1H
	ww��Q��y��On}g�׫TfB��1.�!�(%�s��xeu�dj|$�3�۽ut2q9�s��W�[��[O��whٱ�CI 	L� �    m�  "I�����ݹU�[��p8D7��3��3��O�|~���������v���W��N�x�mZ1��]����ڡ!���΂Tu���C�NMꈜ�C=��Y�gt��r��p��ozZ<�A���ޯE��%�n�5�;t5F̃��n�oj�G7DGv���o�n��{��x�s��E��	�"�`*��
	;��{�]�W}�ߵy� 8��B���*�8u���W��=�f��^j]n�u ��4�z��Nj	���oQ�k�׌�]7)f	��ݗ��W�&����xn]?FsGp��� 8�&�%>�.�[���tߪ���i����~��+u9����o.�_�6냚�e����� ��D�Uň�*(�X0��U#A1EQXEA�(�aM� R(�X��!RSU����EDF(,*0R
�����P�C����%Y��1unB8�\.N�3Z;pR�-���%.jOFrf�e iP�㔮0�����l����35=6���Ǩ���f3.6��3�>��9Xj��:�x��7���%���ө3_Oc�����u]�"F���� ���9a�5��/E��Ȱ�ma�EO^j+d��%W_[���3��W\�rG�Ye�D�]��=�}�RW�Ϯ���=���{�+Pb��V0E��QF19�s��kZ��*9�U�n�k����pY�ٳ�����\o�̼  cb�\��ZW�}#�����oz� 9��n��5���5ۛ������-@���h�DgA��!�9��=T�����c�����w���n�������s:����`��"3�������U����+^��R@I9������Y�z��ﮯg.�����Ъ%���� ��\��]��e�/W��{���d[�p�
�SsNċ�l��l_nn@��
gP�U���i:��&N�~���*Jy[����u�v�Pg;Q=���rx�FS,7<v�=�y����.�>o��~�HYS�Ǟ�s�π���?|�X�  ß�}��(�`�PQdDUA�����}�٪���fe�Q�S;���Ӛ8���݃�����P�#oq^�8�ϸ��ۦ�j��!=É[*{&�YyB婳ܗ�������/>��%�׍��i�r�F�^�>Ҟةl��
\�����֣�{N��+Wz%�5��}��fT����z�N:"cMv��Ei�h�h�W�
�λko�u������ā� ��k��5N�vU�eq��G�qS6�T�Vu�Qһ�Q��V���X�7�u���k-9����x�Gp(�tW���g�)�-D�v�}����]�G��.f���jo;����gykc�����2ϰn�;Zڋt 2�-����Wo��1?Gu������""���D�H��
Ȩ�#UA#';^����.��)���j����N뻝}@���y>�xmo�_Ә�3�s��P{��'0:;���}�t~v�'[�ë������wzx:�<��/���D��2�����	,Z�zv%G�g����os���(���;&���60�*O���� ��xJ���8���U�6$�\r��r�gdL�����J��1�^��v�XV��_����x���>4����K�ڮ.�ٓ:��������Q!��hF�d]� �uo-]lW}��i�n�E*�uS[�:(Hr�iK��	&H6�     �  M���$����j��qN� %ZQ�\�>�G�9��,
m1��t5�-Z~Ù������<��_r^�A�Z��'�\ۙⷦFq�Y@�U}9�+��EH���`� �Tw�}W�������b�cX,`��ʭN�4��b��lw;��$i(�O����jzӿe!��(�����c���3OTZ&z�V��*J�Bj�M���j�q/K�05�z���;�IkS�7~�[~����V��jȽ��M��ͬ����5�ʜP.OE�`$��UQ�^���_���/ǻ����[Ro���m�N@�-I��]�y^k{����ép������Zzj�S���J��ڒ�"'K	���g�+���1�����Oe���L1�ѭ&�9\bc^t�y3���:�c���*0Naٲ���G_TdS6&�,�H믞Y�M7}��&H.��S�q�<n�:�Rj���ר���Wy�|�s��{W�������������(��E�XŊ�UF0F�XQA����Z��<&�AM��S�b�I)�b̬{)��G���T�;��׳��{g8:�&�W�vl��8�����4���^�yS�~�ŴHZ�z�7^ί�Hղ����Ϳj��8pb�����Q��r�� �)�yk�����5^��9�f�7��FN�m� ��.��YԘZ�;:�d�c�K��ܫ��vM�ݠ��=��Q�O���%���q/����S��Fv�O�+Q���=4uǝF�y�sG8߮�)���s�����ӯ4���W)u�5{�p�<�ݰb��4l��t����{3��b�r��@X*ҝ�8�Di<�!ט��{Bs�
0���;ѹC^���m,�k8
"+Pb ���$Q$B,Y$W��S�ޏ���:�{��� ²�p��j�k���xE��nv���~�a��S�i��w7s�+z��FWޙ�Gt&z�/=��6���Q�^���Q�Ec�צsw��  	���!�aR�[~��"}ks��&��>Ů|�vQ������}�v׍o9�m��,H*(( ����TTT�s��7��X)B�<�>�����펜�Ӆ�m�K-	��q�Z��b~,�R�egg�!�ofF5�Y;{�ŨorN�	�w�6����6C=W����85	����݇Wk � ~tE���]��r��Տ�9�����Jm�o�N5����E�)��޻i�o��vt��Y�(O�/+4�Oq��%Z��Y��x��f�l�� � ʹJ�?�E����	@V"����$��"]d�EO
�k�����3��.��D�v�8�3�(�z%$0dP�
'�ة��[ڵ4c��Hʜzs�x���z��/(��߮�u%I{ɨP�y��L���ڈ���/����i�D��o�V�eZ	���m��/��ѩQ�.�	?|��e�ދ!u+����aq�릎���{AO"��V`�漨�`�힯n���1ӓ�v1b�J{(����Zս�G������� �	��G-��oTV�{U�Ȟ�v���Y���+{/r���U���=�6�T�o�O��I$�	$�����HHI?�TB$?�� ��$�		�� �!BI	��$$�!�$@�s���	$��_� @�I5��	$���x?������I'�k������K?��� HHII$ ����@a	$��Y B�����R	$��?���Y @�I?�}��?����I��)�I�	$���B�I��.�$�O��vk������!!	�, I!$�~ @�I?������	$���I'����/���������IzO�a����w��I�L�I$������d�Me���<�S~�A@���@ ܟ}��s��y�P���)I%��ӻ�קU���
:�fZbٕ4�cTj��Rm3��VUP�͕k�鉥�v��׶�cvl4hKe;f�۝J��*P�R��Y�6�m�h��U�X�lZ�fUa�Z�T�	kam��j�Z*��h���e4�Hfe+kf�4�SM�Z3R,cH���J����]V����ݠ���kd�۞������W�޽���p{�����o���jn�{�g�yۻ䯾�{{��3r���n��xwG���+��W�m�o���}k�7W����.z�կ�m�l����c��w���{�t���+-� ��P�s  @�;���B� (�� 
(z5�9�|�t>���;�x��^l��p:�=�v|��x�^��8�F����w��xB��Ɗ���Xx*�Zdi�����Z{���{z�	���^ �q�����L���齍x���/����}^���xsl�׻�^x������>��x��>���{�J>��������|�}�ٷ���J���Zj�kY�Т��n�Gl�K{���^���_{��z��o��w����3X��7vv�����7w:�=޹������!�ڱ��=��n��7+�^�9���Nw�Q]5j>y��+Y�[hcf�F���0(>���h�1�sS�@C�|��7�o{�W����9�Ѽ����l�����}<�O����X��}���n�7�9����[4��G�u��{����k��<>#��Gn8姮D�1=tv��T{�����o��OXѺ�������x�m�e�y��־ڹ��i��;Q�����͐(�l�<��@Hy�]��n�pqt3׾���d�{����=��^0=/y�ɢֽ�E�����z��uOM��)����l�klh���u�v�Cl|{�=����0g��o|w��]�5kS���O��[�g|�z>{;b��÷lw����k������}�����D�F���k��pf��[Sm�:ݴ�:�ͣ׻v}���������n��ϯ{�Z���s��>���o���z����z��<X�t�c��w>�U���z=�[��}��@y��>�����|v>�c�ʹ���o^wm["����u��w���e����>��we��}��={���������=�uy׶�>ݐ�n�޽��^����w�g��e>��:�������/{}�������=ݼ�Ϟ� ��L2�T�  ��A�J�F   ��d%*�� � ���RU@�@ b�� Ѡ j �iL���4i�e?������4~���f��v��<�����5B�k8�Sii��sZ��DAC�� HI%�I $��!$�� ��J�?� $$��jI$!$��!$�d�BI���_�����ո��6:��n�'.���*Լ&��L����2�~�\n˘ƫe�o]1�'�t�ȩ
�YM+d1X��×M5�¦�^KpYz����j���5�*Q��m9n�E�*���0��씾̛�n�lp�5���ڿ�}2M
�����`�5n��K�b�$��&�¶L��ُ)Fn�����V��:)��#�/\����4QI���dc;�)�'�u֊��,��s&ŀއLI��P�H�fJe �XN�+q���OS{�����6�X��*�M�8��X�IYKh,�pt�V�r��k�sI�e�6.7�o��Տ�lZb�̈́kG���� ��d�ܢ��y���P��Ɖ+F}�.����L��(�>�npX���)^�U�L�ɛY3(32�З-<���������7�0m����lWV�f[�
�-��e���j���`��k��kM�0�V4�`��l�HZv�e�C������S��oj���ڵ}yi�q�t6XH���.�)Owj��z'�i��Y�@�l�}5U�~�qb�˴6�:i���3j��N�p���An�%be�Y�����R�k���($L`W�
�l��.�p�<~t�^9HC����TR%3y����-����op��m���̸���#�d�BDenbӭ+˩faȶ���p��1�nR*�+�&�F?�$��Z��S鲣.i#M��Y{-ѥ�:���+$�V`���;N��e�#2 �(\*�RaX��������.���ܭ��:հ���OR�����aʇL�0n�St�Ec'0�~C�C�K1�p�t�PU�K�C:�n���'k"���vK�e�M^>9J B	]�t�S(v�A��j�~�~�e�lb��Ԏ��U���iRL`y�tW����-!U�Y��P��:��$���q��i�Um��h�3$̱�Vh��"�\�-�2�Ֆ)���T��)#X0"wz�r������w��v�J����FޫP�Zou��So)�xLT�N�^-�ް��*�.�Ʈ�Yw��5p�H�]]vP6���k.��#�,=��N֜ZU���]7F��diV��r`RX�EP��s_��v(��)�G�c@�����È96R'-��3i,�͗B
����Wέ�ɐ
`ee��ԤR�XЖBùl�q��0�����J�,�hA��YTZC�	���Z�^k�k����-^!J��D
*۽���e��-;eC�DL;��	���h[CbL�١����oe'�j���\rf	��)
;H�)����1�`�y����h.�k�ڠ�bX9���6Y :�M�{J�R��]��n��VK:�ku������Ŝ�P��)�Ѹ�����^:��xI:�t�U�*՗m���=9N��V��x ��2�n�N���r�@aܶ�V��F���AW��@o(�s���1P���ૠ������vأSq��4�����v�n�ᤝ�g|i,8�S*'�Skv�H�ٵ�-éF��iL�3s+hRz�4tHm�u�4D���\љ�Q�6�6�K{�c� ���ud�U�Q�A܄�[6�\Q
*���<) bj�Q4� `H��y���T����b�6��<D,ҳj�eٕ{X2m��)�W�ɺ	��{��c:ӕs暡G/5�2�H!�6^�J����Ǹ�а���
v����f��X�h��oZS��1�#&޳����p=ǔ)�7�����]���=.Q{��+,#X}^�1;n��H����Z5(�a,յa��B��m��P�����Wg5��j�J��������(8��ة�����e�B����嚋(9�oD���f*VJ@Vj!�u��M�-
��u��q�0��C�v�溷�º�խ�2���q���,V��]�ڈ5�;�1T��\*����i��D���tFkd*��Ib�yD���L&���:��um��n6�˟  ��^��
�5Lįjtj�U��}����-��K?sciռԹ���xzA�j�)�-ut��I�7��Ef⩁�d��#� �r
��l-���[J�����raW��/E:*��OiQ��*&1��R�k�Z��i��K׃gr�δFl��o{�(�vu���mضM��DK�7$����FӍ8s���ym��32���2�s[�Y,Y��.Z����e��ϰxje�;,�+�-a����Q6�#6��wC�f�7�EmI��X�JfX5���76�4l^1r�s]6ꝍ�F	�P(�o^X���u�w^�A���e ^��e�'�*�4"��wn��n�Ұ��q��� �-陀���g��D�*��MG�l+��ͫc),��ʴh7��v<�oe���c)[Ł�FM�Pd�P�N���MV�dA�����+Yr��X#jxh�M�*�ŦM��v۱h��?3�J9{I5�u�D�E�S6Dw%�f��x�Ь2�!
'(Rdv$Op��>��i
=�o�����yG,��d�,��M�����H[M-n� �-4��0n#�d�Bz�r��Ym�m�k����%t��v�:���ЙT+�+\���-�v��=oU2�d�@r�"�e �#J��<�)6��G5���r:��fU�S�;OZH<7`��P�!�פe� R�N���]�gi��b*K(�Lډ����ŗxIЭ���k����<ڠ�^&r��U[�f�)񶍩�^�"&hIh��Łc] 7���/�6��Z�?�H�D��K\�3w�y6�m�4�fAx*�X���͛2%�L�̐X�ڿ��� ӸO�	w�}�i�sIʕ
�eQx�܆R�KQ� %6jn��Q��6�ݫ
$�p&��Z��(0k\)e
�2����f����mU�b&]��l}Zl1[Sә��u��|�/8w_m���<�nb�G4:��I�a�y�'�T�5�Gj���Ť��������f<PDr�ުG4��1���;��4��[�K23RֻcrةX�`	��IB�Zձ3NJT��Z�-Y�R͗4��SM6e#-�,/2�zǑ��5n8skr�Pz�M�0�B�[5z���k�G#bjs5��u.��F�/boh��&O��S3Kk4%��(����1GXp����9X�ݜ�O>.d�f�3�Lw{Mpq��^ۖ��R 6s�M�w�0�Q�M�Z]1T�� ��T�O^�6�J̤�j(�$b�+8HY��:�G��ᗛ&�jsK�[�}�Y:��ajr����yc5�ي�
�P#`1[���f9�5�T��b�b��r�E	��V�.c�����2���VY9��k"��`R��!�{D���B��?Ѫ�2�r��+�كb:����.��z;�ef[F����f��X��$��VC�����Sωfs���V�jlyr�z�[7TqR0}�f:ګGzK�sg����Xy�0��v�5S:�i��ous��
�6���MxaܽN_�/
� � �8��(����Vf��A��R��e<
����%�?�N��=�'TE:2�Ow���aEu�m��V$����Z�;�W��X6�ú^��
XU�Ɇ�4w�3[i��ޭ�.���P�+�R���2ܗ�I$EF+c[�$�qU�Cj͹��zft3;@9y�̽��¨_rWե��5��n�r�a�v��y@�ZJ�Ph�2M�����@�u�Y���D��e6�:R�!�+
�Ne��< U�X��޹ј���z/����&�gw
�FO�i�I�Lܼ�X�����p�E�ۭ�X�M�a-��ٕh��-��m�3쨣��̬��TM��l��(R�n�P�7%9�rGneCu�ܷ�D�u���Ǥ�y��sZyvn�aKw*l���Uz�4��F^)��g��+K4���n��;���q7	�`ef��DyZT0ѭ�݆v�W$�嬌ԕ���zE�HC:��� X��T_�0%M�EHe͆����Ĵ���ҵf�Eo\��ش�Uݹ��T3݌�j/-��isn�؄Ǳ����*�OU�Vc�\4쒪����4�U�o�j���W�L�u[{P^&��v�=�0qN�S�!�թ�*�Uk`�e~R_
�mѯ�2�:�9&#�)P�̭���w9� ������W��|��9�Å�3SĐ�6�m��}�h���8u�����CQw[�%�	O���R���>n���Es�4r���6�.��m��74@dĖn�(�3[y��̆���R�i1ηo%�`b���;Y�Hcr�6��Y�H�tF�l܃V|@����V���$�0$�2��G�u.�:,ǛM�uk��ˊq�9v�)4��̒�N�f��`�����t�ɴ�%����@����lķ�'i���s���&./���-��V�������q��*,o��5;r�6�V^��9o+�K�8��p�@�X��oz�k�`���L(�����.kFa��j&I!���5�$�=�ml�%���+����6��hǷ�;>�7�/*Q9�$w��#qƎ��Ӥ��ٻd�Y{�3y�����ƶ,"��V3J.��T��
7)/ia�P;ؠ���b�4���Eb�n
sX����fR�]I~�i��>�f��V��2J7.D�)�7*kiPi�	<Y����+��K>DSy<�.e�v3՜�v���ۙCLA��)�i��	�\�򈗏���&܌�7ef<x�7��V��$H�Sj�[)�Iu�w�M�4f�H���OQ赚�M�/�.)ҵ䭸򂻎�-�cY��h�lW{�3��tzZ�݁L���) z����ɘ@;��F6�3F�����I��n�ۦ�r��>�=aNn�8)��v�KFڡ��2�j�B�ɉ I����0J�Ȥ������yPMopVn\����5�'���W�5��@�^~���t��5I`B֥��1��/1囫�̡��o)	����ŧ�Z?��#�4���Ka0VǶ�ěڹչ� ��ؤ���7-Kie�㗉� ��vд!��'(ƵU���K��"�� �:�K�Te�]n���Y��ѷJ�:xԅ��E�E��w&�YW]f����UZ5KU,d�������DM�1U�5����sw��s���to�,2rx����z��,|G�@�Q�tV(��5�G��i���l/N+�!2Xj�Z�y�t���+�k�!��NʐV�a��7т��U�aӹ�;��b�U��5��ג	��%3	g29�uR�i�k��I=8١\����z��UX(��Y�[��l^z�Bq2ff�	#�gE�J�E7�F'������y��P�$mY��R��%�Ga|�-ȍ[��3�4f�{�[md���#�e�3x��O5ܔ�G��*���Щ��IV���%��[�Ϝ��-_L������{a:a8��3p�G��У�j���[E��%�,��zå[l�V<챻�����&J�[�%d��2�n��Y0��xȘ�����⊄ۼ���J{�Vjh�WAl�)P�mmӬ��N�A�5�)J.�E�tStn�^i/�,kz�$��{����R̦U�;�6D�^�Y1WB�*Z�H��0T83F�d�(!A�YL�R�Xm�-C��U���]]X�6"�l�BYp���3�����"��j��v�$�R	�Xn��2�e�[gf���#��텨�5a�c7H��1�[�-m�cv��/(����ţ�At%Ƒ�<�ݺ��2T�R�/^�T�������n:�E�M�dVzC��Y�d:U�flY��p�չv�L^��ZLj�b�Ba�yX�bXu�v�d����XX�q�t�n�a�.�
TU��wbts8��.Rɢ(T�������J��Y�"˺JTq����<�N���f��P4]
�J�.�N����ՠ>겵�lݪ�d�>ݰ�:�+s�B.���M�����be�D�5�	[�^2v]kܭ�1k����p$�H�TI� ��Lj�j�v�q�Y��Ӭ]j�����=�Y�v��a�gM´���������<Ÿ���ʕ.^����$p��30ʦ,�R���6<�`B�y@	Z�č:7ʫ��髼���M�m�Y��#�B��w��ETK�$(�4��<��b@m��N��u)��JJҝ��E��we�
��<�0��6�W�<�Xؓ�
�*������&1��M�P�������%��4����z��`�b�)�q��z��_/��	+��T
!�DDm0d2.e����X&�h�87cݣ.���R�{�\������Ar����f9�8����j�����B��i����2�&�D���ݷ�ly�0נ0V0pí��f�БVQ�^q����o{�� h��:��C���VP��Ê�nd�[~ȴ�m_�~t�1 ��W��z1��3�7������)��2?���9��(J�%[�o���tV�i�.	�VVX�-4��PĮ�d���c�^�F9�D�t�֓�Y�KI�O(w��VT'"�ijy��A��� ��t�u�͒�Rpe���*EB���:,�����ee���ϊ**5afG�*�V!�.��w�Sin<7�-Q:x-ڭvS2���N�n֝^�w����$Y���a F�f��j)�Qٰ�Ӻ��m�*�Kmk�m'���^iu�[�b�n�R˼. &�P�H,K�^Xe6�P+������E$�A`[j��i<��<� �n�k���]`wR�������E���@�-�elM��5
Sk{�3�jU&����1�g0�Z�*dFXF�|^�(��$��ݢ7�e�8|�d�ձ;����DB𔝴���.�үk��c{t-�Jm�9��Vm��9Xbf��ǛB�.�����7r�`�@��� 2Z�j�X���ҬJ�<�G-*0����U�����l�PI�d����mH��A�d��t[m�ۤ� [m��e��n�m���M�I&Im� �$�!�I$�n�-��m��4[L0A��I�$��4�)"�4�D�m��m��m��m��M�I:m�)��$�m��m��-��m�Im�-��m��%��m�II&�m��-6�m$�m��I6�m���L�N�M$��[A�m��M��M���)��P�R�R1,J����H6�$���� �Nd�%��RH#(�����K(5�d
`:-��&�m�jd9Rm�I&��%��9�E�!��h�IS�4�����URHȠ�9(&S30�L�	��i�!�D�D�I�L�Y%�:6�)]��~'�ݨfl���٫���I��2a�7�#�\퇝�B%2MSt�HD"7xr�Ε����E�2�[vga>�N���mN�r? β��XR�u��ɯ�����;�D�νp軭�M/����դfhX �\aJ� >�[Řآ@�oq)a�;$�7fŪK�����)gv�(qur$���D����ռ���TMp��c>2
\����f�	�j���0Ԇ�&6�Tⴒp��\-�׽��'I���Yy�ml�8Q�!��짂CB���ӫ�	�yӺ�K
㴱^�+nrF�W$2�R�޹�s���D��V23s����l`�M
S���x�nP�Zt-����Zkl��+q�̋M�U:�}D֓Z�Ä���gf=e�k3'Lt�]�mK���
mk{���أhlеq�#�#��B����˖��h�d�k��5�7�7��#�&�m��ق�L��O�&��Qh������]�J�x��z���}#m��6��N�76��1��B� U@a}{^lY8�;{�Z�r<�.�4�4^����DZ5�j�Й�3cs�cX��q�"%:����[B��4MX�s��|o=�����n��Պ!���n��ԕN�i��ǻEP��t�EPl������F,�.�B�xĮ���2�5:��738)����mf`S��d�6��b������&��ե��y.�J6ҍ�ܻ�ph�k���%�R��:�1�8:�!P��ۣ�s�������w9[ut�YˇFc���f�h\�1����`����.�-�7����V�^kEQ6��f�u�NJB�9�Bn��g�"nD��ns��{����k2tAS$��}�/;˨]�RVK��5oQ4�nL�*J��E	��n��&9;�^CPw�h�J)f��5��m�*#i�f�En��aeR�^�Y6�]N�T����P�������.t����_�f=nj��������6�G{�����x����P+'�tj$�t�d�$�$˹-K]ji��d��C�8��@WJ"�Gzo����`�{I��{�˛Ć�u�9i�QgB5K]������kKiTf�p,�ǬN����u�o�S�u�23���k�n��&�K{5Vt�A%wY8�L֕�/�t v�.������o#�!�*-S�>6���|���|�8�=`;���'a�g�4�ν�lGB�����0�V�|��܍ܝ�Zy�>U�қ՛���rd�A>�R9�9 LE�3	}w8�&q e��Sobf˦��нZ�I�w��q)؎_O�NӠ�f��Eՙ��WeȰ��%�ӝY����0)����'d����"��`�j���'���ܲuz�t�x�Y�����(�#Ҧ��#7�v���o:nָ�Վ�z�(���>�ı�`l�iŢ��b�˘��F��{��:��zM�#WBw�w���s�6�3l�}Z��Z���͖bW��� f\�5�{l�o6��t>��	��lĮٿ��|��"cL�Ya�O��'t%�l��{��l���Q�0�5q�gtTR�`rL'4C �&�:[�����5��sn�r�x�=$�I�3�MEn ��#q�,�1��{��h��С�X=�LuF�_H�P)�\��ُ	�;�KJ�b쌸��8-�-�<�7CM]_A���-TagR�]z�]N�\���R��zu*N�ٕ8G,A�P�Dgb`�������"3�ղ�"����N�l�]�[�!�V�}R5:hR˶�c�ݡ�4ŕ�E.�n-v��4ڵ����
�2[l��V��(X�r��P�[+`L8vc6!=����;d��#�#@���0���p}�x.>��iD���3o!�B�aT��i�dm��.ʸ�]�&۪�I�e�W��,�xfsq��6PS�hPo�"���4��٥������_wK�Y��@��_n�E�'�Yu�D��m���uB��3���j&��N(6<���p���ͽё���2E�5��;gN訧ѹ�j����WSIT���]�i7F�)¯B��1ko���w]+1L�]m�&��{h~zZj�	�ۯ�v5t���P�Ӓ��tM��WQ-���w�h��Ms���G���r)z*aub��o`ḁ�dU�'�0#h�}�:�����ꙷB�B�=�^Ҋ�=�Q����PӛW��I;t��~4A�P�%�ot�{oYі`"�-�蓰\Y�rA��!yy�/EFj�y���f�Io��w]g`Ȣ�nie&$+zf#˛�S�ܾ�,m��LOw e%m�oG:����k!"�:7�M<�î����%�(�Yz�T��:��L�e�Cg�<�kO6G�7i�4�j��ؤ�T���F�T�d�\p�=�'�p���Z�y��;�L�K;�p���P9��2h�`F\�[�R{T�i�5���Bڈ�/V=�ܝ�'t��O��6�-杼��'8��7{dt2����hih�l���~V-J}b!VVj�Ūn���U�Ƃ�75��D���]
t��]��y�J̖+gt��Mr�#�c�W��7Df�deۖ`�}|(��R�7�b�Zޝ=�5ֶ�kl�mf�N]��'>[ؚ=�B�i��.�3[����('u{}�Fw�-�ʎb��[�.ѱ�ȷ�t1���/;�b�]�!=�T�h�m'Sx-�};oZ&� �+u�"ՙK#�9P_;�`Gw�����i�+D�#���-�0�z�唙v&���gZ#]��p�Qſ�Nt�t����S�Aʃ��{��L�'$��U˝<��V�$[�Y��H�K	+�<6�s�0�f:3�%��ƬRE����yε�+G^;��\kϲ`���if٤�)����4������Сb�RZ�r y�:h,Yc��yi�[lXjĹr'�3^���NP�uw�\�|Lh��ݳ|�h�R�:�/w��B���B7(�Q�8�f6��w���k����I�.�u��3M����Q;����eUǗ6,̋t��a˻��ѝ�4N���&�1�7	�M��9��-�ŉi�6��0X��ru���%�ssz4r��y�q-�vt���J{�n[t�3V�R�/W2���n�M�X1(��ˋn��(_ŗ�Wn,��_>u3p|�2j�ۨ2�j%��nrX��Lk�c:����>��*Ƈx�֗�bF;��܀tÄ=:�
i�w>���;����x)x��n��]Z�4>��K�b"��7�ص��*��sh](�VS��!�7�,��x_�Y�|�7Ѕ6����nw"æ�go'nb�{�6�ǋ�����_:��5�-��iM{5;���a��!�(�{h9"��w:`j�h��w&�hѰ����C��[խӑ#�W\s���V^F{W+F�n������n��%�fh��2�n��"�s04�%޼[yGRs�b]@v�ga7�pl��.�B�/s>������pY3q&r�Z(�g;;#��-E���A�dIc���ګ��
����s���Y�L�6cL���X�ʶ+m:(;��'@s��'DZ������mң�^�����T���6��ʒnV	W.���>{���X��u��o)-=w���k�M
W����;�8R���"WE��q��b�utd�\]�j��[���b%��>���X��X��+����&ʳ;�!���m@a�9�8��&VJ}�P����ܷB؛%��X,`�1'��Qt{����fxc�DEz*G[w1m4MZ} ��6�ػ����U�i�}֏k�2R��
L�%�(���bY�)hϒXM�;�P��G��ZJ@]����ֱ��]�У)��qVh�f,FW"�������kY����ų�bYۡ&V���/�>���'7u	�(5m�K�_n'w��Lve�|>��f��4,��!�h�Fc���n�)���8�T��1�]�*�.���������K��X�<�;pb�,�k����e�}�R�	��X3��6�?�c�z�Ю�	�7<J��\�]N
Ͷ�ۖ1/�� ��q�n��H!����ճ��x`xӠ�Qb=�[/Onһ��u�4b����+�A&����V�Y��"X�gu[��LR��9+�[��ܫPP��P͏�H��e�1�Y��]\I\0��d�,Su���6��ꊞ�b�����n5:mv�ʬ�x(�!:��e�{��#��o�yK�M�L�.g�u��n�̓iZf���o�M������).]��R[[L導d�Iw<�Yi�j�޽�9�ayY�D*��ε�:À	f�<p
��[�#�q��3���P@�������SJ�WJlC���F���6�ve��$���dJ@��tohd�ͭ�9uc;�j�Z"7f�����Q�o���+k�gC���,�k5��ۭ{��K�vj�ҝ���"\b�E�����8������> r�V񱝤��������q�r9���Y����]�/�Ch8�Ǚ]��V�α1q�ѐ��`H�2��.V��5�y�	�������+"�\[)�ry]x�c�V^7q� L�m�3�fY��0vގ*E{��W[��o>�t(p�r�,�ͮEK8�<�s{4��.6p�no�GxZ���V�"弰m�h�
Û�]{.���]vLj��C1�:�;}���\�n���QF�ռr�Wi-Q�t]d݄���S��[NGf>8�$u�z��k/a�x����-r��.-��>��m�y�-!�"[ ���9u�5���+�J:�Q���H��vp�,�O^��xf�oG��ɇ$U9r��k9��|��	)�f�D�xف��k�e�Mf��7��n�2��	�\Cr�\Ϯ�V�tI���E`�6�,.�3	������Q;�cw�B�!M�����¶ol�G}eL�"�M�q�a��5�g`��ʔ�HϥR��G�Nx��:pvo����Ė���v��6{��2Һ1����v����*t��j+�P+6h�l��>u���n(.���cu-�YA$V
�}���tW�����u��U@4W>����cl#�޳55��ՠNЏ&���q�[E���pa4��~6���|��F2�ә��j(M/��mr��ѐ�eV0 FŜ�ˢl��>u����<��X�:�@�K�b�b:��f+�(�^D �o��z,�����Į�ąiYn8bB.w���4���{���t��zS�>����++:V�LIrٗ�m�-,R,P���]b{.��܅[q�4��M�k��e�Yeԁc"wen,,�
E��{ԥ�0J�R�1x�)t�h����KŁ�-���YK�Z��00jpY�Ʒ.1���ʭ�/,VVG#�nf���}�R�ǝ�am�V2��rZ"n���W�s]�/��u��e�3
h)s*��}�	Bv�ݰ�Ɓ,�Z]u���*�r'�T3X�&��]�د���]{�fb8�f_T�"�ºS��F�h�o��$I��gssj}��Tt��tr��e�����3xGR��ʡB�*�5���op��k[t:P�f�Svj��i�6]����k:����yu_VQ3C�(h=���e�m�s��'�3�ʝ�g�!D�ιu5��U;�qB��N�C�Y�(��t-��i�:Uٸ]�tu�k5�c�{�֦T�o����^��& 3 ti�`*ٻ�Ht�)Q	b#Wkݬ�W����0e�W����:� �
�h�yruf}�t����Wi��\Y�U�仕in*j���H|��,�r�˧�v2Sъ�9i"���}j�L��ьB��ֹK��S��X,J��+u�������Щ�7����%��v����}ݖɲ�ƹ.A`v�:��|/^A%@V󿶐��H�S��/��}lֈc1��m�]C�
��l�n�w[�}�]ɣ*h�ʣ�U��W#����]9�aŗ׵/�L�qb�Kn�8�i>�&����]���OB�	���uX�6���om�z.�xx] (�
�8T�H y5�m�.ы(�����c[�<��nl,�1+�q��ap��i�h	��.���|z�ecr��̂���ˎ�n>\����f���Ѽo2��c�w-�I�
/B���d0�䭁�^	t)���=�1��6�����n��F�#}�V�
, qA�Z���Wb�� _����9�)�4]<���U��0�/BC�XWRk�tZ�N��\���N���4�3@�vԃ/�8`
�
y�����K�2���k��1F�z�L��F<(*v�5r�j4��}��n��-C�8�L��M]��R��fm `ĶZ���(#�࠷e�]��x'����x�ұ*b����O �����CU8)�ku�*Z�?B/_L��S���'vU�+�sz�UY�thX]��]�̾Qw`�w%�u���W>��^kĐ�kճ�`j���+~A�\q@dCx`t˴����5�:y���d=�Yr��D�t�
J��ʡD��
1+�o�y�_]c��0@�Y � �T0*G��i��s�kHU�4�"�$x���8�����!$��BI4��@�~�BI��d*@s|�ӆ�Q(�mi��X4�m��m�-$�%$�l��Mh��!�DY%��%S%Qd�M�L��غuc�.������L�a�Y�ܕ�O�j��o�̫������� ��p=ͼmJT ��ϙ[z��y#�k7Tvu�@!�_3�͒�\��)bŠ>5�t[:�3�+��Ǎ�.����8��,�&�)Ar7}	��B
�Rm9&��A��9��f�\�T\y�o�q6���+�m��q����Y�VL8\�`���1���sUe_lV��vL`"���j%������s��wQ�9<�w�e�d�bL{�u�w=���nN֧p5`���`���;�&kOc����e-[��bIY�o���J;͹'��QRC��5a����)��s��ݝ*"�]q��&��i�!ڲ%ۦc���t�)���$w2�Z��͉�x�b��W\��mn��]6�aŜ)� ԢA���3`�pF^���T������+��U���y�gf�q��#x{ME�"g\t�Z[�P�<G��F����n�(�R�鵇��GX�M,�9�݀oB��r��XS�S���x���P�N�'R66����1`6��&�i�Ɗ��R�7k�(0�M�:�=,F�a���gz���8]��^������p��A����JBf�W�c�w���^���ӝ"�;8&�"�D3y�`wL	���ך��μ��
�'VU��(��N)�-PIqv�
t�����*�:���^�V��-S�� �ןB��w��9}DA��cVkQP�0D�sY��[�zq.LG���L�����eپ��2�Q��wI��t��B�J�"a�gJ�f8q� B��z󢴥Q1�Pe�A��C��Ֆ�ݨ���� �r��é9x���|%4���:�]�&�+E�rQO�wV����/�l��Eu�L�S�u3E@çF.��N��
���@PE_Sb��b��T��$�|Z�'��b8+��QN���P���i*n�ѐ�5C_���z��X��@�܊��}V������ y�W��}���Ū�˿ӽh1�_O�}�̿aC<t*X���]zK�7��VW#�e�q+��
�o��󬱖sƼ ���Ԧ�`�qڃ@�GƝ/-�����-�����Sh����= C�U| �`�أ�^��۬�~Ά�Q@�L��E}x��*��Y���T0w��f�l�n��]��y������R]`��S^�2+Yj���-:||d�
i��C�%�k���{ֺn�~�� 
{��r�����Wc�A+
*p�~�"�gښ��ňŒLk����h`��D�bt���� Ì���ש�+9�Ly�2�G���g��ިFA`�(��=�kX�=���ٚ������b#"E(��F���*��F���Wq�0M�=���YX��р��m�e%n��q�Di� +��N'�L�m���5UV�-���:��b�#=��l�%�!���X�;[,�q
K��})��
�X��o�ܤ��ӊb�w̝JL�W��-�3
h<�����7�zHok��4�㞼�;Pԉ��o���E���:�5�x�A��{��@~6(t���}��;\����gZ,ze�&n��P�

�tCOyW�@��~�Q�4I�Vo�4��K*���<�+U�չމ�Z���^gs��ʾ��-Ǫ�L�(�)����b�w=���֡Zh��{h�G8g�e]�8q�}�Fk'���6޸c���ai����|8]�M
V��GN��X���XG�PT^��@�<e��ߎz�K�Ԫ@6�F�����+K�>�L�X^.:D�T�|�a�ONW���yr�d�}�o������GF�UZ��K���u�@h�X�N
�ߧ)g��<ߠ���������cW�%��"�>�U��`]׀�ݏ0�q"����f�!"�LA0@1�/|�ݛ��>�ep�M�ۿ<�ѯ_� ���!�7���E����6q�	��23�g�vV���{Ն�v�R*����}�]�ۛ��7a\,�'51�<e`�Eg9�)�p��HFc�0�ŝ�c��)X�r'��Coe\r'�eM�H\}D�8��D�d�}dK?�xw"���.���4}%m����QC����.�6Ӡ���<��ai�KOݞ��#/%Y����U}+*Tش��g;
�x�c�ΣWLe����u=/�P�?3o�{�4y?2cZmx@��O�u��\>����::��;��B��s���t}�0�A���!g��~�����5ǥ�[̚}�d�}����frk������5m%��v���;L�ҹ��Ȍ�W��Py���k��^\T�W��(h�bm��r$;�ɡ^x��yt�y�L�$��}�{3�X0��Z/؆���p8��.�t��*��o�W�߹HȢ�X)X��X��ADbc:�!2�"�)" ���޷���kX���Ţ���<��h~���v��}CҘ�4i�^�b͚�þ@S�Ƒ������Wc�^\^��R|C��1�@�@�ha�;�]w�V=� ��b�����]�\�>��X�D�v�d��L�z]�{ �j\��սl+W��N��8Q{��޲"i�B��:ins�ր@Kry��&�u������Q�z��.L��}�]��ȟ'������;��1ֱ�=�w=�*dߵ�h41���7.E��I�a�e	(Nܠz_��k.��z��U%L<��b����ɏ�a��D"0��3�g�5�]`�r,�\��|��zy�h��4)�S�t��{�]j��8� �U}C��W��M��A�4�OU�L�`��!�inu`z&��W�;ڸ�od����W�_*�]�il� P�ɝJ>�HQ�p���,\��>^��{��ׁ�=��'l=�^�ؿ ���[�_`˖�F�cA��,P��DS�ֱ0"��c~�wY��1{�O�nI�(��"� �2���w��V���5~����
�R=�6�l�Y�U��W�ˍ��l�=g�W���<���x��*��篙��G�̉�-���1UM�E����5��`a��@�`u�S�:�8��t�`�} �!����A
���:h})a2�|���}1`�A��_]�]YB�\�]ZO_`��I1����M��P�K)�6� �k��r͇ߤ4��Ѯ�U��ր�Ȭ��N�8��L��ТT>�b����x�+�4��Ă|���S�ɴ��x2�p	�<�6Ԩ��G��qN)K��|p@O��b
��V������},CI�A�X:�=՛�@��@`���O +I�H�T�D�LR^����. �K9zJ*�^p�z��k e��9�2��'դ�0�Φ8V>�R�����>����w/w$~��D*�n��b;��~�J��]�bG���d�{�r���ڵ�}޼
A�}�Ț6W6J���f�� x�?V����3YĽh�/@Y,��7|ޒ<j����,��O­r#�I=�o: eu�����g9;{#2��
0Y�T��X�X�SˋȞH�yKhל�C\����<>�i�a�VVz_ �P���B�ۥ ��z+Ś�L�&��Ǩ{0��a5��f�2����P��a�ò��3����L�uϽ\�F��wkP�b"����kG�,��:늞�#�Ȟ̓1� B�S���E���߸�:����*Q/4swӳ�+��d>��R��y�}ӫ(���,r��%�������<r	1�bYa�V�l�s������/ı�k�ޔ��0���u�4|xR
�5�]��趻��W$����������q���	 $��b�}��$�e�oNiǮ��| �EM�\��	;#=��������˦yp<+`<4����۩�����(`�����O-V��#�|J�-8`�X��ݤ��%�"R4 D3��#�u)��,�#+��f�RD�{j�cQ��n�p����K!�	�cL�¹����y&�v��2cD
#e9!����F��<_���+��Ĉ�b�*�AVE
*$d`���@QCr�]�K�g��󏼇S��1�49��K��w �0#@ "*�t���ʭR�,юV��.x/�
���+�s�h�K�g+qæ��i��-.4T�3(Os�sְ������Xv�s�����v7c
#u?+���'�~�ב ��[�*�OKoa��Y8�k�rY��u,<%�b^ʹ������׈��H&���:�fC#l��`� �`-��$�(��v襴��1DD�>�m�[L%`��/�L3��Wܢ�١@�Bj�u�ڈDXˡ.�,]��fte�a^�<��J���ߎT���P�-��Uu��y�E��@� �&\Dr�� 3���X�.�]�[�ߩ����Y��O,T�${εi�Ʀ�-������ة�1mM��^N��M�p�_
��s��W���8!�27��Ӌ*�P:�.7��#��?W���7JK�������99{�\�c��wv ����+�T��S]��r�J����G:;��Hw��d¶�u���ٳ�Ş�K�T���e.h`�DbH,E��b���Vs�ɘ���F$U;�w������4�U�Q�:��O�@�\�DN<�M���u
h^E��G�~|�?e����{�!���E�q��:|�٬�%q�ӷ�� �^Ҹ��������q�XEpNH�eL��E����$��~�It� �5��o�7����^{�yΙhLS|�Ñ�Mg�89�_�r�2x�$��ƍq��Ns�����=u�w�3*3����eu�+Qa�j{q���س��tҩ�,�S����H��PTs�����[k�^�o�8nwU��R���P��*�Uh>t���{�c�383ΞP�z�P�!��V=��k2����s�M�|���ΖU��xQ�.`�� L@b0Ԓg�ܸM�Zl˚sƟޗ��{�eŗʯR��: z�&�m9�DdK�T��!���`����]�䐻�%�LQ�;��6�$��!�e�w�d�si���>9�Q�Y"�;�� i����]WM����+�����Vqp��d���ץ��@U�U��h���Բ�g]����㨭H��3�RH����"�p�QFdQTX�c#�l���A",Ȑ���0Y%AE!$�b	 �}~��4���o1f(~�+��Xa�O��8� ٚz���o��,��� 47��^�_�$ճ��М�tFºV�$��4X;��.�;���k�6ǽhM+�Q�K)�`XY���M��x��]k}�¹=�q��46*ǹ��n�C	�g��b<�����Y~V���쨣�o-�@����)x@ޯ=�+�{�s�r��U(��r���wv�.y�V=���Ya�1b*�m�m	�\�B�#��k���#�T�q�N�L5�[��ƍ�M�_>�5�����@TQ�͍�x���G��iB�X�r�t��O\������ik���Z�Dܒ�<D��j��$)$��:.3\�E�2Z>?�
���BF2���g��:����G�/'�.��*�v_���i�[y�c =j�:���u�Ӝ�`D �D5�$K{.��[��[.�P䲼+�Y��n`B
��)�x���:�%3HQ�H},y	���]���5�`*[#��=�U���.�r+�S�VA\H
dD�`"��k>ǹ��l�!h� ��{��U,�?���,?(�E�VmMm`� n^N�J{�o�Z˴4d�=�A~�� (X����B}�%��`k�첂:v�S��d�#m����D
�B�����N(�����Z��SR��
���2�R�Z�(���ɶw��kGl՝��K��ت��dl�v���-J�u�ʧ�8�����fiz ��-��^ap�#� �)�8K��;�UN��L*����򕸴�wD_	�FKьU��'_!��ޑ� 	8���n����'K����*�7�:w�`]�� �.�kq�M�U����4���xlɶz��C��r�ݾꥷ'�'�� ��nl�Y��Ƅ�aܹxxW���S�m�%��t����Ka��;ON-��x�Ż��+��Ż��W+y�q<*����؋*�`��P���҉�=��Շ��8�+8����=����Le��)f�"B �*�)�*�9�%�@$B1 �kכ;�����=k{��o}���42�ڈ�bܪB��i�����~\"��T^�I�l�@Tf���#=C,����,A��.��0zJ���G�0(`ܗh��ӽ�t�;�]�� ;����W,F�
|�F|Zܬ�b�v:˭J[rU��/�bl����<�+�. 	ޒ���c�)GuimA� �6��xd0�䆪��Ο����jx��&LaƉjrv�F/f�f�c�e�<B
�U װHLq�7f��<ｙ櫖.=�xk:k�y�f�����z��� !@��3O
@�%\��X���%���2�
s=JG��)WB�0��jn��u�PT!@�5.��M�+��Yx�:5@�tN�kW-�&n	ǔ�|��G�2��e�G ���sM�ê��@P������l����#��x�D�~�uT�i͉wvs�|+!����e8jv�+R
��F�De`���9)�Z��
�N���rkT�}D�*�g�ң�����.�y�}��@�Sh�oe!�æ>͆�rU�f^��p�n�>y�J+��irA� 8TY!]	
��{�R�{Υ.��6O��k�Zt���V�v�*� B���{q�+v��׽&�1t�K��u�U���84+�W��cƫ��Y�Jq'���]�&��Gf�V�f�2�^���[�Z{��̬zw�]c�LSr�y� ��܃^�Z�hJ�U�KY動Քu��.P�:�j�����q*aB���6�[sf5�v/�I�.#"l�$�*���h��4� T�� �A�!�h�t�6C��B)��D�d:7t�!�k8�J�a*""g8�4�jKl�s`f�A�:���n�Q4�Գ� (^U�J�3��:�"]�5��v�B�Lv�7���_;x^���[(i���$[Qk�` �&*(
��h�/�F��b��Uq%}HEv�#�0���ha4,
lL�h߫-z[��0
�� ʉ,��ԙL�()ծ���W��Y�9��Ԯ��Ql�e�2��@�φ���R#z����yv��I��-f��-��>0���b%�,A��-��Ax1lCkn^� ��,�S��V���o�����z�ʹ�=�7Ӵ&���w�s�mo�2��6���!658f,I���[DU�h�y�&�Ε���(�SE՜P~§Ʒ��;%��s��l�Ր�.�8�[;��::�0j+�sL�;ל���h�f$�F�Q��-T!ރ[�b+u�� �S�V����񖳓���x���9������j�:�`���x�J�.�
ˍd�ڙv��sV&s7ѹ�2�֒��Һ�ָ�9�M/�j����<���rӴ1]�IZ�x��
��:����(( �M��A�u�M`�x��g��(��5%���έC���W�$���E�{RGx=�[6��:S�w9C�-����̋�!B�I��#w�n��+fą�L�W����K*�q�	9�&���M��ҺNp11���.����L&�܅9bW
���Ἱ�U�X3��r��;-�U��;U��r�96�x�I����#n������tӺ|[��C��F�t��� ��ޞ��T�h�z�a[��<3�0�f�f����S^\m�[N/,�x�q�ȧ��<����IޔN%�e�IL�4�u:�	�Ԗ�j�hn���T+��6�!�s��|�hpaO�l*�h��x��@�)��>f2S>H�u�[矊q�:��L望�Kp�;�`2�tO8`�ϱx`.�6��Xi y�V�p�ܡl�s�0�y��0�[��0�y%0�|�fS���}o�}�����e��h�M Ri�V��qC�PZy��2�o�~�́������%:J������Pg�KfRx�"A%S �Z�� � �M✠SL�|�zɷ����TX��T�0R"�]���(�XDC�u�}�}��^8�)H,8�KN'�dƪ�
u�Ʉ���KO�RG��!��Q->�BФXi>�-�C��Lv��Za�)��L)-�.~��L��b��J�ӕ��֥�c��ɔ�Jg�P��U2S�8Φ*�O�T��Y�a���3`a�N2ٖ��W]C��v�P9T,8�N9f���*[B�4�ٲa0��+u�}���o�����5�M�RS>I�a�;�!Xt��K�{�2�%!�P=��h�a�V
A�x�0�l����D�s4O9aڠXğr�!�ɢ8����ƈ��;>���u�m�Y'YO�	���"��I�a���'fS*�k�M��!\����I�
�d��
�M�0�y�wSI�-�a����[`,4�no���~�]�_��=��J`.�����2��ڽ�t���îYx�@�T��-��d�a`R#�$���i�%$�TY)�}���XS'P�5ʆ]�!<Q�@��F�_w$����]4�X��}�g-�Kgިo��e'���b��h���JB�枡�- ��u�K@�U�{�10�C�s�{f��b��e�"���Aw�r��mvn�,�"��FH@g�ႂ�Ч��pq%03�\�0��,�:���05Wt��hy�m�Aa�m�5�MHo4�dj�f{D�Ki`O��̋���j{����a�D@$`�^O�N�zM����u�^�JscrtW����lxbSLv����v�C�4%�����R���w[�_�N���IL�
M�����~�!�3��}����L������@Y5U��<��5)>g�'�Rr�XZN�g��[%&Sl��}�{�czZ�9U9�	�
�-�@�:��T�!8�Ԕ�h�I]���j�u��(a�q��a��F�ci�E �!�U=Ve�/�oh���ÿ��	n/��L6�M�D�1b*�"H�Ō�̡H|A��N��nu��-<��e0�5T�Ri_]d�y�n��2����&�|��O:a�T�m��_{ݗ�s�x���d����
]�8�����Ϭ>c��@�wg7ۇ�ZJf�A䖆�3�y^ѡ`,8Û��T<��S	��d�v���Y���%e�cZ��p�i:�٦��!ߨ��$�l�c�0�IHU,>I��1ۓL0�>O�A��B��v�-�-�3[�t��!:�����{���������L�I�L��g^y��;e��3��D�|�Hj��RB�wmNn�!��O6�1`a�aOS����M���Ae�gɆa�m01U'Y^�~�~�c��z�Hc�6̲.�I�ߘi��֓��|��|�a�_U�v�)�II�<���,˄$�-�IZ��@�u��a���`(�����(y��=�����:)�HZ�[�'�e��m��%�@��:�0�O̜p�Y����J��S�
`c���������f��)���DE���N�w�}yyZ!1dx����i�a�V�p-)!�ahRm�}��M��)���P)�
w��O S�<�&��ai2�6����c��u
M����}�x��z��-�wrɐ��-�p'�FP-��;�&X[>II�8���_�!���L��4!�hYL1tLz�8�O�Zγ�Zw�&0��): @�d�@�ߏ�ӯ�׺���[�4�5´H}_}y�@tQ%������{�:
#�i�u-'�6��c�aw20+_+�zM˺ô��qd.��F�s4ʫ�K�3X��g!SPn�J��j�\�N`K���s쁀��\)Y�a`5e]�6%t<^M�E�U-U#'� ���>�4��'b�Sw4�6��&Z|��d��	�,&�jÍ�U)���KJz�!�TOwU8�0�
A������
�H�",X�j0AUD"����� ���9����Lb�L)8����@�ױ��(R�uD������u�sXd��j#Q) QU���)��E`�B�M ���*5R���a%��������&�m�4���N_2[i9��g�I�h ݴ|G�$�bޝO~�쭘Aa�j��o��&R)�}��P[4��8�M!N���$�B�Im6�Il8Ͷ�d��ѶB���h�@S(q�s`�d��3�o{��wﱸcH�j!�|���0��oY�c�>�L��&,Xxɧ>B�B��Re+�{W���C��GD6�i;�Y1!
�Wɖ��Il>g��D�����C����0(�崠F1��6�a��~d>C	�}�8̠(}���$�n���0�
m�L-��_y�+z6��h����&v��:>��e�i����K8�N%?!�^7e�(~C0ϘS9u2�9e2Ri�K`���i!i��l6�aL��-�0�
�0��L%���������]���a����m�^H,�E���@>�a�y�{�N�
��o8���5!���;�wti�~�آk5-�C޻0��m���Q-"��|��R`"#*��)ٺ��X T�,��h�-�2���~�Jd�}��b��̶Ц,�@��xd0���آ7P5T{tw���I)2�z�i�6d�Iަ�t0W����j��=A~���s�g�&� 	(��q�hQ�s�l<�0�6�0�<�Wh��i ��$��;O�Ra��hSI�����@Rd�_�m����[��8p o��>�{|�z�@���i�9P�N4Ͼ��e�->e�|��L$���������~�:�@�L)5췖d�%�E�<�x�\$X���C,��w�뿣�ӺҠ�3DW�
�gQ�TEG:���iHV�2�l�f���(�B��ԖtL�Ut�!]O�T�aܹB���(�5f����/K�3����_ �@�]H������ƨ�p�TJO!)��\0�6�[%�����2ل�|������0a�!H{��$�$*��L��3vél�4b
E�PDPQb��
�f�RH�̴"�E"�ǽ�{���}
i���6����O���r��_O;�+���E+}�	��N8O��z��<Bж�_!��m��&~�)�B�۩>�����S�}�g��}�y_]�[@Yzɧ,)
C�����ZO�GP-2ɤ�T۔0�O�f����-�0FANUe�3I����n�wf��<���i4��2��u�]���W�l�r��N�<�i>�8�6��9�%��S'�I�,�,*�w�8ӆM&�A�2�m!�a�f�d�mZn�:�`�LY:�|Su����}�^^� I�	$#�fB�HL]�SǬ��b���w�vN>@�IL6��'��Ꭺ�X{���,��%%9��2Ͳq-'����L᮫�����<#�,�Q�|�O�[l�%>g34N��a�[��S/�-'��	�� �Za�T���KCL��JBЧ���C��i��C,)
K>=$�.B�k}���t�cL����[O$��}��Q2��4��䔇�[g7Rq)&����=�"ş$���i)�R�-�Aʀ�G� F�$p�D����sg����
O'Pj�,0�!���� V�^!O�>�?J�ݾ���*�}���ϵ���tH�x�"���A�،�~w���Oc�B��NL�'^��}Ә���^;���^��D���b��y�{r(��{��e��}`�D,cb�
���$b��[)Eb�b�
�f�k	ˮ����pݬ:�`�-%6#��((
>k�b��':�\r�Л2�U�aG|
yNgAy���W�K:}�a�ܱ�e��X��Ǔ��I��=�8�? �q�I�1����wƻ�_��a'��+LS��}�a�e�L!�ym�*������C�g���H���{䏀'\���>Z�X
_޿�
\��%�	�>*�Ǆp��uw�?K9��U-�TX�I��	��}=C+@�e�6���wǷә�7����¡�]�� 3e�ujf�t)Q��&5T����@f�2����f����?M�����Po�f�j�E�'O|��""߃ �$�d���d\5�����=�q���MaRX��T��nn��+���j�#����K�
��ώS+�k2 jds1�}�BStѭ>�3GNvO��,�H�cfل�ʾ{Qɞ�&���>��G�;0Ά3_:\XtmT�q���K'¬���ـ>����7V��K��ȝR�g��oL
S�}���T2Z��"��ܿs���[��iN�m��̢#�^�S"DX�Yo��h�~��9��{��Q�CQ"��RDTi�H�DEH�X�`��DR*"�#:o7��~��U�V�W9�j��U��k���H,$A ���9�_n� ��e��4�z�ׯ+I��I�����4h���c����yڪ@8G�l�9�HK�
添�^{���;-�H�=�ٱ�ߦ��78�i|nO"��z�>�N�"�zf1�mmaݩ tc�»�E���it {�����7I��Ȗ>}y�_�L�ΪV;!|����8}��[���.]Jq�d#��?b(��Tb��O�^�B�.���!�����@���7#���-�]�֗ٹt�w�ү}���Q~�ҐF(�� 	��)�����h���!�c��)�kf+z]G����fUR$`||τ����=��kJ�]����/	����>��%{;���yo�%�}yD��������ڬ&6:��eS..�!�����O( {�&=�G�H���e�ه��	���Ӏ��X���v�j��o.�Gډ���2�iM
�7��Vᰯ~�vЇ�ܝ���#H(��/;��`a,��/����k�DX��)�����jo�C��r�n�rϛ�C�k_D@� ~j�W����>g��OUD��$�� A�f.C2��n±E l�Dq
����rE�{$i��C�X뭎��u�:�.-���95H袡�ۣ���V54�����*X���.`�gʙ�i� ޫ(0k��9�`Ʈ��W	4	"ʘ��>4#�"%%o�#M�J��M*?`���|\��UɉC:gD:�&0qZ�=z�'�B=s17����#ۼg$�� �Vo1�;�6(Ԫ�F����걲��Y���ͩ�1�A=B��bt�[3'���:�����'m�Y�x���s��g������
��
��H� D� D}r�q�n��n�����ч$Ug����[𛔝�r�Pgʅ|�$��=RE�q�s�u��$w%��7��Y�s�O�:A��;��ӣ�{:Ot�|�jIO!� �:ٿo��:��yC��1�� n�^O��d^��}�r�F䠏H㎕S�{���g�X��5%I�d�>��x��X�rģ����Rc:���ȑ�����,g�{<�PI$��Ċڑr>��J��2�fD�^L3HI��=.V�N@��+]�"m�(]O���h�tơ��� ��ӹ�K\�4mx�A�ن8;�5�w���oɝP-��u�K�=�o�|�}0�a� Y����8�`i���tj�=Uj]xfg�_Y�nof<���	{X$y���K�ݲ�Ύz���4A\ѹrC�E 2��6�_��/ƍ=��%O�@��N�����k�^�ž���u���k+uݱC����g� ��!�΀"v7�}w\>4����0�>�瘗the���3q����*k�t`�˪�����n������Y��w����g�QR��"U�@���*��,��E�7����k��:���s�t#�dH�r�,U���"A��K��H(��}!w�F��ڷ�Ǜ�����4��s_��^$ ��U̦X�Q�7'��{��f ��8�� D}Y��ݎ,��Vr~��ʧ� f��|�[Wue�$�`���M��^����s
�l&�m5��+5}��}!W��7;=_`�Q�s��x�F�]�^��{.g#a�Mq��+�QMK�����@���CX�X�B!bdC�Ϳn���޾��s�7Y~��Ԣ�A� �F"GBD DG�_Y<��&�mc�s���~V{����Y�grXۙ����R�,�>5������Z��^E�FiV��@ϖ�T�r���ۥ�{o�^ק5}�_��w�8`�� .P���׾�(�ּ�nj�����Ya�+fg+׹y'7��g6I�ʔt�*��x�-����[�saJ\u�W�5����7�H�҂(͛�F�K�����E/�j��.K�/xn��b�\r�ݎ���]3��¾�ޑ&�d�]̸������
��S�n�~�#0��{K>�j|/=�����}R���q�f� !|"F�ݼd��bq�P�J{ٵA�UR��$��f�;��1[�͇evUF�CwL񁥫�s6!ʔ#z���OI`H�x��T��-��X�_�6r��}.�+����ɌK��"/�\��@��'�Zt�_j�h�'}�ב�Ǚ�+p��K����b&�"�Y�o$]Ӄ��!��W�ӭ{����jE���o���'V}2E�/r�[��L	F�� ߯� !���(�1c"����P���$
BP��IR�X����5��j��/.q��_D����� vf;������c�+j���&R��D�Y!�]�+�L���>{�U���Rt|�]��24�D�i�	-߮��.<"l�׵T��� �đU�OxSE��)�Y�������'sX�O�BZ0���=�?z]}{�6���(F�0�@ T�����~�]"�ˋ�L�t؉_K/W2���@��U�!V�t3�A�P��(�[Rnq�34D��5�q�1_n��U���\����L������F�?<%�7����Y0�t��~>�]�,��7�}���D "A ���ZG����}���Ը��|i��K�8�Vw �e@a+hӷ�v�v�=� �@Ւ{ʆ�0�߸Gr��ε�x�5:$Dh�R���]����c4�lO��VT��.L(�x�d��14������ 8�ﾃee�R3��w�~��Zd@���շxm���,T��}O�]s��d烚��o�E��<���0ުpJ�������"PB/���q}Z;*�DAPT��JХb����λ����Q�V���$� ����IL�}��+9��̐�*PMΌ
��Y���u��Q����Az�d=�F��ۨZl[�Hxd��l�!��;�"cy̋;���U�ݗ��тe?P������z�]u��Ǘ_ 0��}���i��Y���խW�E�u}���0X-�/-4���e�Vu/w<5�/�㖝M[s;`�xa�~�l'%gW,;�� i
�#�:��Ҝ�����X���Z5܉ji��Ƅ6;A�*sX�*m��Q�Z���f�`�"���ē[Mޫ@�߽JV�1h�z� �n����	ՀS�d�;�,�Ŝ�_$ڗ)!t�
8��K��ʼ�`r;�r�o�Piңy�@eȃ8�֌Eަ�䫦|!A]Lޒ�i8��5!���[�
m}�MK���R�Ү�&��b���)utv�a-
�)E�M1�B����!)�0�v(�gu���<�. �0Ně�5��AGD˸��S6ޛq����W���-f��:xr&�
�jL���X�#��悵ԥ@p�g3�\�<�:�ׇ)A�)[4��X�HFwV����VJr �6��Υ���ힹ�z:4���Y��xbÛ���2�����B���;�A,W[y2��7"�@�"�X9pʅԕ���e%o�
����x�)ka��XgX�t����s�*�5�U�e��1�6�'��L���5UV�}҈��1u.�Ah�KZ-�Xs=B!V���.���e�׀�8�'5fnթ	V�Z��$�\:��n�J�fd}-�A �ºXu[�]������"e�2�0
B�^�&lKZ�TU_�}:���4P���;21Er�`Ϥr��J�T�� 	�39�򕦣5X+4~= $�|�M��@�l�Q6�,�Im�m��I0��&��[`�>)��Qm4�!�A�(	�6 ��{�͙���ЕI�ϙ��f���3�[EhF�h+�5u�� �YC��I��G7a�5��T�(�>���Q/!�b�ܴ	�[��Z�U�;w�Uu�dD�2�M~��+�+�AIvcܱ)(����h�%�	a�X[��!��na���xS�mh29Z3[nd������F�]v���)d�����bͬ��|a��2�����`,�����N��u4!QΎ�f"Ժ�9�]�w7�����Vw8�d�RVv�T�-	�ܷk	$�yQY+	���H��|9���`��DSe�G-�`0B�c���yL&�A5�pS�W����Ǧw���9n�te9SECJ��Ub뽗R�Q��5ҭԸ�P�OJ��͌Z�ƍi�:��v�*�s��o]wj�1Q�'X��WW�J3��^\RWr\1��utv�Q̬Wq�i��2[4���7*oV�i�*�D��Z|�7�u2��g��ͦ�T�V�l���`]�۶P���>;N�MQ�b �j]^a��ѫ�
m�c�Ʋ���:�f7��߈�\�	V�Eњ���b7�.tnq�X5܇�s�r�����F�h��=&�2.�lٿ��|�L֡��ᔅ\�����J�[։ѕ�6�K�P�@�1S�9'�nu���ݥ,�dڒ�M6H�5�M*яN�*��m	zŜ.�ՆQ��E|RZ�!�!��
F�;��r4��h��̪�p(��656����ĸQ3kBr�V�43.�Ñ���0]gj�`Ya7s�eE���xU���r�6$d5�6D�'Ŷ�m��t�tW��s�X��&�%V�9�#�_�u��
�u��9�7ߗc�z�tC�B��|��C�3�m�jɔY=�Qj�����r5wv���ℝ}ݯ+u�=� 
0Qc�At�,�B�S�N=n�g�D�]��K|lJ���{t~]j�W9Ϭ�o= Z�ʪ��	��J|�f���O=pT��%L{r~�G�^�w���,�<��f ��(G���*�/t����<IR� ��jC�Zk���9&4'wH&jd�k�k_�O<{�')�/�@W��f�"<׽�yڬ��M�!�W�_���3BƜ����*�~`
#|��w�I�B�w�� %��1:<�~du��V�m��������>� ���o�b��~��7���aTF2Ab A�~�@�f����[2J��c:�>~ϧbs���ͱ��(��Ù��)C�X��jʿ:�j�F#�vz�����NWֲ������)}��� ���OזMou|�%vx]ec�#3��Ѱ�Y��5N����k�Ic��R�M*ۨ�Ϧ�s�~N�Mh^8��?g�w�����+3�W| A̾��׫V�(UDTAE�1"��,PR*UT������"+AEF
"����Ѭ�w�X�sw�j�PUEE�ED�"�Xi�DTU�9�EEE�F**��C5B�
s��}6�uæؼ�u<�gTǜ����N����
j�
r���Z�"��N(Н��u�
R��v�o.h�c�]��,����W�#����3��yֵ<!�#�wO�h���q�J�<��g3��/=XT<�$f��bA�\а,`�̦|<�2�"�K3�1j�{��gݞ�r�g��fO��)�&l���A��S����B�e�w=;\�u�H�,��u>���+Dչ�v1}����W�崝�I��: �0���*g��E:괟n������y�;��|���X� �b@E���UF
(p̈́��Q ŉ"E�#*7ש��|t��Xe�g���1��Φ��:�,C8�,�O"�4ط�=�@�1�c��W�K^�pg9�n��[0��F�tL�6��Oq�dQ���6�Jy�{}ݾ��s�|]�t�DDD����(qUi�q�xh�9�����׮���ݷ��G|��ˬ[(_c�Gs�����GC↔e�+�W�⢌�k����F�1� D്r�:%I�X("�3@���u�����ݿo��n��zN�P�AI"��~��1�pkX�K��Ba�յ�@2Ԩ�YlW��i��U��7F����=����I�m���Af�U��&T=� �;d/.G۰l.tr���gH0��WLzʲ�	"�,��wYFE���E0P�0���Իf�/##��+'��������}���/i��Md��G�o2� T	�<�>��n��=�O��1|��v~W�ֳ~�g�V�g���3y%U�{�4P����G	�g�|��+#7��=�ظĜ����t����c�����`L���*�1}�:�w4ۓix�w{����wS��lyE���w=��T���V"���D` �����m�/z�l��4tB�8��4���ۧlŵ�����}�C���/E�mH��A�rhF�s�E�~4�Bٱ�ו�"�ӛ	\�s������_�/U��"$n_�59��{=8X���}�5�����}��s�ba/*����l���P��"�șS��b�H�R��3��^z����ml�$H��ڎ\��k�G|����҉�"#���uDD�O���{�ܦ��Cu����9.e����S��[�6������Aa3X��V��V�f�m
Aa4��sx����kY�;7��o��wv�������DsJª�j�T��~7O�J3�)Qgk��������Ĥ�����ǃ��BW�b�='����n�3��D���c�~'�iB����Q��n�^���}W{����^��������ߖ��[�P3���Ӳk����C������bN�r)%�
�o�:�&*�<lVwJ�N��A?K�m)����w)��w��[��}�:�>>
�]�T�cx�;�,c���H�����ڕiܫ��	������b��X��dD�|>$y�E���}�A��T���Ľ1�/�#�(;�f��|���c�l�Y{ݼy�N$R3vbtN���Ȭ8�zj���6|F��_y��d�^�N]�\m�=�T�ʪ��C;s?;�\N3����r*�aH�6s>�b��ϑ���h���0T��q�*VY����ͫx�n�sykȫ�ײ����;@ *��(Ȍ%}!%w�����2V�O2kCFGE��s�\*\���'�7H�������:�̢���ܖ���<n�^#ub� Y�H�|�/���~�5FsCP>a	�ioSiw�c2ZH��m��SҤ+hW����i�j=�!˞�Cl�@�ZM��YLDѬ.96+�&�k3Z�/L3'�pޙ�Kĳ�a�`�ƀ̢P�O��jv`�_:U��N���T�A�� �&�������t�8"���UaB�N���N<#(N�,7���>��+ꪯ��O��owk���Oջnyo&�Q�r�5JO�uh�~�]x�5��XP�����=y��{w΃�0��N���u���I�O�R�mOվ���וFDH�A��2 0PF1H�~��aDQ�4�P��y�g��G=�qt��~�����X�ۗB<������D�8_���{��d�%�^�~��}�~[�9קo�4F��FOy
�mNٕ$�M����!�#�d\o�#�%�����.�b�U}f��V
����~�ɫ�o���g�5�:Ek��$}�1C������#��7^	�ԁsR뗳eͿO�ѮD�ۦ+�J�j�z����$�\'	�yRL�+�z��#S��WB��{��2��Ԭ�X�'k�yhCx�����~v����3:�cc}<�������ӵ$|s>dW�'1����y_�]�-=ƞ׹�^z�s����Qg� �"#���
�0`�H���5�����q�]ޝ���� �u8��TUS�!ʅ"��毡/?w"�n�'�{B��<� e��\&X2	�s�E�D�F5��vc\z�Sa�v������<<�t��Vc��ܿc8��YƏ<M�y�X��X�d+5|`��a����W|;��[���6�!�CZ��at���=D*���"��1gՋ���0�@;mˮ�^�\���ӵ��� i w]DD���n�N�U2�:r�ꯎ$�������ax:�.�1^�/M8]@h���V�����0�(ǰ��w�y��Dd���u�FP����!��i�Tw��O�b�͍����<�?F.�"�����'��=���XG�!3��x�b2�2uT���0���`�<{�t�,*ĳ}�[wGИ3�ձss �lOt�4l��r^]�;���$���Oꗆ7��`�0]�g�zt>� I�c�sfhֵV���J�mk�t1����!ۗPփ��4�m�Xc8\�HL.6��g�d��������v�mK����9��%�ԭE�_Up��W�DF���5:���a�#��#+s�&0�Lb���a9zױ��є=v B1р��J�пxߤ�)��ͩ��麾�TW��ۙ���{w��ޫ�k��-C�"��'ä��鄏��Q?P���N��+?.>��D#w�Nr��e2a�v�˽Ox�����ˏ1���*�Ɠ�Hc	;��!'�Z��� "��:�]�O>����(�A�bȊ�0EQY9�k����Z���3.�1O�QR�K����A)�y$h�.|ҫ��k�g�K��;�g����ګ��b�2'-L�hl�ra�U�=�#b���sk�����%K��`��8�#�$�Ώ5,��ѱT�^��:�H�~c�ɏzq��j��p/�_�N�tY�����&��k���U粣g���dY�c6e��5N}�ط�kv��^+ou��BG���"ȑV1�X�0��.T�Ǵ�ZW 0G��y�����O]����es�>:x[���'�G��������:84�E{����xh��sj|3˫ �TKr�ϝ]l�K#��U�*:-[����N�NY������N~����;��Z�a�����8V����c�T�j��~�N���
H��ԧ��u9������"�I���\+難�M��{��k&�;��-LO��&���oi�+��f,�Dk��WsDklSʴ��D#�4��fN�'ʾ%�4�_C3YB��
�e�ȼ�g����s�s�}ۯ{d���Qb(�(*"����(�b1Pb�^r^"��1E�����:�菔�%��9��a(f5��?�4��
�ļ���}���x�D�b�ī͍ߢ�Q�ۺŃ��/�&:���;����GϦٮseJ�3-P
�bMgN%��ݷ^&���Q:#Ds�>���ѝ�-��_��r�F)uH��"�t���_����8z��8+��=Eog���pD�}^��c�-��sħ2փ���>8���=⏳�]m��^�u�׵_b�ާ�A��DUE�H�������z'��H�8~�?xp4�y�k��^'FF�!�AZwb��5=31���_��(ר�X>�(wv�@���s��9ɨ�1L�@�s %��B�6a
�N����*���̟mVv�����;u�${*XjT��lD�}�Bp{���Mʯ]��-�F�)�X�J槶��"<�>�Xu;����$:�DP����)*0`��DQ���"���g�,ޕ��B���t� �EQsz��]�ݴ^*��uM�Hi���c�[��WGx7+���X�s�>��Ip�Z�lvOt��H��*�əb����g��r��t�7�:�h�f	XF�� Zg.�.��y��q"��A6,��@!o�o��;
j'G9U~���=��s]38���#�@]�Y�m��g���aK'�P�{ӷ�ln�P� ����%��ȱ�C�7-K�7So����0��R1�ܘ�0$aq=�3���Nt���=��=Z���Iׄ(�>����H)L��9���h��ϣ�E�_b�gQ�Nz����a�$��$B�]b���⍘��
p��:0!#lĮ���վ�s<k���zv�?v�#� ����N�Ȥr�~��g^�>�k��O´�ى1��7�W1��6m�����"v���@�鹐�'7 .`��U����oU�O�s�Ȩ|��ww�/\�͵�}9�֊^�]�?�,�@xhl��p�2;Ě@V*��4�Ŀ"��6l��ɔ���}��Lƪ����w�}�2�;�7�GC1���*�-_;�.�.��:���X��^���R�8�BL0U��,�}$#�����<���v@�H��F( (,"�T`�@R�����יֱ�w�裸(iQAA�Bm�A@��s���n��N权�H���f�^�ݽ=�3���ĺI��s%�lc+%h���e�f��νc���HG��ڭ�Ѳ8���RZ����dUQ����;��͝,��v�4�9.�$����w�&�������{�ffn�}��]�N�dN�d�T�r,�\g�祂�u�/z �F�yYy�H�0!h�����7u�Ǣ�aX�œ��= :Q�Zb�bi5��9�ӫ�տ�`|0Wx�����D@����\-^>=�������t ��i!kn�wv��{�=F���[ۺt�A�	g�mHf4R�ļ�U�4���{��MesCAҖ���ų�¼$�����5��Cü*��D}��vg ]�Y[S,�<m���������Q��DѨ�[���' ;�u����<O�2ҳ<��J�_����g�;���%
|P�$�7�@!�=;�\�=fk�`�FAdDcDEAL0�"
�3yw�o8��w�� �  �DG.;��s��o�C��:m���E�#���w'�B��*� TSq�����'5�E�\��׸L!h(��=�P.��B(y��	�"��	�f�'���d9���кM��U*"�L�Hn�5���"�}A9�2|���� �� ���ύN��e�;�U��>�n��L�B�������uR�m�YW���(3���ֆq���k��j=�g6�^��8M%L���C(�2ƢDYtgi�=1%�l���D��+�8�HNu�zݕwN�dFl:4@�3�*��8jb�;u�*�U�x6�X8j���
��t�_b�7�2�]G��rV�*���V0�X��ys��@�k
'㽡`����	���w ֝��=�X�P�	�u�!3���,&�.���w%>D�F�)]��u���r�4�;�{�Cw5k&rn�:��(S����F���IDG݇�^i�����u�:��sZ�au�nt�:�}�gyd�j�&�[��*eS��\~b	&	F7Y�q�s,a�0ܖ�ع*��R��4V����g.���*QiZkK�����dyԉ�,D2�q�I�.D�T>�"�����JA�:T�{�'a��w<;�E|����j�u��fc¦cV\��:�*��㠨`� ���7�42% I�I���C�Փ)�0��SG/�J`��4"@@�J���%� ���e����F��H�ℋ�ˢ2=�P�@S�d��Ѷ�a�	W[e��C���8�����j=�Oa�I�k�.����^�ԁ]9�Mlƥ�r�N�>}i�TJ^mJ{Zi������ͷ��o*����ۭr*�Y2᫾�4R`��w ��-J�u��k��*f����`s��i����I�}S �@�	������Y��ہ\�H]�Ov��
�{�I���"��d`�鐭�C�,E���ɫs��7#�EnP��=�ز��W�B	�*��[CI�c8�ߥ]���S�2,P�}ŝ�̩��Hn^wm����E�湥3�*�j9Phcm%��m��Ƀ�us�:����~6�[Ww6�뭋��������b�+�%s͔6�^ͤ�m+Z�+ٹXz�'Wpi�w����q�ʽK�g��C���^ƥ]���}�
�d
���Q��9O̗�v~u]AB�<��Ke�=�ɽ��������tEgv�i�|�Ψ�ά*��n�}�������'"�Ӓ�(�v�6��eH�t;rìR+Ovd�Ջe�Pz�keJ�c�Fٺ�@�&�Ĵwˍ��츧pV�M��B/bf�o3�-���+�r�tκ���O�9LZ�[��T���^��˴SxM�<q&aԯ���s�s�t�D�\�T��kKN����K��A���+��������6��yEO5���jΈ��\�eW��π��S,��-��xЁd� i��O�4�;�<�ٷ�}
�`P̓^)FǢ����Q,+���$+�HPz�8�r�G�άsr��H�I�إ���op̝������~�UOS�6k��<��}#n�s����$�f]���������"j:�k���*O[2�u8���Dh���KRQ���8� NֺW�������o��eئ#��@�zs��i%�L�|���B2o��Z,��D
�����n��Y-ŝ/5�h[+:���P8��3�5DEǱUgyk��&�g�X�0
��]'L��	�9~T�M���)��o��yZ��@c`ě�X$e�*0N��t�;�pڽL.>����V�����dU����U�X
0E������f�t��Xxe�.������E�=媖������{�2w�ɇE�M�wgĥ.��k���Ӷ����, ��)��aÍy�q]ҽ�ݍ0 � 	01( M�{i:����b��QY��V�l#��Mrٶ)<�'V��v�������z1�FaX�')H���׽={�bj�����;F��yI���`���#D, �{k1������~[�bHw�E{�u�+��*
}/����<;�a��iV�Ҿ�Ԯjw7j���=p]��Hn�S*p�S�b�'�2�Dm��>�
������+��MmH��FI�޵��縭�o�N���4*��Mg|�� �ͨ� n�珬לo}{'E�Ӟ�Ǡ�п��K~�gGúS�h�Q��j��G�]*�����?�c��0��<w���S�X�~�@��ﾭ��}�&G;J�0#yKS?<�fv��^����L9���X�lJj'�����9�m��W�7�*�/ �{���~�jfa�K.<8������������w�B>��J�%N���հ�E �D@I�%F(
"Ѭo��Ϣ��[4�����#vbq��"�k�l��2�têU��b�e4TP^��T�ܓ�".�{�_:��_�='�V�jy�߫��;�wS���)$ˤ��M�O37���F\�4`i�@G4M���m� eLEܲ�W5x�dF��v�wmgBC��b�M)F���&��'l�����K���&���(0.��gv���n��ԥb[O2r�9�vrS[9N��d�.
$$0s�O�|\*�#�g*k��3�Sf2H�?sFZb��%O��i���#�$]t�ݱ��UlJy�Z1�
��F�~�]�z䜔=';'��zEuǪ'�D�z�eku�>�5�d�?��H0"/�D >����~� �kFt��� o�>�������m=������]�|O|Bu{�����0��81��]><���0i�<k�T��G㧼Q�>C������[Tj%�!��lr�[jr���ˎ��3���~����E�ݧ�>VEJF����:����`/_�`���k���
,����&�x�Չ�bd�Y]|�	 ���"(1AbFb�X���\��^��Ys�R
H�Ȩ1�Pō^qN~��o����������>��x|Q�S���ى�j����Տ�8|���A�n,�!�����^ީ����q������z�n�֝ݪ����pO9�k��w�t]$" N�z�_�6�M������^	����0�L
`{�˻ӎ����V��Rn������F��&����GB�3u
Σ#t�#*�	Ci#����u�rΏ�u�xeܮ(Z� >�Rb��K���a�q:*�Ё*b�=�#e�g������������䎤����*�7Z ��S{
��/5(WN?z��>����R2Da���wqi{+Ս�1�q׆D<,�h��z�xƎ��w)��xG�nFA�����
��b���˻��y�%_��&>��k�o��֏�����ܠl���fק(U�O���G7 ��xж�p���tC4(�}GA�Hv��<���mF��Y�����>���=O�z�T���c���A@U�`
����R)~j ��u��Ս{#��yUϯUxVb<˙+��U��1^f�T���l	"G��Ёx�9�}���_����g\�s7�Ϥ*���9��X����P�p#�1ӓ=I���5΀B�Ǎ�P����rdЋb��xyh�ћ��!�q�Kҏ� A�Hv�oT����_��-w@)�,5�%y.4������s��{9L���lx��2r� ���9I�j�����-��F�V����mN��Ye�胴Y(��yOC!~P25��:ה0�f��(tl�MJ����[�8�D����F��ٓ��ξ{���Ό-�/��
��3靼��m�Y����w��ov��A��Dd�"�}��������}�L��Ҳ�[X�#Fݷٹ�����d�HU/a���M��	�U��pA_M�w��r��=���A���\��T�+�[�ze����o͉��
��^�{�b�>�N�Wۇ��qz ��,2xšn�\E�];e:-����G��CX3�r#�w��f��z��O�\����y���ܶ�~�e�-�49׍ �MOx��|S�7$��@h#��B ȰU"�7�5X�����dX�� ��b �O���������u��گ>,堶���i'�
1����V�z�c��9�W�������57N��Lۣ�ȹ��聧3E�S K0�K:{���}�ݟ?o�\��C���?��i0o��خ��2=���y�l�x2���~�3�k\���m��+��*�aŊ�*c�ژ�3�%/�.�����"8�M��}G쩳v���hōH�~�հ�j��������=7dGd�)sI}Q�X�ʙ�\���g�s�j��3I��vi�*�-��2�n�6/�F��K7Ju�C} b Ɔ3M��=S^��1�]P�y��U�����5҄Kn�)�:a��8�k�k��Nc\� ���|D��p�y�Y]��m3Q=2����f�S�����:G<���s�N����툀8�Eޜ>u'_>�ه��zj]���6Z:TO^,OF�Nfh��E�Xt?d��7会O��__]}�ff!��A_�/WZ�&�7:PE�H�  @ ��"�b�D����)��bA�����:������Y�W�
�#2���Z� ��b�z���_�&�Uq��cQ�~�s����^��/19W�J�oW�R�UhЃ-{�
C���1�p���L��LL2>���K�ｯ����~]�3Ǆ����]���*X��E/�r���'���l�_x��Ԥ^��:,`��F�'�8z��AG�������WVbz/&}rvH]���|��*���}��O��׏�݀ �}� g9͋׿s�AX�z�qT-PR�
�H�"1Db8�X�Tc��DX�Tz���f��^q��\��9��])DV0X���A_���:�,�.���L�2�Y���ag1t�����'k��|�N�H.�\��:D��W�S�<k0��v�P�u����\�rj��J�{����)�0��]�'��PB��b����٫:UB�I���\�S�Q��݁���fa>e;��lj5�����'j�#M�ø����-�\[�ҽ��_f_��N�����*��/�l[���Ň0E���e׭�ա������L�����c2����c?��j<�[x������Z�1d�)�tJ�(�Q�'N�����u_S����Eb��)b(0��[�*"�w=�����~Un��ﯭ�域~-�$��I-����_v��{t:����@Y{�����J7��p:vh8� 1����B�H�,k��d��q��̬Ͳ�F��u�rc/�!��ɺ`v�&b�bg��֟'+K�C�%�.`T�~jw��斺0X#y�z���D��Y�mry�H�V�̛j�#��8����?�Hr+)]@�~^�S,�vEN�>�t�$AS�f;�t�<�} נ� ��I�7\�Sr������U(Ւ����2~� [�wk��[7�<<`iu��x�$�(�j��}��ʁ#��;�G|���L��%�8��yv3���]�e��7�lS�^�y�p}��hlSus��C�����]����脜ǰ�26rE�R��}�:����a �Y����*�Z����>q*{k��k���YZ�yO�������f�a��E�|�����-u,�`^���sB�(��9�Zjz��糽[���� D�B1?}�� �U�E�:|�$@(N�_���_��<ܶ9m
�G�ב����;�;귔�ix����L��������<�Ӷ���a���r��a����K�����V���e$iZx��G��ﾃ�߇d5S2�����s�7��nN��N��c�өƯd�����uLOc��B_pf��?��w���Ɖ�����O���`� ��(�*�(���J@��U�UO���4�Yp�R�ؓ
���P��i�nn	�?��ts����x�їb0<߇��yz" �{,�X�o�ܟf>@ H�����u_UJ�*\a����7��j�G�Β�4`ΰ�.O��y�ي��������ơos&"�&8\���Ϻ��/����Յ�6	�HƢ����>��	au�}�ob�?bV�}�X1|S��Z�Xݻ�?/PQ���e�d��y!wz���o��PY�;��*�Nt��w�PQ��,Qb�0]׮0�
TY
��>]x���N{���QA�I���w�]_��W���b�"�Dݲ����D��p�tz�h�ճ�2�nEB��s���5u���Π�ݪWV�FY ҟ={�'��qm��*{��բ{���脯=�U�������p�^.ٺ���:������'�:�8Zo����[��9��Y�+�ʽ��=wn&�(ތ|0(���I�[T��}DG���ﯵ۫�o�z:�g�>]�;�F�u||�2;��2]�6z��u�����#�x�+~v�����Y\�yg�z]�D I��dz����6�
�>����#��*[y�O]˱ee��mW
��ƹ#�*]��^>@+9'4�kW�j�"Q��LF�5��H�3y|߽?G��G��:�S�)�W-	8O�S�v�m����ڍ���^��*�7��x9O�WR>��r��AG�y>�I+���ŵ��_Mjߟ�*>�UW�80�W�@�����}Y����& ���+(���E��X_>�Lc"�$�����=� E�nK��ڵ�n�S+a���Yϔ�x��3��N�@����
Z	���wK�=^~��o� �,8+Z�7/r��v���FN�݌�ލok����:�Yf���6Ug�ƪ}�uz��)nbQ�)�<���lڳ�:+��!�FO��Y�Wq���l8���� d��"
1D=�ߦ{�{�w�_����T�u�����m���޽��}K�.���{ܕ���]�u�0�u��kp�T�c��.���ͺ�~�c����]W�^��1����+�u��h�
�O2�h*y��yeeϽBRC,�u�)D��h�����ym��q�]aw	�pN�g����ef^��H��Wz�7�w�24V�kquvڔ>�n���53�*�y�g�ZJ�9u�*�#+�oʱ@.�]5H*�#�7u.���j�*��Zj*]l5��E"�#I��33RW�����UkEs�a�:E �'��őS���[��h���A;�W��+�,e݊�FUm�a97�����Z��v�X>���R�������/옾�
��!��V�5�VPX�8����S̈́��T[V��4�i�X�Q>�)�mV*����T�7TɠS�}�;��Y�)�XA�%r3�ǦԸ���u���D&'eB;.P��ާv(4&f�F@-��+i��G���݉�J��O0�e�Z��~	�)�+ ��aΠ�K�E=F3�tq��ۚL���Mu��B�X���T�)���H���UU��ٜP�}�o5j��+�IE]ݣc��[V3�K�PJ�"�A�5��dg��e�D�d0�
&E�D�5�0ɉ4���¡�dJ��!�r̷Xԅh%Ѿ�ID;���w��Yy���(w+��wk${��q�w,�[�ʬ�d�)���P�٫�$:Nӽ(s�	P�6T��)�U*��Sᛘ�-�}�ΐK*�ΥUAT!���D|]-�c,i�u��,L}¯G�y%�.�F
��Ruv�\�kjECg	�#��z�X���D$�,!Vi Z�I���m��iSI6�m��m��!0�i��4�4�t�A�)J�� ��F��1�	:U�ۈ���̇V���C�:Imxv;;�T�B��"Ҵ;j�NSti��/h]
ٙ}�����K [if<�^��۬�]W;���j���穇�&N13pW�T�T鹴,r5�'�)j�8v�;�S:��3��$16
C��q��.�1�}ͺ���-/kE�E
���!������&ΗV����Q�Z*r�N�"��ő:5��.gv�8��Z2K�h!K��r�]͎:S�[��I�b ��J׷�+U�i��r�9+rK����&�u��h��'m\�9�!a���X_w�']m=R�e.W�R�0h�'>:�y��LM��v���fϝ�K�<Bj�&CGy��ƻ:�;m��J0�P�6Z8s�Hy�>�-l�.Y��j��,����q��G�#���G'i�Sx���T�T����N�5�nV��Օ��U�(52A�j�r��.���O��V�t�`��¥� �n�X78iZ��KR���8�N����z���Ӣ�9�i��x�l@xP�+��%��;N���S��J*�فP5��'�hwQ́.��ʩX��XвH�D�\Fъ��н�q.#M�j0��Ǆɦ�C�Xw��(��m[v�WS�Gz�R��[��Bh��Ҡ/3y,�zw�dZ6���P9��G���Zaܺ�qD�*>g���f�)�>�� ]jj��J�u�	��w�:
��d�`:���v�P�9XD&#�q]K["�V�����;cڌWpx��K4)ZJ�+VV��@;��D�A�I�S, �-�QM0�4��.��doV$��S`�����iv<:A��j�W:-n]d��)�e0&�v�F1J�;0#��F�i����<�/]`lR��y�\7�}�\�Ad��M�))Ц�V5�z�6
H�ӭ7M�z^Oٙ��?�-�����SY9��p0y�Ϛ���y����}�y��O������r�i�Y2|>�+��B�����Z��,�H�`�Db*��K"AE	-W|c�u��v�g|�|�;��7\�)_JL+{�El��n�g�'�z��f�W=�RX�g?84�!����{��7��s�F��"�<�� �r�/1ɮg�����.��o�Uu�Kl.[ӡ?Tv۬�Wp���gBb���i�ޘ�];�.��2����}`O�0T���|������K�s:
]&���sw/uG�?1�:IC��s�1�u��:�o�} ���^X�c#%a��� Qu���9�[��~c����k��8�b"#UW��fz�3h���'
]���(�<�{}ANЎ�R ��� D�}$�����[���(���)]Y��X��zI����ꩫ��:�h�ݤw�h�K[f��%*;�M=�a�-䞵��0ܛ����{�w���l�c�������zǱ�i���F1AE��*6�C�P�DFDX�]�������>�ڝ��A@�#����n c���s_?N8��w�y��'`�����a/�Fc�Z�q�ey�/�*F2�/������'Og7�:;_H����7o���ᙸ^��cC�=����֤OZ��>��O���ҧ%V�mf��T�P��x)v�ε���γ`ﻷ��+Gޟ5�I)�aoR�Qneo�y�_u�ns#Ih�ķ���[�=�c��u�O������`:V����ۗ��p}��'�/t�����V�H�^��1�">�J�C>���%^���Պ�zh��]c=´���w����.Q���Y��=��
g�{v">�O��c:���Ѽ��4���r�ɫ��
��=Y�$RcװI]V^VVaP� YqJ�7'���I�Ұ�\s"���͚f`�y:�)p<�Ch�krtH��r�߾�w���>��؂FX$`�Z�!���{�c��K�}����1"+*�U�Nh ��j�����P�ص�����N�=w�Er��R��u����5�}K�}��$쬼����M�>��W��P/AN:G�B"ZO���R�z�+b��b���e�ϧˉu�2eW4U�	lcPʾ�e��|�Sf�^'�6b�̧,U|=��N��W�OS�1��j7*3��=�c�s�wm�M)DAI �n�G�%�S�;��;�\�Lŵ2� �.3qϜ�^��.�OŽrS�}5��>�6�g�$vrMǽ^N-��#ްǺW�;�*�ꌇC������ݟy��ϸ�����y5�V?��ݚ���E�蒢Y��n_>�wUO1�wwo���7]�/j��+[3�;��|�}� ��"�l�`©A@Y"�hA`�)�LEUA'K�}���k���u�e��"ӔP�V�}P�Ev�Q�;�c��ư{i����,I�n��4�N���,����c4A����|��ɽ�;o�r��]�oZ���r�E>��é�-���D����\��aO-�(�~zwW�z*�gjk^f�'��v[^δ�{p̹;�y��x����+��g���U�)��퉥���Z/�@���K����~Ж�;ov����^t�D��wc�v�F�#Y�EJ����;}�z�9Y�ٽ5��N�^wg�8iT�Ξ����a�K��"D}�'{��	B��뻹�f��9y79\.z���G��C2k�<�a����������:<��?���]OL��צ??{�l7�%V�.^�����/���>\u���'{잨�W�ڣ���5���Z�N�_�أޙ"��A���)��Va�ӵ���sS��W��%��"	$A$�d"���oݸL+#d���gj�쯔���{�舀9�_��0�<^������v�����>o[��o�u�9kU��]fY2���$��L�H��;
��j�.��z�/�,����ܱQ����V1ĬO/�t�u�f���H��0���nS!滫�s5�w\��Pa�B�Z�Uu����#4�c���0醚x6̼U�S`W.W�}����}�{�셾b,4���:Cw*���ȻY�{o��w^��ߴ;X�`}V���|%�)�;�'v�b�8�^I�o݆����X�جG������ou"�.���fʬ�<�ۮ�5��=^ES��m\y^tû<�P���}�����"�@e69�������7x�ߤ��x�<�%]p��������V惶=��Oۮ����2��1ӣTW5��p�T7��]50v�t�DD,��Yc�7���'�}�+q������Ϣo:�}Qʧ�u�Z�?r�y8�=��Y�ե��g����'�	�b��oZه�cw�}��|�ߖ:p�0"���%)QJ$�B�"��w~��s?W�HRP�DQX,dTE�U�(�4"*��DX�A�DF t��s��|e���ۘ�e�{*�#���>�u�c����u@a�ګ�yzý������(�0$�mm׆�^�1��z�[�忞�Kp;皥B�N���#CS���:{�,��U��amqa��sZ�F-�����w!g��j���~�=DEn��Y����/�u�eyLx�=��0Yx2��֧Ϟfo�{ݙ���_�9����!߀�����-w���*/ء~�e�}+x}�s��� i������z��t�
�\�$8����]��BY{�W�x���u�W���j'N�)��Y2hc��é��5xW�����A<sTk�s�I�B60Q^"��Q%"L]mZ-��O�nc���}��!Hɬ[g�ū -y����λ�����1Z:���eeCܛ�9���AK���l똩 a���U�(�(�P���0�nX
 �$�b(�,bA�2DA/��s6���޼Q��ͭ��-r�9P+we�W��q�>�.�m{�v��{��Ok=߯�W}�}ko���F!����Լ�Y�bȉ1ύP��>�n�G3�2l�:��帵~�8�؊n���S}���Y=���^̘V�smZ��|� -�oꪥ;r�F�}����/$��COs�WGz���
o>�ݍnz�{��8d�b^=��5��l�<^ek��旫wX��{��X�x��DG>��"GI�3��yG��}�������Ԕ�j��0ׄwBZ0V/�ot�(�k�_���tmNq��=y���\LӵUZ�����ַ�l���������돣�.��Ɵ��׾�Rk���ϖ����N��ѱ����q����暑�:`�7��c�~�����[�^��g��6�X��,�
��)[�j>JT�9�g��5i�"��M׍/��P* � ��#'} P3�����to��o��1�J�=��u��ꀧ��a��~�̗�v2��_z�r5��8\�8��`c-+�5��s}��g �Z��<�⚘���c:���E}  ��g2J�o(�ɤO @LT������N�9u�svsN���\�s}��+W^���A+��ӛ��H�`�/Ǫ���r�:�O�����g��bn�ގ�z�4���*�x����[���L�"o'*ow
��o�r�c�(�s�>��~r�7-�G��}����A���	`�s��b�����;�4�el��]��Z�����7뼔[��vM����Щm��Yzi��k��5���ߡ)髑]�����y�l0����W_�c�n[J1�nq��1��ߪ����q�J��Z�b��'gW]}ݾ���{����Bi�L���.��%�nMC�1����<�E+ݔ�WW߭�I$̫&X��#���H�+������ٽ����ǻ��>ω�$P���#F�֑�A ��f��g���e-�����9����S�q�]2�w*����v�<��n�:e]��,��>������գ�興���Ƕ�c�����^�Ҟ;̇����=�{'js[2_���"$X�)�]��.�93�fB���a	���h�D��!�D2�.�T�MA���QԻ����-�� LgL��:����sW;�m%���h���W�/0դ�R��2W[Ȱ�"��ڹ�c�%����K&�\y�	ҵ�im����A��"��;�w^��M�3f�~�Q��S��7rc����cظ�=�ike���7���V�ݕ	l(����������|һeh:��U�Ej�Z1�k�7��j��ީfI�.g+��2�u�~���q����x\�B�ҍ�Z�S�H8���~|�,g9l�OB�8�L~����n����+���EP���LNS�ɿ-�w��S��}�K&8;���\NTj<��S�3߳�d ���S0UDET���`)�����9潗��W�Yn����G�m0��%���ۓP؇�< �P���~�l8�E�Gu,�)���9�42��߷p�b���d�������ﾛ����ĸU�T�lSv�N}�^'+h�����g0Ҹ{W�=R��aUg�:p}\�x�0� .Hk�%Lؽ�r��h���0��"�@�sO�ɕi��V��V>5�9p"Μ�(%���̫\}Lt��$�w���1�8?	�;R�+�f�����u�{����d`��#B,E�c��9q�z`5�n+����|v6��d�	W�b�:�9�k}�Y���G�ؒ���=;��/�E>��E�Z{�OC�z#�y�5�>S��LlfGf�{c#t��؄9���`ĥ����O* ��%�8P�;|��lZ�_q�y� )"���/���¢�X�&=}3��k�ן_=�}z��PXLfBs��p����{�����?����3���-��Oe��$n]|}�:�Ŋ�O?O~h&5��a�8ڍ���r6���fe�M�fg��̌m$gwb�ڈ�������]]~�����F�ъ��<��V{N�j�>i�#�3Q�2^[�G')Vh�J����g�;���:�i�����"z��OR�2��)Z�ޭ6�AcV��o��NW��u�ڦ*P0*�X3�+�����_e�V�R��u �yI�'�3µ��rǭ`�]az�	�R󒞚�ޤ >���g�^���(��T����f��3�r/={��#5҆�\���Lmۧ�٤�A%H������$h��`��D-��^�u��Po��](W���H���Fqb���,�=
m]�)6`_�@Ԭ$�����.El@$-PƏN�VL�R�U]�S9|�&�h�Ԑ�+7�D޹3f��<�N k[�<1�
����@�MRPI�H�@� �~AV�Ӆ���IHP�,נ��68
��]*�L$Q �+T�K�ϖ���3�8�20 8��Fzr��n�g.~\_ ���M��ct��	ثlB�{_���]����jۙz=�4mM�k�z0|�y.�~�q\9R�>�Z�����Kw^�n�x��v���h�]�-������3�F�͛W1�%X�R��l�5�d�>�B�`9� �)�z�L�y�@�G�-�m�2)���-Xb��.d��j�KxS(:�����km�*��%.���1�^3�B�貐Qee":�C}y���ޭ�.�3�bQ���&�ώ�!D��Լ��G����`}�ܡ�R�7ۏ�Z��5�hy١1�����;�#�q��MR�c�f�Z�L�0a���.�UJ7Z���u���:��ؕ F��F���^;��n<�FZ�EIHK7T��R���i^���u�ký7/(����	���_k�F�	4��Z�Q���_���=�}T̕��V{�F��c$,\4�ڒMg�X���0J���@��ۧb�WJ�\��Qv���F������_oS���Sv�v�P��.��Pm^��qZv�\�w��|��C8�05K6f>��&��C3)�۬=r��3&f�*b�4�oJ��|"�̌�0k����n�V��6NϷ-�V+��~���v:���[�qM�'i}�\.�D�2g^nm�}¤1��\���h]
�ia�D���Xȍ#t������z)jt^�9�h)�;o��K�r;.�ř�h�� w��"t��,Q��rF���vE����'�{@î�m��ݹ������v؄-L���9;����t��&�&���J+��[ٻG�͆���3�aOOfqK�M`Ú�׏v:��+*�~]\��	C�4Vp3�8���J��.�K�ur�{�\�ow�J�rkK�ָ6Wi���Vs�l�6ukW��ˑف��==��ɻ����mnmL�!üg5A>쌬pGz��hN�т�7��?�ҷ���Kn�<�̻�2\�'�ǮS|*\��w[Μ�k:�6���˛�\xQ��8-��:Y�uܸ�i#�rW)�S�u��ZoR�:m�#w��c�q֗�o�y�pmZ@�\b����O?�q�-������ۇ3��S�����c���9��u�}�|���>\�r���*�?`�~�fR��֞I��2�x6<x|����}Q	��t�׋N<��ӎ��D-��v��l�r���1�}�;��O��\=��|���r8	����z�ۨ�F��%>���6�مk;<w�����?g{�;��f"#UQb���	X+
��bLQJ�H����ꪅV��O��K6�������]p�Nn�{���>�_���cR�s���\3�F����{�螓p<�^.F���x���>��=�<}������N��n(��s��V��D�>2��y-ٲs�f�l�rB��(E���3��BX#�gf�����=���_�7�	�t�G�DG�G������IֺK�)�O���!'��zμί�g�� ��u6�`SP��0�W'^��[���r�,�r��Y�_F��嶒Y��-s��Gi�����4������r�g����[~?�?xg����^B����8����5���W�8��������{�}sD�}UF�|��n�!��3����f���l�>N�V��Vo��{{���n���?d<+&�D���zs�ݝz�
�l%�
[\�o�#{�@�lݨ��TlPR,X�1DU��"� �a�1Acg��+����w�� �A#""���i-�q�mO�'�9i�p�E�k	��y5�۔�=�������c��z���8��y~M[���X��lS�s��ì�m��0��}������w�hf����s�s��o;�ڼ���Kt8���R�F��ΗfgC���Cm�1�}��,�A�rރ-H7n��7��P�̜�k�� �dd@��s|�z�[�p��ח����޾�d��]���I�:4zg_��bgq�`��WEg�x��f|Fɼ0 �f0�z���m�� $	$�in̮X�
����o5�B���te�XY}Q��Gn +]�$𩻪�L];���n����3�������}]���V�9�$=	�x�U�o�O�!�R &�B��li�m��N��6A����+u����}m�I�Z�a��>�yn׽׾GW8�#��i�^�w��ۍ����/WwJ\*�noY��ʌ�{o���S��g�������e>r�b���b�H�EQb1d�@�a(b��3�gx����}y3��c�����}�BN�Ē�H�Z��Y�ך��׳�(���J瞝^���w�[y������_F��|<����4|\�5���w�3�9OI���C�I�py��-F @��O�޽YW�/��*�O�}�%�74��&9�q�K��m�Mó�S��V�}�a�Q�����J�b�3����b#� �p<`:m�$̅�k{~e�4|!���O��Q^9�"�;Z�<�s�Ѭ)Kj���^��<�Y^������g�ἐ���C��D1������c�����١M�d0���TxŘ� �z�ԈY�CW����r��:�[zm'�su��@Y���g�Ɍ��%����y��(�1�H]�z��ɍz�@]y�}��W�;!_w�v��i�EV�-�����U˫Y�v���Z�m7B�#G�[s�iym`���#�[�7�X�^]#�i��o�����,��/�ެ��6�վ��=ӱ�U��DDdb�E��"*��{n;yj�x�ɞ��|�P]�{\m��%���ܹL���>�-N�\���P�W��8��w/k�ծz�+����q��������o�JK���<Xd���}����<��NBT�C�J����y�+�C��sw\��^λE��������7�w�m���D`�#��d9�Lg��=���~0o7���)�����x��rT:���m��;�ۥ�ܧ��0
�&��W�/Oh[�G�Mc��,�$8N56���pRj��w�h�����S�?n�o<>�q��0�D)`S��u����_'�b�Wk�n���M ���`�gbʛn,֫E�,�4~�[](T�Lf������2\��'|���uG�~X{�߿N�tW��,)��sy�<�8���euv���C���,�ݯ���� � (,NUAQH��V3���BΩ
��R�(�dY"�:�c�+3���|\{�����0#�aM�8j��T�e,�;P
�{%q��8���ڈ�ˮ\.�ۄ}�
�h���b����>��)��"�������_�}�M�O<�ns���^^zT��W�{L��8���o�sԝ�������y{Ѓ�q7w�W���<,������v��)oX�� "d�n����}��0�E��[��ݢ�N�C��?O����yF:\�ټ���W�z�ܬ�I}y�ۋ���O��Ev�r�=�Y��҉������[�-�
�_D}!Z���t�O�g�qK�4ɾI*��>���D��^}�����9؁�L�"��-��F#��ヱc�H
��sZ�9J\w�_n�|�f݂"�#Ń��̐����bmv���V3~K??/vI��r�א����r�Ze9�� �@�A�����C
��@���{�]�9؛�Ӛ���F�dPF)�����* �f�u��Ef����g�*x��0.fck�U����������O�ލ'��Ҳۺf�iJLv�r������}Mv��9���M��L�Y�Lz�$���}��8r��nH7+5��\
�S׎_���v!�ϳ���1=��	��ש��diɌ�]Dxͪߧ�&�::���":�}�֯/�󏾏�"��\�{�a�oY�Y�͔7ٞ�I��>�W`l��i��z?Pp����u��q��v� a}���?�ɘ��ދ>�KhJVؿ1�F;�G�\+l��v]ev�zw3ܻ�Rs�*�~���T�Z����~��s����ִ�� ܜ�/�H\C���z�@� i�@�ŷNUj���N)��hb��jjǱ��+@s,�h2��h����N�}��L,�Y �d1��3/������,�m�T�0��+��Q��c��E+�Rb�V�;w�Tʚ$@�.�F��d5��#5��%�We8'�+��nNn��t��Ѣ���}�X����$~��}���X���b����(�@@��d��P����� "+��meU��ŉj��s�Vg�y�`^B��׮�oN����6OW�ﾡM�x�2��B�6��t6'�[�9`-yߤ��U~ɵ<3}��R�j����_c�~�t�m=ד��9���}xD��G�7����L�7;����[�+�l����o��C����<�>�׽_g�k���DD�,�`����]oު��=>�֎�{�������d~M��k�ɟ71���'�Q�^�/�6��7hjBy�������xL�]z���>��#�s*�(,E�	f.��6k8���t�<�W�g�g��ˡ����C��D��z}
o79S���{6-=B���K�l
�����߷�1��FkW�#�`��RJd�,�AV9��S�g�{묍�7��RL�AAd3���`�E,P�����z9�7�w���qj���`��Ή�+�8�)�ۻm#e�]����fΙ~=��_s���1��u^��$�(*K�����Z�o>�ˇu<��{���k=/;�k=�9�!B�)_5�8ץ��?T7Ǧǧ:�����λ��+¼k�GյL��X�s��0�H��8;>F��6���g�0$.�}�d��n�dk���Sr��<��x=��Z�6�Æ.�5����>��� |���q�Վ��9�O3g��'{{���-S뱝��5�e+g�;.����`E��`���g�$���~�˦2c~n\���t���~__�Jz��f'�E���-�m������c�C|�K5!FT
�]����d'�O����7��I�CF�-�Gg���X��u׽�*�BQN���?�T ����Gg����#�^�/���,`�E�I��b�B�� Aګ����[܇�����" N�޾�]c�|�w�7Z�H)!(~�ǪN�˲C���$�ǥҬ����_������ĲU�p���s��W��\����{n!��?��~���b��F��nm����]8c�&�`U�q>��&��2�;p6�j�On�_٬Ѝƍ�_}���}���n��_��=�y�6YDK�)��S�/l*J�»oy�mF�h�_c�c����㷹�~��\dO��a�/�}��Ԍ)��gt+H��|�7���db�X(ȀȒ?j���]2�$���c�ah��ǺpD��D�"˨�d�}u2�_�r���fg$x&Y�*��-E��FmT�ڗQZ���*>�"s}��R�z�4b�-��<��t �^(b(�RzKGb�V淉�z�Gn����N𾔼�aGMg}�w���׮��k�<�g��b���a�|{<�f9���Ѹ1DA�A@���P��J
2�[fr�{:�8T��(�׫��7��8�$�H۽b�菢�G�A��q8=�s{׎g�6̡0�6�(n��y��	56�ɳ�=*��"[����.�0�%�PH�F�<���r�klm�}R��W��y����+��ү~�9hJ8�]Kx��ﮕ����[��M�n����պU�[��Vc��y-nN���2ZU���ly�^��ؤq�[X�l��?\����3�7 y���W۽ei~®�O��omݿ!˪>�+�ف.  |�L�y���i���ҏO(ۑ\h���G�;U������J�BC��b�g�Vh��٬�|��b�������;����\u��؇+舌 <���}��^��xm�4��Byo�2�[��y��J���| U�W*y}�9�f����w�]ӏ`��t6��45�^����dECy�
��9x��7�u�n���e�I+���T8躌��k��8��Q���a�6'�7�����[]��[IM��mWz�t9Z�y�>��:�6�D{���{*��6~��SټiCe��VN\b`@�������*�J�d�s{���`Z��0���q�Ȟ�Q�o�1�Ҵ��>g#X �1r�u�k1ӣW\xV�AC�ZOhGZ�@0D�`q��ɴ�ɺ+.���W3`�a�Sg�f�GF��t(_��n�T���P3M���J����u�f�>���2��'mA{(R�:%����D'n�c/Z�k���ڷM~Lҡ�#8��/)0��w��>�WV�i`�.(�D[������a��jS �&�y�EV�$z���:����z,PY9���Zp'��Hzu��x�gw!z�aux��	2]5��X���x���Ib�J� 7��p�q��".�E/���4��L6�n�)ª���)��5͛�]���EF�7*��_�U�r5m��vε�g���Z���Y�j��˷WL(lR�-�\���}u��8"(�b�?1C�ɪ-@�lU0"��H(%6���H)X$�&
h0I�J0_�ׄ���,UU���gЈq�`# �N��e�r���xmN
�I33E���^JL]⍈���';�e���S�4�5�3�Q�)ɯA��\�1:B��nUc"��C�	ٯ�����dV��n]N�E��"\�PgkM�^�qL�b���NN��uKq ��_`�pw��vk�y ��Μ��-q�(V�3(Ӧw�5EZ��%�h ( �"���m������%&B,"�6�)ӣE�4�TXd��m�&�h�(�J�6�*�i��F�h���wI�P�uE�xBT�x/��ʑ�,dP#�칏@f��:��p����y2�咔�K��3/h���uӻv�&�����^9��>瓯)N�n>��Ջf'�|��}:�7��k�ZҘ���Z�l�%���.�ˎ�����и(��ڷ�N㢞�ie�c'&uf�X�k�Jѳ�&XN�!�d^���H�DѩOE�rvEܸr"���|\kq�Z�DL.��t���J02��wA���!l<��ݹf���a�MQղ�rʏ3앓\��1�Ci5�Z��u����Uݶ��D�6�D�E�|*.�ƻ���^�������i�-���=���m�d���Z��q��%5nU�ʕ�b%<K�r�y5��Y�۳m���[��Q�9��QӮwY{9��0o��8�B���CrZ��pք�[N�$��?]�5������/fY4����;��E�bP���p�ZۊցW7��_qA��F�&u����.v����x|�a�ns�Mrmc�ؓ�b�I��g�R��U����O40��Z9k�\��+1���Uۖ�4�-�6[QIy���W�Ҿr���3��:�����2mGD�� ��Xk+�A�=�bAV��3�q����ڭ狁/��J�ٿ��=�#� ���j.+֝,*�-T�أO\��#x�p��SN�L��b�jD���G3>wh��mitr�$�+0�G�p񺾽rV*��nT�W��t3cpe�%N�K���gWn�/�Gp!�Xo,���e[�T T�
�,��h10���̒��Q�JE�L�����ي:�y-);�����N���5[\:��c�n�M@<��*��N�7*�7�F,]'ڹ�����y����.�n,J�����X�,:ha��lR�#�=����5h��lr�����D�b��>���8��k���k��[ȧ��}>�f[.Ʈ�/������J�'�[��S��|'��ѹչ�/v9׫�hã/EC�Z�j�6
 @ |��PQX(���|��׽�?_�����>�_�?��P��	>B�� �bѲ�p�(w;f/F��9���qu��dQ��L�y����}��ڷ�Re���u��3Y2��LGяy�>4�N�鸝�랖3V7���\��ow��M����b���O���y�Q��w�jZ
 �PV""��H��>�T�i�^�;�0��i8��#~T�"�'7� M����7ڽ���X�gy���� ����}\zE]�{г�Z&uc�zZ���~��.���ɡ7�bn?M�����5Y:��FD�䷽޾���w��v�����JrJQ� 8��}�~nۙΡ>z�Da-$Q��� ���Yy,j~>�q_MSٕy�WJ�����w-�^�t7�;c	��9~{�j��MM���f�DK� ��~�x�碬�rfY��7�]e�K��v��ȇY�9C��gU�ܯ'��V��u���]�9�������na�� �D��@:�PE���{���7��f#k<���e͗��s�?I��u��B�k��r��f�v��h�ϛ�ӹ���u�]�S����b�������R�m����[חq7�ܝ�ki��|��#\bw�%{-6��{��d���ˀ)�e`F�P����
��w&`
����c�7��#cVUI>�	�֟p���X**�FK�n�̨�E���� �ʷ/Os������g���~C�и���ú1E��x����ܻ�t��u&�#|�R��]{)�:�qX�R1uq�ҹ����u��C]����q�ע���~o���Y��0��f"�|�)�������5�h�5 �EU��Z [{�6��:"���VY�Y1�VA�Ҝ���me]�����TS�8�ZSu)33�l�x�^����a�CV�����	ֻ��[
߶.��z���؝�ER��sY��u��~�F
�UC��w�o^1{����V�Y{w��~��f)��Ոu����щ]8m:;�x������Wԗ��p�г�����Rr��|�e�D��p���[<sN@��ud�"���e��|-Y��<c"�W�{#_!wVfx����<��L.���yp|9����n���g�_u]X(��Q�Ud@DNg�$�H�ŀ�_/-i�?{�������DGd!f�`i�Xu6���r�����5�]�7{l��� d���t6=��~�<���%X����v\ǖᚮ����9�dG��t�b�M��.I���JK�����5>�;����d���2�Ճ�ʮ=�"#������MS��y��b�U�EU%��O.���X�ܼ6Ї*v,Bk;��f�-��K,$S-����1�L��+��#1���^��+������6�eEJ�<��)V�c���=�

 �+8gX���\g���ڍW�X�A�Ԍ����3Y��w՗����w�u9���[29 {�؀S��(j����[	�9=}�/W��l�Q���gw�}�#���L�T5߹Fh�Fz�B��6���
{�ێ����-�����;���W�p�XK�!��8����D�.�k�]¾����_�دg��������uY�� A�ޒ��>߫:��|��w�>�pT��X*�+�B��:����hQ%���x���:�[YLg]�t�x_%��Pz{��[�$m5Sۛ=������Z���˾��������>�Lb�Q��]�
�c�}Or�y����˪��>��]�K�JB����7�w[۴�yP�ź� � @DV#��Tz�k-��E��(�PQPb�*�(�t��D�~S&f�Ƀ�S윝kUl\������Q��X*őQ���ZI6ѤYAM�ПJ��n]�*��2��wS)]͠9�>���9�֩�;7o�)w˪n�e�'z�k �O�˴;��`m��n�+=�ZU�` ,�C�RXs�T6���)�RKWD6Am"M�OnhガV�}��9���8+׊> �� 1�'ۯk�9^�-����}�!G��{*n4}8N4�ľ�o���X�q̊msk1R�߽[�ݝY�]Wg\��kY\���kb"Q۸���㪆_D���f�w��]�2��ʅ�\/-hw=��^;�V�T���K��y�`3����-��]0ϸ9�	�J����Sy�DB���H21��b��UD�(,b�0PX/~*! �Zۉ~���;�������R��������ͷm�+y�uf�����R�|$�,��*Ƿ����s�]����Cur�&�^
w���o��|]x��X"�b�}�9HW���L�$�>^�Sr�I���u2����fL��{|i�-�{�����CRwt���	�?{wި�Lo���{|�.>���}�
|��}�����1G����`̤'�>I���&L�Z���Tyz�T
>0LY�!�f�3S5|���m��0��I�f[(��&"�-�LckY7a�^PgfSQ�z�2�v��*Ek,yv�R��w����U���=�9 5w��gj��Žr�T^�7#��s�Sj�۠��v�;���DDXB��y�>��{�{-Rs��P��z;�5�q{VOw֥h�Q�9�T�/m�fU��ֱ��Y�e��ԇ��s��������
���(�"�U�$E+�	%���IU�ǝg~�:��l�D�`#��"�Z���:����j��qM�UL�̜���/5#y_G&=��2oO����{B�k�l����zC�/���Œ��[�.:]�w��5��z�3��2C��}�5|}uOk*u�ѮC[[*� 1�bX�/�u�<���NNB�g"�}S/��+ٜk i�r�:�6���<p����	$ �AI�;�7�M��[o�Op\<���[r�Q�3�w���F�k^� x�Zy��+�˳���>Ga�D� ��/Sͣ7c[/D��iVr۩M�]J���r��
(]����w8����v�ƺ�ެ������?�]��_1ur�s���Rcm9�����Ic��l���"�WYz'2���8^-P��:3�Q/���HOs���)�/ tȘ���z�}~~���k��S�BtW�s�ڼg3���=�o������22G����W~}z��z����� �TUEޫ=�I-�(���7X���~�a�Pqr(|��X�5Q��V鍶yƴک�:��Vw�7`<�Vu�|:����-N��7*�';н]���kU�B�^���[�Dp���+��y��2����wxzn�.eiܾ�}�"��N5K�G����
��{+��/p����ʽ������vw�������h���" �M��R�.���܌W���)��޺��o��5��9��.���1�1���]�� ��i�K96	��D`�_Rf�vs{:N(0D������t��C��ˢ��Lż9/%pMЮ�	�u�&]ٰ�*�gd푻��.}o4o�@w�]���QU���cV.��^������ٍ~�)2�C��E)��#5	���L�/
nϊ���%��� \z	����=�D����I<ޯ���k��������$Q`�EY��n �F"("� D~?�Gҽ��Q�����Qѽ�+!(͂ڲ}����>�U�J~�	���,�����S�	�k�{j}�u�w�=��мqn^FN���k�|Y[q���D\/ۊm��̅OR��>�2���ܿ)�����Mo�Tn{Mk�����.dO�y��w��:5�y�z�����^���6�����d �'}�}�}���Ohչ_]�>���5\���W/�}+t��=�U{p��g#� =�tޫ6�^���I�x������-�����j�f���"�d����O�y���e��_}���B�-��b�&��R��f*�wD6���6\#�S�Q���-��!F��0q��lB��K˥��C.�� �(eh��{��Ǧ�m�{$��2y���FN�Ƌ8��E�NKa ����Q�IMѣO�nL����ȓ�˼���s�����o<r'���ߵӱyo���m�Wod�/�u��wo�m��wF��cܧ��'�7�Fϣ�AE"�1U`�F+�
H**���u��+^�y��U��=� E�#�&1	����1����jut��r�0��n�}|f���\�ʣb�u1��ۆ�a�(>o6P(���Mf���}xc�3���`����>`Fs��&�b���Uz�Ta�/;g�,�1zew��\����O�l�\�+U�/�mM�Rb��S�OQ�Hy���^�c;ϱ���&���z��P�v>�?j�uz�wn��nQ@�߶I����r��Fqj{�IQ���E��k�=Bk��0�S��)Z�)/P�D󇰱l���o]��ͮ����{ҒI�|dMDiPw|�Rcxv����{sn@�� � "3�n_�����z&�O=^�q`�Z�b\iȈ�$��wg8�㦹=�������k���;�����i�H\��ݚdL����I����o�R5bl;�Ǝ�;4`�q��\��^�Ν�W�~8��꼻�ʐ��}����ᝏ�	��+�N1�W��<��s��E"��1PEQ��H�yD- "H�`��7�z��L֝��i��N�=��;�W���ͥ�6���p^�ay��;ܻ�j�m�y�������[Ҍ�E))\�DB���Y��S>�3����/�q��}G%�֥`�����H���kݴˀ��t�m��7�^�Z��}�խɟ}�319Yx����'ZܣH~��6�6���}��C���G|�g/g�_<	�o��Z��{��}�ae�=�<�{ºL�����_c����^�^כ޷V_w�>;2�p�i�ҏ� ���[�r��}/3�{s��jϮT��<�^N�y���bש��EmGڼ�+V������`4y�W��_�ru�R\�w���yN(�+������2�鵙WX7�u���;�L�5���w~�p	�W�e��̎�Qu:\�0V�G|٘;3pOt��_}��tj&�06�@vb�,�*�{?_m9�XxU�[L$��e�WTQ� 66-�4\1��I=²��Z-�U�>���3���<p
�F^R�\�>]��S$��4p�/�#u��ܔ&���U�eAZ��bK�-W�+�+���>�*�f���O�Պ�����k� _I���O�_^��I �شDI����R](�L^ތz���U�b�`�,�&աN�,{u��A�i�*��>��Q[x�r��ӧ�XEhB��n	�%�C�B��:r��X7 r֎ +�(뫛�J5ơK ]4�i��(Mt��۔�ۺ��;��f&�H�������}Ni[�y��U�Ӣ(�N�@��8�`���M�����	�$0T�MH4%0I�$6gKi���"�(9��Dka� ��2(BB�����{��Yyi+xJ��S&�X�A:����,������ܢh���S@3Y�;�m]J˩��9G[�Y�I��ʑ�Li&����*�GLУLf7b9��|�� H��1�s
	#�\�O%��y�k]�+�#k�wUk��U>����77��M;
�U�s:� Tn@+Uh�׭�w�z��X� �Ɯ���Ș{e��X3���%%	�t�b}R�ܒ�3F����"�`V�Zw��_h71*7�B;�����v
V9!�\A��1�p^-N+cV�7�Ѿ���3y.��j�]i��31�]uݙ8���P�٥�X��<��@��4�#�ڻ�b"���j���tQ���YW�X�ĵ[��9�Յ#O�)54��/��̓t�j7�|,�����c/�w�s��w���chj�D.�]i�z*�Řݣ���E���s�C��t������ifH�Kѱ��T���u/��wQ��j`
c\��4��VU��	m ��bWFv�2�C�MË��-��3^�v�����O^l��w\�)k��̕Ϡ��f�I�<��F��l��ֹ�B�{��e
�yC�gq�r/��{1��{�3]l��Egwʳ�sC�JȲ:͙PiM���4��*u�����CN�Ny^�k�!�>����G*�{s��|�=7Y��<G�smk7C�G��λ�:eJ�[tUq�*�5���Lu�T�H���1��꙱�'��-���)�+�bb݌�ќ�.���N�ޜ�N6�WmI�]vuj�4h�&�ss}'j=�����_�1Eo*�-��k~���錚�'�ܒ|���$R_ݽ�QXDV&�R�A��>1   �>��mn�׆��A{��Gb�X��{��}�W5�~�S]�e���v�ͦI��=�w�ov)\U���0�C��u�Ϫ��_����ݦ<�c�R�}m����
}P�'�~�����p���蠠=w��q�C|ʆF�ym�v�����1g�E
Y�~데�~���}�z�Ǜƴ(���e��G�s���_i��$�Ѫ�������<y
��Z�'���.2N��Q��vQ����K�5�[�!<K�)Ro4pާ{�O��ь	��F)YN[�u�����F��~�>?[O�b�V}L8���ޱ|s;Ӗ�G���d��o��}]�;�v������ɡ�F �REE)�]�u������Φ�'D�J*q�\�IL���X{�o���OB��cmJ<�V��B��_d���O���t)�9�a��� �C@�MY^�Z�������;�� X� b2)Y`�("A��ʎ�/�c=Y9*�):��F[ɾ�6�>�W���k_�3QY� *ھr��^?,1J�E��J*�!A�=D���9W0�ŷ�No�ZN����"k�I��j�-Ljn3֒��g�e�{��[�U����[#�J=����Z�v}�ٵO71voz�w�����k\�aLK��FO���y�EA7�d���k�_��J�t�s)xg��f}]�ǷOʇ�l�mb���8{�{��z�9:gPp���7�������R�Wx��u %��~�")�j�%�\ϓ���/��Ǔ��&�)�������-K���6�rB���@�{�ݐɞ�/ivg�DJ��	��*>�쯾��Ըw{x�i4��DH�����DF1b�Qn�����\�uX��
�$�ʊ�����BIk)��E
*l$�2x�xfG�p�֚w�gu��C`0�����M�w�ų�����U�)��a1��c=�!4Ļ$^nȮf'.�pB��1��g�.�h�6�S�z��"�HR�L��}7�n����Ӛ�9k��������o���V���p�q�[�1	>��f����ܞ�]�������.k��4+�n�����Xc��%��-���3�~u�=�a�R犅$�������w=6O�k�OJ��]��]޷�U����{������CGV�ͥ���y4s޳X�z|�A"	TjUE�3��p���c����R��i�}�Q��jP;�c��B����y�ң��{��o�SIc��wk��O���ߗ^vWuiZƧ�U7ܻ�������󏾓[���2�HC'׊����r�2OM��͛�X R�N���<��Tevؖh���,u��K��˘�^��,m��1;�[��Y�`Q�����{��s�2F	"őQ��"��D@T� �!"�#cHSR+e��bKs�Òp�,r:�+�(�xK�c��~h�/��ù� @s��\�wu�_�oPUGT�%/�<2S�-�1,/]�{S���<��*]�92�MS�����Puct����L���"����&[ÿ}WZ�ù�%���r�/{�Fi�M,7^֢N뱎�Gb�1�4�ae��>��A��sHGA3>�d�a���/n���T�}�.�3�]�%��
��e�'�1nid���c��o�ϲ�6�gU����(��5���AWϦ@�`�0 ڬ>d�'�y.}��5J�{���,\C-�U��,������')���΀rS?S@N�L�lWy�]��"��uת����}�T�OZ�c��W����D@jݗJH�gNǬǏ�޻�h��j�	��z�+��d,Z;�Z���j���0�B��2���g�0����|��s}�V8�E�cr_��Y�ge�ݬ��.κ[����Q����H�"0`��� ���%+0_w��k������af���6 EZ�_Dk~Y��b�Jrl,/N3Nt�����KV��)���,ʼ����Q:pP�4�np!ֳT��o�g���w����������Y�����V�PT٣un�]X��"�N���&򡷸��XB}aX���Į�Z��怖tf�a�ok��7њg�t��.�v�8���b\�2'��x�5oW�]Z4YeJԼw�"�I�7�P�A����p��2N��gNV��^�V�Q�u�e��#O�Cԗ7�\��Z�� . FM}01 .�C�/_�b�s�+��EO ��W�I�'��y��
鱲ܙ�K���N���tL�+&�/F�_S8�³&nX�)�s(��'x��1���bNc���&���^S�g�1��̆^b������o{����uf�y7���,uk���P�b�5�_!�P����h���C^��=y��A��~��"~nͭ{K~�L2�T�G��`r� �Q�S�\Y�*�A�H*�Q�1�$��@f�AQ���2w׭��9U�Uk#kG����NZ�!�=s��2s}o�aD�T n.��]����%1cd�4!�_U�(o�>��<��SFء�x����-
d{�~3�ժ5�INn� #������W�wX�:5�ț�.g7?u���@�M�J7nIų �]�u^�Vh^E��K�W+�ZDµ��L����ò@�l��%��dc�KGdǓ��������a=r|��bc6A�jY��,�(r�Ls�ؘ�p}�<r+��%Hd~�_�2�!�܌M��}��o��5N,P`�
20��]Wg��AN==�{��$ѝ��e����M���[tqG`~;f:��N�U`ML1��y�n-xŝ��&�c,��n�yWq]{�J�v~�ڨKfE�-�e����Dz3)QZ��B(�n>���sV�O*�rbl�,D�?y)��s;���N��4,���/�����o�R�wC���?��!��򾫣��g�K2�f�x՚�.��n܆�"ň#D�"���(�b"����A�1P���w���b\1��`mb��(�#��Z1aIAn߽�~YSA�#�}>yN��=�݅;�k��ZYS��lǡL�}���o9�	�N[/ }Y�����LkK�y&nN�����H�1��'�>p���]SEz��m�f�@2L�R��L@F=:���x� 	1&�T��%�KiR�A�?���;��/j�iL�R^erP^�jĝ7]'��(�l�J�M@*!��7	f3�f�7�Z��I��W�8 �7������`1CLU�jN,I��.PP��5(H1��_n�L+�t{�>d���a=/_L�5�N����5�a�%���7y�_~�����2G��?	�{dYq׳x#���T���	 a�^R$�ﶅ��Oe��s�y+�	��R��&�J@Ɖ�=1ya��^��h��3���⻔��=��s�:|bT�q��,�&�z�����6_���͋��Ⱦ��O��
��ɏ #Αɉ�4+,�
ܔ��#�G�m�U�L��������5�5�Em���m��}!c��c��1�x�)#Z��P�+`�bE"� ��D�(�|�Ea�* ��{8�>���
����_ŷ Z���~�9;"3�_�ۺ�/rbt��B�u�v���9kD�b��<YXU1��EL�$����-g�^��Tި�9���¡D��X�Ki_{���1>����xO�+�r��C7sڐު�)���vI�ӝ{�mD��Q�=&*���c�U�Gld�l�H�G�D|���sg3���k��p,d�0���i�U�l��8˃��I���*M�POV�V�[���\Ht�Dm�Y�;��/))�w/�I��/�'{��jY&fFi��UG-���[3%�/K�?i�u�I2��5{�=����߶I�$����{���=���lbΩ��G���\�#�U�CVR�]7E>1;2�E�&B�հ�]?nZ������ޙ�nO����ki����ž�[s5��ڱW�aD⺙��́�{�J�.dxx��Ѵ���Ū�G���<Lj7���H�y��h��W��`윷��ɥsZ3���3���.�d
?�*�*�����F���"��}��m�g��9٠�cH�F
/ڰ��0U$�G-��f<�Oh�7���;�h��
sD>�IH�C�����>�l�L�i�,�!�c:�����j��5��u�i��4��Rڋ��#�%�;UK�*�c��_����jƄp�vx��Nˑdڔ nO �uܻ�jz��kB�'
�<�,��0��=�'گs÷]F'�xR���!#��!Hg]�zG��-�<�u��ͭ�I����V��<����䨥�r}��[�I���V��U�n�YN�棆qġ�3�V�fC����P�#��ߜ}Ip��"�I=[ǜ�{��*ƩSPp��鿻6먭�.�z�nB3�hͭ����WI̞NF����`�gC�~��]�Oj��z�Pˬ�	߭����:��NҊ�����:�~"�I��-g��y�ݞ��Ut�G����
�H���z�=��y�!ԇ.��q��˪�y�K��vB�iw��l�fι�u��-U	*�NV�oOY��ɯ����QTE$UEX �EX�����+@U�T�"*2EQFcP$�$ %V�f�s�u}캇�L��o>& <�}��O��d|�J�yGJe�#�*��?tG� ��WZ=fY�3�_]�u�(��a=�����<�]��C�}`���̩��FK����#ݔ����b�V����}=�v��q�C%�=]����c��w�B%7N�2���wJ�̊��8(nn/t��_{�d�ς؉3�;� ��DD>����A��Ð/�SΙq�Q~ib**2 ���E�1#F}U�a�~�2Zx:���k��h�B�
 p5C��T(
�����{q�s%0���2&zb�K2~�4�]k�-]t+1X�kô:=�yjX�vTPcz�v��!f1��I�1����pfύ����G�$����S���wH���H�r��{��3�n�Y�*1�gJ�hh��h :ޝmb©�4�3��(�x��n@�[Rvc֪�l��B��='ȳp�����@6�>ٌ�:yQ�&�4������#��"�߹��X�T�1�X��"V(���H,H��b�A�Dg~��;���f�O<�ϫ[�{�mD�Dr�g]�?hR��I�������M�¼�:��x{�zO���)�S�CA�Z��!�?��!ߍ�GbL!SOΫ��I��!a���|g���O�xǬ�tt��#�O�*����#,�}7��vTڍ�����;GO�B�QV9�1��Ώ?wE`U�{��9��9�Y�������7�n�}� Y�(V�Z2���r���<a���'�n��};[ |�$ A,"����L1�u�����w�`�E�$���ks�^�<�/-ԫ�ˤ���I4
��S���bP�X#�DC� �J�i�FS�zP]FRv^��n�b����S��q*�=6̩��ntxZU�U���T��
5��}�ɘ,1(��Ku@VF��"��4sz���W'G����ٚoV�(T@*�4��<���NK�P:fWkn���B�]gɳ���>�d������]
�YQ���,ֶ6�_`��EtR���"(iӬA^Y�����j��h��Ƿ!vI�ȥĺ������tV@sv�_��%1Xc�#��5S:8ܡb���#��}F��C��������cmmI}[|rE�\�����~��84��9XuvPa$��I�~J�:�8��`� �!�!3.�4�s���/#�W�����ZL	�����}��x�!O@*�������2ee�|�k�/'M�C��A�?R��Y�J��Si:m��0)��(�2~�1
J�	.[S��[���b'eV�@m�]���
����_6[U)1T)���qf�5�P{�OxL�ݎ�.����Q��#�Ҙx���2+4�c��!�@�Q!�R�X��xj������A,G�oO�m����f��`L�D2*�TX2&,�˺�VR��z�*l)�(��!!� � "-�k�t]�����E %�o� �uЂ���E�+"���6�ʨ�-��Q� RP��(:"�lKm�?�'m��m��I��%�L:$���*d�`2Q&��A0� Ц�`*O<#�B�KQ�-�no�gEt����j��bWq�H6�jlU�����- >��H��6Y���d���w#<����U��P�|�}u�tB�dL)}yf�.o
A��.qe��v�)ˑ����v��d��l�|���[u�䂃�]��A��6�U����LX�l�(���.h5*�b��$^�C�VMsl��ongr���wݩ���^qK���[q�ٱj��d%qo[3��X޷-��r���MǺt�֊��W�m�:Z�E;xW;Q�vN�*V�X˥���|3rI���J���G��}�|p,9��>�yB�m�{O�h���&Y[���Dқ����*��6������0e���ri�/W��f.�[���G� d�����Ğ�Oa][4[����j����o�KJ_nb�t7ٱ��q�����yS	�\&
�V�\�ܮ����U�(��s��hNw�)�eTsf�i��P���z��իjxk:����.�a��:�×4��W+(c���6e8�\]e��`d�������p��O���Ǖ6>)�?o��y�{K��-]b����n�F�+\h(p�7h��hD{��	�*f�t�M!k���݅�A����.��]y;�H�_ה���n?'DD�c����+n��t���J�@^Ұ*��4B�]V	��e()Z7�У!����(�v�61�gd����%��`�'q����=A���Ņ�O�p�4����d X����A*�b���H�*�#�crS�q�6�M�}ٵ���
YJ�ۉ��2Q��̺Vj��3+��z.�����2tW"���7��l:��gT~U���w���e�D���9(
a�$g���$X�������Ipl��7��x�^7��Ƣ���;ӗq�0�!S�Z���~ź��m}�UT;&zrci�R�"�f�ð�����K%���`�t�P�|��venz�p�G2d�ޗL1��fw\kʖ�ژ<K��DȐ�oݭ���@`ਜ਼C�r��i�E���bdW!3 �FEA$��3��:���rvр���DD��۱UH����������� !wu@:o6���S54�����<W�pͺ����ㇿ;�7���Y��2$8��#[TC��Iq���>ɐ�z����{y�iO苫�!��J@s���!�#8�3�J��j`*k����k�Q%���{�c�_L���!�㈦~@�C�1ʶ��GtT�Y�i�[�`REԱ�x�6$���^ԋ�F(��~�As�N�J�Oq��;ɺ� �b���S�4����A"F��#��i��vS���bl��Ĉ��}H���D0#�"�DGB���ͷ~��`E�di�D@k>�z|z�i��6a��v��>��y��%�6�Z۳(9N��+�ܹ{nBc����u]Ν�M{�X��}߮x���u<��K?D@ʜ����Gf�Zg�!Ci��?.����7���	���ecS�u(�q�l�R��^�!'o/��<¢Җ'6g�~Zz�l==��55�/�^o%�BMb�^&�	 "	$�U)^�X���=�u��{[��uPDHUU������2d+�=ӂ�{ӡb�"�ѩ�r�����t�~��D���~��r�qw����{s�\C�c=�1��xN5�}��)�g/xy_�K�h�
-b�a��W���i�7_8��Ɏh�u)�d}p|���l~>Nݰ���jM2L$W�f������ɕ��2UP�
X��6�j�]��ێD���Y`z�CLw����3��7U���v��	=�I���Gw��Y�v���U�;5�9�2d���X���.�	��@� t闳1��O�?-~�2�_^��t�6}�{�=�q1 l"�hn�kH�g��>�+���B ,�ƷX,�̙��1�ek���H¾���}؂=Dʽ�k�l�G�dMw(Z�x�Ǹ�:V�_E��%�6~�#��%��S&�НYl�����Oۀe&�̂sE$��������c�uD�澁o��-�h׿a��θ����u-�8<��r�~��R*�(�!�HR`��IDM�����!_��c<�!���70 �@��� �Y+���;�wW|`��T�,�p~*� ��-��r�Uۆ
;H�)+K��U����
��+���7�\I�����!�MF{�҄��]󌛀}~��×uN	�>�4���ϏP��ړ���tm�^�ͿgW�+�G�h}kN�g;|��P���ƍ+icoy��=���O�!嶛8)�$/&ckUTq�~�ٱ��B!:��/;#���{���n�I20PA�`�}}��r���m{���^���R[��2�AK��}�l0K�)��~v��~֜�����8����Ozp�ˮ�当�k����T(La���=��ƈ[?9����z2GȀH�O�wP^Ӝ���	��!�R٣'/7�����\�w�Bf�u$ؗI�d5�.��
��y]�Qީ(�ē�.�}]���7�Cٕf�{�˿Ƅ�^{Qҧ��/b�z.;���yR�e�R/zj��}�g���֣�㫒�f��#�y.����r���BB����^�[0*E,TH�"*F(1N�6DPA~��3~~���OX#���x��w�@Yޙ���]1�cˢY��9���q�w�t\�S�d��p�HrI��m�� ����A͠fu���{���7����5.M.t{�`�	��!��n�es�k�v��^cB��t�� G��4G�EB���=�}�T�36i�t�������8B ��ʺ��}���.�H�#�:��9�$��x��Ke'��e�p�^�+�u�&xP�a���Չ�S[ܸL�'g1��=[柫w����=�@N��v��9NY��5���`�a(��'y���+��!���dLW��jCɄ���K�Y��z�>�O!�@� o?}Z_�[�+��""L@� ���)L�P/[���-"/��b� �9���(P���0\#�:��-G�rm�����տ�7I��@��������A�ݯ�h�wAXT�1��om�Xm�uy.'�7�*�H���p�˫�ݻg�	�|Je�����n�|:U
k�{��L�ݭ�QP�b-���2�H��� �X�}��*Tg������w{��I$ޭ��d������<Z�X�A��/y�{9x6F���iO�y,��v�$v�9��zuxO<���Q�Jn�@>���:��\��eo�^R�x)A��\��9�K�lǱ��<9��h�czft\��R��W��C}�9��F�����<,b>L{���T-.�ʼ�9Iq��f<�׾���eJ3gUP�ď%ƽ���"���^`
�Dc��^~}�\D�co}�s�%M��a�L���nX}��$�&4�����Wǔ��������g�q��7����5/j��g���K���^�V��fdď+bmjۚ1������1���H������'����G���	��DG��\��Ӧ�vQ���ײ�u4>a92��ع\������J�"��ȤYV�1�P�`�b!�b³uek���﷭oջ�"�d�4�T4�L&�\%Eb(�F
�c �s�+��W� f���x���7�	f�T����
��f���5P`v�/�*�;IN��M��[}���K��R��ٽ��{UIY$�! o���Fi�����=�#@��U%�K�s��;�y�+���;���9�V���a��ڙ���0b�n&��b]�����'����^_g���3����Q��@��&)k ����^�'9���������l�>f.�9�NzGi��Hk�� ���w=��g���Xkap�������]Oȶ�lyWw��<��.ʔ�C�xS��M3��Y؈�5σ��݈v��i��ߟ�0��='�� ��l���j��OZN������e"�����&��o8�x��h�:�?Gn:��Q��ٗ���%[�J���}[5f��G8�X˛'Ѷi�1l�+s|�������<�^� 8���X&~���Ou�U�!���Xcx�Hn{�W+�*�.�kDż+K%��T��;�FuE7�����k:{t|��,���	��#* (�j�Uc�+������ⱂ������T�JY��$��`��5Amm)SiB�
��()���g9�����	Y�����܏o�bE�ksmI8nTM��"oM���Z͟K��I&	�������wU�*�@�=&%��<Ҋ��r����.��V�H�4g���X��V���}�1�힯�Us${
�Bw�uݪ��J����g��X���H`�����Y�;<=���<R����;��0��}�f{��'�"�`�;G�j&WQ�dB�IRb�o���7H����Ԗ׆��r��hjnO�M���6ӜZ[f �����DEl�k>�<Ifɓ�LQ���ޝ��rL��O����#���T`5�~��ž� 9�LR�Ѹ���T��I�!r�:bn1��%3�9�Ě�"�������Mk=�ô��J����j���y3V!q>ɵ"|)eW�S�\1��;�B;�FD�� {�bƌPdA�l���
�U�=~̢ڡT )�� �U��yv�2�bAw�>Ͻ�V5�w˫;�`�$�F �P�&��|e��^���r���kK0�#���Q��^5E}]�X���0'a�(�$�8ɞ#�w�r�E+T��qݯۈ�	]nT�#>Y��� uӭ�@�0d&
�A��r�T���9�Z=�+���
{r�XDu}[�������f
P͗I�M���Kؽ���3��d&���-�6��O� (_�r��d����,[�B�0VjM=Z�K���R�T;x�:J��0�I��UB�U�k��/�{���f��2�mU��!n߼ن-��Z�F���Ny5Q8}��}���>��n<�kb�D�0z�RN�Jp �{����J*�1�
��lwkx���y��U��e������[��Џ;)"�o�{	G�Жn�,�>���<%��tv���5���x��1#��}(���EǤR��篮?�/���2�(��׻S�Q����Ixl��,.��xNq
���,�Df6�`��!����gÙ�"1�'�	q`�0L�_��Qg�V��H����R
E"�|��{ٸ�ݺ�zb���	��(PhtΧM�#��F~���+���1 F}:Nv��+�, �a�M�@�[��#�L^1�c�)S�J��ʻ+a�{s�ġ���v��NDWNã(:#6i��J�NO�b�h�W��u�`_�g��&ɗ��Lޒ��1���Z'^�1P�}��eG`�����&�k��e,�Шk�B�@��{�b�HgN�*�Y!MP���r8�"�Ar����?5$�b�,��F|��Z;|�����^�}g@Fr����l�V�����o�����Tn�Z�~�N�=|���OQ�#%͈��Q���4��\��l*q�=u�e��|��[x�ڳp�W�1��������hk� q\�PRP1[W�˭�2x]�16R��V�,^_w�U���.oz���u�'��MC�M�>�(VFt����*C��I���d�U�yJ�G��p�-�ř}��\��V�w����X�K�O��"3T���Z`���@t���Z�{ί����n�Vhj0���x�	y`��{8�k���5�MC8QH�1+$ �E��Fd�δ��Q�9	���)��i�e���9h�Y����������ԯ�w茠�P�����ީ�H
�Ef}��S!�L�Myb�n�^6!IJ
��@�#� EMs��O_��n�m͔j��,���>��&������<:���n�����dyX�w�Q�WS��F��[-�5�����\x�5��*�N�=��z�4���<Y��G���~5e���ƈ5j�7�.s��ٸ�����A��ᗀ��
�}�f��eب�a�w7��6����׻����Ɩ�G����:	1$}xZ�=ݛJ��h������r�2�?A߻'/Z�<����"=�e��F�3!�5�w^�<웿ݥ7�^�7��|�,Z,H���N+"𕇦NVqA%O#?���%����u��}��ǆ="�Ԍ��V׉!#^�ː�||<N:�O�.���n�Q�`���RZ6�S�>z��8�멌x,M	0��
��1�b�YDUF1��l �W�5�{��W�:��y�>�BD�'~����Xޫ|k���b��5߶�ut���(�@{^y�t���q��!-��)Z^��{�D�d�7�=�.�=����{K2���ޞQr��87��|YP��R�R ����߸a�i����>��0%�/�)��0`?��,nq�������>�[��Nc�d��ᬝ�U��~��)�9l10�<ʳ��҆X���*�r!�'�G��L$M�d�)fT�s[�yu�[%�[@2
���Ȍά:qQ/��/x16Jc��O���pQ��,a�$*8+iZ��e�;�λD����'��u��6���%�I�McT2���耾�n���JkV�Ql��躕u9l�K	g+Y2�RA�`����I��G�����+1C�2�l�"Tz����hwS
�`�K�k�Ǔ��HȄ�yn��Pҹ�42�����r�1�j�z�Y]֝֕�����w@m,N�X��>��rP�����u���1�s�����B�ߦH�5�%�킭uI9�e?��O��O+�ݹ�v���i���8F2�IS��6@��Ypk�;{��]�7�-��Rt9��f�Y.b�cy����S�7���P
#����҂p�Q.����"SFH�RY�dN�:��$���Yvd�"0 ��1�Ɋm�;ZLꧣ��˻D�����J�x9�L�[�Mo��:wG�Z>��&vw�CD.��j��'g��!��`�S'�L���f����N��A�}�eY�TACM1�f�)]��m�����������p
{a�I�*)���]b�Ō�F��'k�z�F��:I�Ğ�{)q~��w+k�h1R�˭�.��5'f�[�&�Wb�
��&�V��4�:��0��@��i�ȑ�Ӂ����x���ڕ7D�cuk�����+S�s����=��wJ��pf�.7��}6�),���K�f��z�B�F������lY���ɺ�&��h5#���N��(ma�w2O�J}�f�F����'V�s�)�N�U�WQ,�e�k1�.�n���!u ��;���,�wBdKtu�9���]2��0�"�+���gV�ǻ�ܐ��R=V�ۂ��j�j�-�´�:zu�ˁi����f���=xw�5S��WԺ���Ɯ=:>�:Xy�N琜��=9 ��&��zq�#օ��a.����3%_K�W~�+-��ʥV�o�;���px]c�:�O+�uc��Z���M�h]�/�c���<���H���t��ێ�-o*ε�Wf��)�Nt�w(t��oi
�`�eX�ޤ_���c��ԏ_ft�F��:Ȣ��r���̚=�;h4��]uK�@�;�kνty^f���s8"��(v�c�{s.*O����ި�JnMT�LԳ��T)$v_Q�w�tH�SL6��ùn�&((����x@�������4�����[Fֈn�"�ݒ��=&�;�h�?��n�C�ܜ�j:�2�u7����l���XZ��z�'��DD�֥,��*z}���_��U��3�k��^���	�51قb�5�-׸L�a����ȩ��U� �_�[ݡ��R��s��}>'8��,�5v�6�����t&�)?5ǡ~�&���+D�H�v�J���|�y|9�"��bsOl�F
B���r���|�U)V��w�
7���K����~-9K������<J��jk=�r�k�{�Cԯ���7���C'��~ot,b�0U��8���uL�^��χ� n����v3���n��@g�F�����~��3��]�I��UoU{�G����CY~%��C�gS$fڦf�^��ʌ,(9���k������_K���A{�:�@i��w�N��޸eI(��@�4�@�²�T�̇��}��0�I��n�</n��|Kx��ycV��B���5Nq�ôVv��ۀC�����bO}�[�T�|���9˚�o���%a�o5X��Ǯ�X^y6�*1�g���*�N� =��Q�C�S�.K&�{�W��	ܕ�\���0=3̃�6�{.�$V$�eWO�@�Q�o��m�!�X�8�*'�����V��י��+j\�����n���w���`�z↻����3���+�'l�l�k3�=s7��1�5$�d��Bu��4����M���^Õ���Y�K��v�z����?�V�w����	'Q## �;�9ȱUX1Q��ņ�`$� ��^7O7v�>�9�>k�����6cI��\4�yTe��������\�+��Z1B���N�Uxv)����g����E��U���N�S]�*�U�4R���O���ݛ�S��O=�p��g�"
;�z}��;Vݛ��E��i�V�f�W
���-<���2��W�?DC1f,�P�3���c��S7�""H�i� �-I�5)5(��d9�4��z�+U�����0�q�� @�ᖒ:(Q�csW̎ޡ�bL�J:��_s3�l\'r���eT��9Rjp	�z����gͭ������@|���\UZ$H�H��F�2�u��&~Q�#�����+E�pֲe�{y�]�2C`�$��ݾy��B�UFu^�f8�s�^��˙�h���&�o�󬯆ä�R�f��><W�^Hy{�c��Qs�gG��d��ӨWuDU�>sFg�x-�g'ד�$����v�.���I��tyo�6�3�a����m�d�Y���M�	Q� �y��wWi\w������9�.��B�� �E�"�� ,!� @�u����v�=���Ipc^�ʄ
ݭd�ң�%��X����7��]���>��J��1"�o��=$O$3 ������נa��� =|�2�^s\�^�D�)���#}��>gz|G��bG����^�AY��p5	5�`��<��c#��b��^�6�x1�&��"M*Y��7䖖<%2Q�t���\����!��C�4,AWԇE�=[W
/�eVx*�h�@����]�Ŋ*�X(���"
,DbȊ"���T���� �Z����XyG�� �5ė~� 
 DU�b*�E���J�Dc b<�U[��QU��|*���`��Ǫjk���}��V�-����ns�Y\��sFq���m>KR+�1^�FD���⾮�bv1$hf��
��{����3J�U�S!l���@y�.Ooo�����31={]p�������̺���`��n�����?L���~a�IA����>h�ĩ���̠��5K���:m-]���Bϯ�{أ�{u�N/FD�s+�ĦX�w�w������lBײ�~�}
�K�.B�[7؋F�; F�C��s�V���{x=�R�X2
,AE@\{��*�dX�޹��zvwy�Y��@�g��h�	�]e�L�o��s���鑻��3�`	|��є�ƺ�N*t�L{�X����l�DoO�-��%w�S{�&q�k^���u��lZ�gK�ҡ�Z��y>�ʭ�!ۓs�KV���K�fd�o�H{Q��	�cd�v�s'�����S�w�C�����.I��� �"0�o'����������O��ħ�������� ,� L��cƎ�V6a�j�ިƤ��M�� +@ H�+�$jӵ��7.�oƝvR�Nv������s��V�P
��YWs��U���/$L�B�.x��zwI�����B7��Dpm*nj��iV2�B���\|@�z�����<Ov�	t�Y(�Z���E#c�{="{D�)]�~���N�Ԁ���4s3�DÇ�
���|Wb0��6//��ȼ�L�~���$������BS��b�#���W1�f��1����d,Abo]���b� ��"7��aDD?i-�a���\��Lӵ���9�Ck=�v%�Gd䬨�:$^[�(BF%B����Kx�>n�0.c/���	��"7;�ܤ�h�t.{cꋘ������դ3u�!s��v SP�V�n�J���.8��-�l獙z&��y<��/���I�_��Q��F��d.�B6�����9f1��p�YAm	����5_�zh�(�[�W^����9�\�#����b��w�����d��gd�FU@�"<n�U�5Y.��\m��>!�_��|�{+%\��澵1�S"��t��<x1l�*��Bq��t�+��1��:\Ð���OL����<�ݒ��wa�xO{s���=�O�X���S����o??���+����,tj�|�O��HB�V�I��H�H]�♡q�.v;��BȄ
f�(�|��s�6<}�܎�If��ew,�X�~�T�EQ�" ���$<�
 ��1�g=�]�R������G�$W�:�2�+��z L��3x�*�ǻ�]�U������3͝�{��P�	�c<jY�^��[y�����W���| 8�{yo�S�����+�6vb�Tg,�رMXM��+j���R�d�zq��s/"��X#����2��Gf�g�
���L���E���/��qi��@�P/@�(�\m׵�������x+ގ���$���A�̧"�}�~7:�ޣ]4o��
ey_�n��|zg\�pU�!� �IO����Z�۪���T���� ),$l�i)m�$ ������dxQ��˙�b��(�M�3Vo��g�9�]��][Y0��ЩV�q�+x��ŏ 8;�fI%hݬ�1�� �Ŋ`�,Vr������a� ��9A����@��Gw`*g->��o b��A��w���`P�:�Qj�R�x�M�'�����Л��h^��x_̈́<�s�Y�cp�̠.
�#��5��I��usk���i�/5��6�3D%+$�7�c<�=��v�#""��"Ȉ�f��.0`ȩV��k{�y�d�����
;v�n�&e�b]p]��G�9�=�!��_*��f���x��P
�S{#c����'���8��U��#ð���܎N�lun8|�G�nK���%����d��"�Y����O_{��y��H���]�������ɛ'o������I���\�u��\�DD ۫�妷�#h.�ͷG�x���G��GM��d{�Z�����ni�}�+�l�e��|G��'ܗ-����R��b�b͑�m�OW����=ٽ���k9�Ö��.��[9��<t��S���I�(��F @�JH�����F{Vc=ƨ
�T�����3Yyn)���rWd�nv()�H���ʕ��m�F�e/o�`:[䒢U9e��{�}��BϤ*��7U~�+Ն�OX�\%�fx�f�$�m��<��{<�s<����랽r��t�<��=������g+�F1"1[������D���y�U?@>^���Y[[��+7}<.�o*Q�ےǦUuάN����Fq�I��JgK�^�~�)��KCXYP��_��%QH�[H
S�g>�{<�>�]��I�0�j�d{�Ak_��le���ZS
C=����~�@�zX��l�#�Yg�{5����[�*p�zdnR=�ϖ]�D���I��Y��r�zߖՒ%^��z���]��@ 4�kO^��s�z`�劖�Ɏ��޿V�<�h h���H�-�B�$M��*�y+u�oO<�qԽ�.��`�e�'��cI�-a�&@�����ڞ�f��#Cԧ!\�JaBGN�Nj�N��R$�vUx� E���fA2�4�MZ]N ]�έ�u�V?l��.�uMm��"w�N�1�b�9��԰���\�sۉe�QO�p,vG����٧�����߆1ۉ��o���;w�����4��Z��>�y���DPX��PE*#������T�M���:�^p��.�7�0��$��3��jx2H��2%+���7�}�=퓧�����w)�!�U�Vj��X�af��v���;������ԙ�+W���üAm���ӿ/Q<F�g�����o�\DF�M_MX=q�-����$l���^�04%rU�iy���~�GR���O��/|����G�,2z���j�ᾛ��A�"�w�Ӻ��d-#(��*!
ϲ�µ�����ƽ��`���V�����M`�����=<��z{7�#rX��t��d�������J���i��UL�O3�zzrK��	�x?K���ٶ3�d?Z��qck�M5���dak�P=��qK����g�	-�8=�Fz��\�{���@��Fx{9tѕʨσ�Ԫ��'S&��=*��wD��G�:���Yh��Klv��!סSn�e����b.����5>���/Q�{d��YI�ì��H*�e{'I�<`&�Κt뛽b��� ��H�c �AZ�	L"*r�`
0g*���s����G=����@��s��g6=�b��h;��n��ץJmt�#�s�u1|�m�԰�[�n �������5����vpG}�5�<*3^7��d�等��יUo����W�X������z<�cf�{C^a�8uB<�<χ�U/�f{�}���}+�N�����b�$�#&�mOX���R:'�Y4 �)�2�xL����%��co/�ON��8��>�n�svpb�~�9M�~;v�į�j���E�����+�����G���|��[5��'$���HMj���aFY�<����W�x�׹�b]�!�A���������;z���1��N��?RI!	$��I!	$�����B@�0�E��H�@�``O�HH@����I^�� $$���$�	!$��y$���k�d�BI��>������BI������_��6~�y	  B����� I�O���HBI9���?�$�BI�Op���$���g�� HI'	$�$����!$��LX HI'�_�����1�ɃI!	$��HBI>���$�BI��I!	$���8_��\��뫒II%�?4����I$�$��*�$���k�����
�2�ΕLN�.������9�>������U�қaT( E �HF�h�j�%Jؓlt @�� h)@�4���h�[@ R@�PP_                                       |�        ��[>����;�m�.��{[���{[`�ם��e0 ���M]���*��qgVm{��:j�盽��lҷ� �v�{��{��V�iO/x :��
��7��D��n���֢�YVo ni"�L�g{���^6����(���{iu��uU��{]� =�j�wu�O;��:�4H�k֕�5]�y�E.��˼�]�L���T!B�    �   �������7^.�ml���I��g�kZ=�GyΪ�gM�w7� ���"M��ou�H�kyܢ��Q6qw���<L��pR�ȼ �lʮ1�3V̉r�   ��7]���y�/=�URٶ׵� ��F�ɕ��f*8�G��Euy�Q�K�wW����4b�׀ ��J�nO��h��{ݳl�Qyb���ytw�(��˳]���@�         ^D�Q��:�t�H�;��ͳ�l^w%Og=eR�� 7Uz�.X���
���M^�c�<GG^��i�1=�[7� ��[.3/l{dJ^Y/^�p R�$��޷��yc��V�� w�mSm��獱�/=�Ջ^�{���[{�wJ�[G� ��k���W��=�y��˻��z�:^[׻n��*�U �         5�n��y��{kn��ݽ�,�3���z��s͌�� n���y��Umi�yc����Ź즓y{���� וE\��ֽw[�u�J�f�n�m���󽎶�� {u�n�˼�^6ovW��𤝷��ޕC<nN��q� ���mi���{��[Ƿ��㖛�Wl��m˄�{�tBI �         7���wm�����uu维�c��x�sݻn�^Yv�g�*� �ގ�7��{;�x�=x�v��ޖ�j���z�I�x uv[ݩ��P���ixǣ� (H����uB���r�I�^x �T��r6�H�ol<0�kŝ�<���j(�� ޑI����5���m���y��UJ���Ovҭ�.� �? �SP��)�IJ�d Ѡj�ʞ%1����"{J�OE(jdT���
U@ ��"�MF�  w������_�����`B��N��9c�+%S�@TӖ7���R*���T��B�R�:T��)A!��/?��=6�v�k�W;|a8 }�}�̋9�>�y4�e.mϗ��/���q�k�w��iG��*�|��	�/��Tv�/���Z ]��h��ʯ���ߖ'QЪ9��5���3��j�+��i9\�|z�IR��n���t��%�e�Wm�,j��'	�j e� n�{rA���R�J�]���k�ߣ�fI�.SR�5+����ɀ2 :W²\S�ݏ��y�i�o��y��5٘F��q�$�KC����&�|7�U��N;�ft[،��1����ި��[C�Yw�l*1o�t�Owkr��>6�!���\���J�Jj���8���X�8N���G�T�[+*(e���[��V+V�:�nJ���d�ʤ֢ЫӸV
J%�� �Y�Y�TV�͘p�!���ykæ�md�5\��7�Hre1mIx�d�ǩ��٨E�P���}��O��weZ�ʠ��!�b����p-�{ӎ�3��X-t�G
`[�%Z}����j�ּ��mka"k�~r�4&c;��jE�Q�UG���f��)ۺ�#e�1��D�
��̙����0:�p��-T�7b��*��M�p���ڪ��Z��ܳn�C9.����YT
�P3ƌ,���f#B�2
�yK���S��)�60`���^�5�*�'e�n�ۀ|/"��v��pim�c��$-8�d���R��hH�S�żj4t���2TU���tٲ�;~����9j�a�!ڎ�J�-��UݫCs
h�J�GnJ���{�1.U:����������l��5�:��cV���p�3��j޻���خ��Gq�7��grc�b�I�.^H�3���;�q�Y�n�s6�ٌ���9v{Oh3.��-e���P��ك6����:��h)r���sW��u�;,�a+�|aTs��1���yA^��bhxP�F����,S��N��E�,�]��.O+V��u�R-��ͼ&(�ך�|��6�(�ͽ'q�y��=�)ĭ��r����1��YM`�.���QfPG���C��Sf[���DKi�`5��b�໐�
�wV` Wj�$lHH94:�40ꘅS�3
��qR9A���b�u�^ύ���S%J]"����x0����-1Wz&5LSJ�ލ7a�\�f�g �	ۏp���f`�7!�p��Sf���L����e72*y )	�#԰	R��?K*k�%�)upT7y��U�nL,Zg)^�)��"�R;R����'4�QM��5�å@\%���4e�v�N�+/e^��-�|����k߰}G���.p'�6�_��@�B�t�U3F+iw�]7Z��mn]N��`W�[P�*���#{>���vK�z��V~��C��Z���\��M��iu���+���k^��2���̦d��|Q��h1�-�����u��TJ�C�]\r���QmiT��$+6�c��D�7R^�z!ȥ��]G�FŰ)"���;1�Op\�����٘7����eh�9@�j���e�rFҩ�iK�kkh
����
�Q�Ō�n�.ښ�Х����t�4�s�0n6��7/5��+U�(�f�wa�5�rp!\߫Er�����u𨀚��(}\(.�<��C�.����˙b'��Bj�{���Ee��`��)�L��T�*[�u!���.�Y�u�(�y���l���-9�� �췗B�����F^T��2�!��7EZz�h��ܻܢ����/R�ɇ"dE�Jio)Ic��*���sfj}�@q鉁>?�`Jw�A��O�<O�#���+7�ya��V[�
�Y�n�K!'��K*�d��n��]S�[�N��(�6��n��:����iI�2�mn��ge���.+Hr�7�3��j����;��M���#:�T[Y��c�%y	�R��٭l��{���TO��Vvc����G��B��u,陉���t-��d�h��1WQWW5u�٥[�gBͽ��^��u�k�Ɛ�-3w/r���i �Aϱ�/��oj)���J�8�ʪ��3����;AJՉJ�;N�^��z��	��y�q�f��Z�v�h�3I�f�Gӎ�6��2VH2Evh��v�c�e��V��½hR�tض܄��^a��e=�/^j�'-hK_mۙ��'���C�����5����6�v�r�Ω̟]�+��i�A�n��ْ��Yט��p#�!�R�si=��R��iT�4dk�x�Sք�h�c��r�K��m��RV�:�Z�8�,�7hfhǄ�Ph� �j��Z�v��M�,Gk�(�n��E�L̳Yno�*�}�aY{ ���oC�-���n���(֒Jaf!Hs��7�iVdL�ۜ8�6�MK�cO0�; 5��s�!ջ��;wA ����ZjT�Pl/t�O(��@fߍ�+���`�(��e���h".��l>�|�Lǩp�6q�*[C-<���ݩp]��ljU�N�)+���AՐi��a���o`Œ�n.kj,����N�v��Th�ɭ7�]�;��8гr2�7�?��pA����pc�n�[�)V&�H�oAVkB�	M�m0չ�1k*���R��-�ĥ�v{��։<F��7�e;��qkI�Qb�lY`��իKf��S�n�B�� Y��GZӷ"�
�]1@�����f��r�3�X.7f�����7�����:�֗{�+�^J̏ڷq'��\[��&33rfg��>��V�)� ���T0��M�J%C	YW|�ȍҜW@�R�.[�l����_S�(H."s��!t�.Y��ۧy%$�6q�[B�;CEk�|bRt]��|n�8qDK�z4\�� ��F0�6�S\�uf�;�u$�[DV=���7[��j���R��~+##H���s�@�Ƅ��&��hr���Q��(��t2��̣����>P1|�r��ƾ4�
mP���t�X��>�Kr�����<'h�З4Z���*�$/3���E��J}�P��jɸ-
�yK�M1��7�L#�Eg��;d����co�!�p1�f�P��ڷ���׹|N�6�1v�����qu��%�-С�i��.�,Ή9p:�q��[vIM�f�=S,ǃ3�k_|V�R����Ū��>��P+��]��rs����߶�b<�����Ji��BN���F���:����غ�ɭ�U��,͏H�q���-�A"K`��q_.����7qUXP�iw�3\�9U��cx�&�Ap�f���[�D�zN��I;�(j-����6����ٛ5P�e�f�ʇ+fR���Q�E��Փ#��i�����؛˜��-탓��q杳�st��n�&�(�Ȁ�ۄWh[�����X(��.�(EG�r�n��u���rб��ӯ!�`X.�e�
:l�Z6���Z$����e�� )�uK�(b!��b@\6���gK���A�Ibu���nn�Z���+p�U�u���򢠕�{p!cv��oc��z��v�h���X�[�ձt%�����Zv��@�:l!��̼�n��3������U�6�]��pˍh��i��ۚ�t�YKF-�1R���Mi	&���*���I`cTŗF�P�r�8��`iX�a�)+ 7B�W1<@kͷM&����d�%�wZ�@o/E<�n�%���f��tC�W�(�Y(nKl�)@��E֫�o�ʴj�'vC�UҼr:�[\�<fee�Z��,�wz��2�Ǻ��ȈU���y�����^K�@f�@aVb�<{�+S�mKˡ�L�d�Gn�\�*�u��F���Fr�,e�V�K��K�7,��f�L;م�!G;m��,�n�S�KZ�N������`�PH�%���3=kS3
����mf@N^U�67�$���٤��N����vc,٭؜�5ˢITnԢ����Y,�}�2�n��H)W�^Y��B�[c5�T;[V��ǂ�;ـ���IC+V��V6���k���8K��LIm��y�4��Ú��c͛X72�Lp���Yۧ�[2�X�p��^�p=� M�Q�ڷIJ�;�ȻW�X�[k,୺�)�y&e%j���-�ZS�׆Hou]<��vm�� ;wW��榎P���ɵyY���h��0J�X���w/�v���l�v�h7� O��@Q̒�ת��5=;���8�Ǎ0FhY��Ѽ�٩�2L.]�j���Xi��I�*�fM�d̓ �Ј�d&� e#l	�O]�I3`�aְJ��V����qY�$e+uyS��0�a�J��A&
���fQ��aV�ʺZ����=����0]��S�oa��¦��%�,���X�4)����L�j���%�2I3��Փ�yt�QL�>��Ih�6��&�V�4�
[`v-YV����ج�[#sm�D1�l�60ip�f��30�a��	G�B�Tt$�B۵2kV��*ar�3'3S�!)�*��>uH���-�e��*Ⱥ�R��u
�(ɍ}���L�C� j���M��s4Zq�FU�V���	�|-8$�U�[�!#���L�kku������h��Rt�����ʰ�	�M���͗���;���x� C�=#N���"���ڽ�s"�>[-c��R0�:��N����C1mvkWu��f�[(^VJ;�Q ���f1�n#���X���;F�]R��o"n��uǙ�*�M�i�'췼�U�=8*��	k����L�`�2��fe�E.���L�	i�� J��/�*lݩ�����]�c��� �b?�0^�MVmf�m���=������n�;du�o-J, 1���䦁
҄�غ�y��Ғ�a�	���������1+0��x�ZoQ����Q�����5���Q's���2�8b�.D��.*D=���H}�heY\���ٹ�k�����Z<�Z�u�-[�u��g��{��Fɔ�+��|�7�dsL{S2��K--�n���̻��+B��`���Y�u�%B�,;�/fCI!c��X{�e̳%�ɹ�.�T�HK�b���\7P7�y�6��ܦ��-�"<���A��
-��0k�l�pZ����r��d:�8�
���r�
̸�\G�b����j�LL[gm�S��@ ����sUc��*^m��3w��Òʵfȭ���{��L����(�{���*.
�Ջ ��i��b����1��Y����,�yg��ܺ �vy2|�2H���'���V~7hk�+]�Y��hp'wO-�"�یa�ZQ��QEuwH���"�0�,�>h:9UB�Lg>�syQȵ^9�4�p�4�e��E\ۻ$��z�Y�&b_����A���n�&R�!���\GA��#F�4��n<AܥWCH�ad��v°\��m��jhא�wB��+t��RQ0a̢X�#3hQ�,�TclS.�j��4�\K�J�e���p?��fɯ��+r�Ǽ��+����k!�;�!FAj�t��+�Hd�{z��<�9yZ�Pn\��	QJ��Y��V�F���fY�{W(!�j�m����qrK���v*��T�.!Uxsi��H���3$��E[�-:��y5:|B�b�+�s�Pe4�;�1݉��!Q�/q�͊�X�-���e�n������8��G`�(Lk��JS|̎�94k�����u#�uٙ�M�x1��yt����v�$��'̫�.��)�`�n�I�b��Zk�
[���YwZ���<�bL#���iD�U���w�������p>�5�~���I��70_,1���C�VF
v8��e�ؽgmYu�	K4�L:�U�0���Y�/"�ӇP;ռUZYD��j�iF���@1b�{�'��S^����og����V������U�����e�q�}�}����b�t������}{l�\�(#h������JV$��Y�ֈ;��w�=���x���wWXn�#+)8���;��Ⓓ���6�I��k��N3F��M�$.+t �N�J�6n���on��٭I:yEf(ј���	�y���M�+4 ��ܠL��ŵ�hk�Gd:U��х�wi�-����]#�ff��`�5���ŀn��ln����(����)Ö�^�̤�������Kc�n��V��^dW�v�w^^iT[7{GR�/-�fe
��t�g3Lv�`ꦐ��q�E��f
��-��)й�ie��ѷ.�4�L(a_	��1Z7J�/U:�8]��|�_n%_P��ٻ]�ʫy�i�s�I&���c�����"�-��
T�+k>o"��+F��Sk���)����z.ᷝO[�
�Vl��7�ni �eavL[�u��� ��2͓Rލ�.�qf(L�s_^����%nfF��#��MP�CM=�ϰ<���qӇ���ګ��حr�@�ϗe��YLԧ%^�
cO�	c{�Bd�-[�5^\���^�	2.��]NZT:���PK���S��4�^��;%k��7��H�<�:�����X9��E.ﱷ���Ub��t�(��YV�%�)J��4������٩�N�$���p�s��XD�P�D��0�!��w���k��Eh؟�[דGb�7%)�;��S���2��4�䘴�g���7&��g6C�N�Ҳ��������\��PlM�����U��t�Ŵ�n��m���GU��1�1��]D���q*��d�� �����QDƢ��7���b(����b��?%n�%哆Ʋ�7����o)W�y�yӯt�9]��[C%|q'�e,���*�*���>ٙ�}}����6HN����U��՛Z���UV�.�
@�.�#���iQ�h��Wv]�H:�Z+�D�4�iX�0�v��Bfև���!j��'v�ʹq����#�{o[�ES_l���u�6�@�g\��cAY�;�ol-:u�0ؼ�6I��(�;�6}��n[�As�	z-J�	$�I$m���Zڪ��RZ���UU[UUUSj�Ԫ�UUUT�YWj�V�
U�*��U��V��jڶ��Mm*�̫U�]R�Um]UUAHURdj���.6�`��k�����Bj��( lV�J�UUX)�ٖ	���uJ�UJ�Q��T���(+U�Vv��ٷi�d���,��nGns�s�8z�Vꪵ�*�*�^���L�?%�W�"���^���檦��q�X8� fn�&�u�u��ZU�U��@j꭪�ꪪ���A�o���������UT
��`�U�����ZW������ @*�K�gN�U@UmuL�;=�5r�U@j��]�ԭ c�j���w�̫ꪪ�ڪ���*���]�g�I����:}�v"n�ݲ�����#��<����u�v��mJ:�g8F�Q6�w;��cy7.[s4���\���<<m��h�8�/�Qs6͢���f���b���J����c�M��̼�k��tu٬p����g���q��9;{�\m��l\��0M<8ͮ	�3��j����<���HE7Y籰���9n�n���\d"��zA��ց8^��9m8�N���d�lm۵!��K��n��{cs�)�V�i�]��T�^���ew\�v��R�'[��#�n=��ap��
���hN��[z2IqA�4gOZװuQ��t�އg���;���5�a���m�v|���{�C��mu��{z���#cl�Z���㫎M���ܵ�Ɯ����wm�a�s�����Zᳪ6WΗ�W�۶c����q�6΋9;��\O.�jݰ��;+��Ì�A۶#nu�ݺ�oF@u�-scN�y:�C�Ÿ��rFF��G�������Wnvy}��>BøG��b�m���}*4x�m9ۭ�m��i�<�m�ɜ�d���pn�3�;��[�j�����C��v��=�'�=�y:��ܚ�,P�8���s��uy�N���g� ��O''+���׮�筚檓2N���N���٧sv����iٺ�:��y�w��p�fom�PN��n'�c)��<oJ�u��=�v�n3V�;��g�?;w]nov}q�a��+�vN9"�0��=��j���qk��y�l�s��n뱣��N9rm�:L��t��[b�έ��G#���'A�����s��l�qN�{����������^�c�;x{��'n�[�۳�t�F0����m���#�}�}���~��0!7�Wo+�����rq�S�g]=�H�m�Ar; eŒ���q���Iב�l��n��eۢǟn�;)<�䐞�G ��<ss�]�U�xn(]J�m[[��|�ost�mr�\o%�t+/guɣ��]a�T�n�Qۄ�cX|�ʨ'<q�9ƒ�wl6��[���β����=���tג�rr�(u����⮓����vKĆ�a�7l�봽�Fwz!�	Ư)��c�e�A�Ãc΢��=���;�\��u��h�\>{l:��&� �<��lea�b�v<�:��7{�X�7<�v��y֪��_=�ڣZ��𻮄]����v�r�{
��=���8v.{3;H�b�l�����ݚ[�8w^x��L�B�\R�*W�`�vwce�7fJ��ou�z{EۡG��a<�������u�v,{=�nٱ�/d�$����g�ǳF۷m�!�>�1]��u�ϝ5m��R��e.�C�q՝�p9�{�\;�֩�h�kkz"u�/)�̹�ñ����;�x�r����5�������7dTv+63�f,uּ�J�?}_�ñ��{&�g��0��+N��.�͛e��[n6�N�-��z���\�1{�;lbݍ��<�'�2�q�5ojQ���mF�.#��γ���w.��=5�]u�����3�<���=��6�-���lw ]Z8l�����l�����v���N�Gn��&r��M[�e"����UD���S���X�k�ݸ��/,�9��{�`�iP�Lóe�n�x,��5�<���sضɕ:Z��:�=]kf��ܣ�ð� ;�ֻ=ȕw`�S]�lx��]�:�����W�n�n=r�;��Jn���;�[p.y���#s㰻�x.wC�n�us��4�<�l�]����uN����� P�<Înuf8��.�7�ݨl�6��>��k��{ge9������s���c����[��6������n��������tU�\��㊴�kl�Ӯ9wH�Y����6m؎&v�Ƚ�s&�B��
)���݂3��юٶ]\��xC�5�:�Z3�M>7k��Ý����|gaO�\"���ylE�vc.�օ�yƫsqv�,�v�w\f�t��X^�m�Y@E�:�o�/d�Ӻa�W�n�J=Fz���<v�m�p�#�vE�d��b�w]5˲���\wa��2��X�p�n�/��Jm��=�]�`��GgշW\�ۀ��3��9m�v5��j����c����P��M���qqfxx�ݹ����=}���mF.�d�M��n��On�۶�<���m��N5'$t���b���j�vv�����ᗖ��v�ΉJ�l��%G�V����� bM���v:�gd�t�����m���vݶ[�^�&��MD��c���m�y�'l�l�p�-�s�r������>[e/e���n"ఽs]���tq��֮��Gb�����;�]��7=�1\�0x��unC�q�۷Ô��r�k��9݇v�����a�5ʱ�w1�>إ�@q�q�qwT���7�{��˷���Psv<�2�8�vvS��6���`�nprqGE�.���������7!�;dxݭι7N��CV�U��]��c��[gcj��m���fy9���\X|��gY��v�^�i�1lò)���˫e�!�W����A���hS�&��t�خND���;�D�}����O��!��uj�Rd{<�m�V��+��m�;��ld����9��u�P:3��pp^k�`�����n�Ln�ݽ��[`w��F��u��2���c[B\c�ca���Ï3sM�8�����&�V` 5t�z�,���<�jv<J%����$�kY�f�z�.6��_;|�`��ZW.g��]�]5���֛���=�U��Y�d����Kq�[i�fn��ï�7�.���u���0�cm��o;��`݌u��y�<�{j'��z
�ޱ�le�\�8�Ǳ���4lz׳��;ë�<�{1����;6:�
�Vs�n�rm�#�ov�]Cۗ�D�o;v��Q�Oa�Q3'dx�oV�g�tc��qcu�g�&���\��6���C�r:�v�5�o�t7N�l�|gI�=��x8��أ'�v,m9]�����כ'�'���w�){q�91e�n�8�����;#��-Rq��p�lr�.;i�{�hz�ۇM���\<ݽ�Lv�;q��M۱���k�N�x�^_�ݺ��{m��ZS�G��}��豶玣u�-��kY�Jy^��q�ׇ��5)�v9��*�1��<��cu��|�)�����s9M]�?�p|���Eݐ���� �V;2��4u�\4�:�]8d�u�KК8�m��$��!n�A϶򼎎��Y�>��V�\*��(���ƎE;rpm��t!��j0Y	q�s�71�G��i9�.n����vw�v�s� ��h��d��[�.7�sV3b�p�+&ʋ��<��������]��익�H�`�nB��%ع����lu�g���o]n�;g�v�i�[-��]��(󻋗�sĜq.���x�[:u�cokWv��8P�s�t�G�mr.o���
�����n�����ћ�;uT�m�p���������T��i�{1���nu�<��ƶʔ��8�u�!���Z%eB���A�3��nP{v��㵮��	���۶�<���n�;����q��ʻ`�n�P�X�b���kF.7�Ȯ�ɷ �dS7Wl�d��ڿ��c	�|e�Ϟ��2�u�i�3k�'��G'7�׮�}]8��}�۷�r'�*��
���d�Nwc������#�y�z���w^k�<���{;L������ݺ�:"�rm��'v箽�C�[+��t��Y�+=�z1Ѡ5�7xt�6�lu�c���l�uj^5�8�Df��8y��Ɏ<�p�[m�X=���U�v��ٶ�z���8M�4��ٰی��:C;v��Rr�첷t���㋭�v,��,1�$���_n�n��*�����ʛ�f^��
:�3�ms�ݹ�� �>n��:{V�nw��& �� 8u �����#�F��Y�:0�cW]�6@W���lM`��vLW.E�]��lz{t���&஻-�Jƞ�v���.����[�;9�F	�۞�b�O�=�q&��;�q�������@	k��:Ň2q�����V��/\�<6���
�0]<��9ջ�x^�v�m�P5۶ܗl�:�W���p[����k�*�lm���y��{u��w��5�Ng��nl�{ 3�t6�mkG6��/]8�G����\n�%>́Nv�'(���0Y�[�h�yX��Oz��v�`�ݓO�������~�&�]xA8)�NŃ���<���b����om՗�p�4A���Gn3 N1.��=�Y���F��U;y۞v$�b��;v���c ��/\���&�v�'��e[ٸ8�����nlͬ�v^p���t��紉i����wN��k��V�ݯ.��q�gt���#x�[m���0^�������A�u1�ԏbz�tG[	������Ah�i�zP�:6�����=Y,���󺫅�L: ݲ���mGawnE�.��-�]�c��.Ӷ8�l�nqh�v$s��\�n�-u��F��u�\2�S�OF8�ó�ugM��'8�u�2�l��ҧ7g�ڑ�;(��r�1��s����{MӶ��7�g�Ϟ��9kcm�;n����+��i���O`��B 3�Ƙ�8;��pV4X��S�\>ޡ^W�/g^.�6��;������d�ܹ7\�� ڝ���{3�Κ{v�u�n�X;g�P��_q����Q���;p͵�3;�7hN�^�E"�:�����k�.�@Lr�mX��t�Z��9Ŧs�Q/l���B��Ԥ	�D�7�Ì�9�1����Ԫ��{>E)�1�v�sZnָmb�()�����+dg`�_.��2`�6*4,� R�U��$94tg�%�9��A�^�n���`ȗ�=R����pbosu.����{�l��zϟ\>9۞ n1��k�0wlq�����\�7u���ۨ0n�Z�Ca���<[{!��8���y�.��c��u��
�\��wn&��>ܳ��aؗ��hj���WQ㚳����=+����۬4��р�nK3ɛ�ێ�Tv��!�vGq��	�]@�I��1�O�ԗA�Z"�}����{�'��\�m�q���O F3�D�f���y/)����pu�˄�ks���m�q�������n�9Ϊ��xT��ll�ø�&Q���2u�g�vX3�8�r]�T�۵۠���E�X��<�vw;����L�]yx�h�c�g��%�Hn8s������������{��\5�ϸ��/��Mu�����3E��M�,��qY��ANDL�S�is������wݻaF�������s;)Vt�����[�g��PV�������.C�N�p�{(���-��g�c�Iݭ�Zr�:禙�W����F�>^��x9W�<vSqs˸���G���y�Z�a��u�N1Ԧ:�Y<N� �;=gN�Ok��q̓�t��c�7fޡϣq�W�v�Ia��8�4��s�=�q{q���e%)�glP^0�F�:5�V�{[n��Tc�;�����7�����*-�ݍ���:�D���������N���a:�Ŭݻv���]v*��r�1�:Au��V�-!�n=�.�k;��ݞ�8�L�3[hW `탪w"l�s��GQ�������ƞ(�z�����mv;����9�L۶�á�y��M��0�xו�"��5.ڌ��vx�^V펍�*�n@�N�Z����7n5���%�<�Ւ���UN�@�9��/ay���\Z�qٰ]�8{nNn���z���9'�^�\h{���w{����w���Z6[��@�ۅgы����Wd�h�ui<��ۗ�F�86���Vֺ�����qˎx��`������9W�ݪ.iܭ[X9�]z�:d�m����v4e�Ih{���N�yx�r�i�.[��S��HKZzy�u��wkGi�����;�)�c���vںN^^F�O���\;v��{1��ݪ���:��	�ֽ��4�-���{�Pn�qؐC��1�d@���ls����]��p���x��Ϸ&��f���E?���!�٩V��j�H�0ք��GT� CivkiJ��U��:\'��1��#k�����?�}��R"!�D�Jf3�v#��d?>\(���Gc�ۼ�Vl�.��|,�T �<U��E����7�f�Aϵ���س&��@��p4Y"$�r3��Y�(Sg��`�C��*�Wq���ƫ�1u�T��l�mdk q1���܊���X��D��h���N*~����ioִD�qYl����;�f��[Q�S�y�������UX+&a������1���qY��]u�-�}z�A�£:��Ĉ��dK�!j'wB���(�,�Y�M�͹:��\�C�"��@����#���w
�8���':;w9��ńc�FL�;��P�u�
^]�w��G�Yj} hI#h�ҎC�q����g�o c�����ח���
��u;�zL��n�Ǥ]�so;��~B���?k&1��>�����z�ٺ<(�����\�U�B��Z+��8��.�.)�f7g�[U�]_L���ɽβ���P��ν��4�ʷ����ݓ����u&(8w��\�/fb�`�+�7w�V�"mR���c�V���\���W���Ϸ����7+T�iq㘉s�Kx����AΌ��O�9N��lu�DUK%�K�i�5��gG��+�!I�vT����W�٫,y�`�x�`@����(��u$��{��&�����u�=�cV2�E#w�y	�fk��N����R�kt�Oc�*�Lr��k���r�v�;W�6�FMԸΔ;/zv���"���������9�&�-���\n]A�ތ�͕@��P	,�+�L8-_8}���{��i�QZ�E9��Gs�P�;~��w!e����(`��c�T�LlV�E��6��qc��<C=�x:퇻	գ-@�d-�+-33�μ�".߭^KnҘ_n�M�M�����4�^�ˋ���"��	�يb�;��Ai��EX��X�ݣC�\14���HGN��ו�k�8�Y�j�����������f�m:衕<[�����#j徺r�D�|{��q,�!v�}Xx��I&�a7���=y1^�c�;P}iۅ�{ΗS���gVoxY���"<����]앛tt��mWW��Y�;���� w�������R#1��)'dWU;ehy�o6�M{t�F��cTvaؚ���5���D�"R��I �~�[�s�zOhW�ջ��#��Vc�����4�nee���<J̋�MI;]��� #-_z8��]u�6KE��ݚ����e��o��^��d6�.g~�%�I��G)�xS}xYܧ3n}�i��p��J����dQl��蘠�q���X�Km�\��˕���76�az�c������6�B=��*�sE�_o8�u�egP�m�
!�L�_'2����A����U:�����OON��Y�ؠhg͆𐊁9���kvZ���gI�m�4�Bb+���i��o���с�k�W�5�n�k��./������ߛ�p���+��QE�&�`�Z�;�;=��}[a�j9����$Y��2C̫�M}\�(�&u u#��
å����OR�0 ~��#1��\�̻y�`ćr����x�1a	�{�fӇ��XXۣ��hW������ֽ��Lގ�����/�vΫ�,�5�۔Zʽ��:����z�F�!׵����XȎ�N���SX��^f�$�y�=(I,��RUT��F��-%}�\��]�t�����uD���ڲ-�9��j3J"z˸�CR���yR������U�$��+�M�n��q�g�����pz uyn���'l���GIQmN�hQ4J�-�ܳ�Su����T�M`<��f�Rވ'��d*��w�LΆУj�;C����V$w�p�Y� ��pr>r,6��U}�߻�V<03�e�XC7v��J���$I/�o���t����zHr�̱/tp�Yu��S��'pApr�UN�Ru
	)�ЫO�bo4D�\��P�FUv��{1Q���v�;ۡ-�x�8-�0ݢE�|��EEL8�&f�n�*N﷜0#�A��ʛ�Ȳ8rی{���uL��[�_r�Y�^�,J�)I���oQ���`�C(��4n������^�=�9i�]�!�&e��U)3����Ņ�#���ݎ+��{�wr{�����Aɲ�|v�c鷗��+'ƕt9� $js��܀XE�_u�,�%dؓ�t*_1�4�d�+e1�}�]�l�f���0V�fz>{��Z���u�Y���jݝN���C��S�8⸭b{GB���E��"�u�|��-z95�nm��� �<��v���y\�2WX�uq�׆��L�����J׵�ք:�m'�s�R�������Ggr�x`�n3vUvN��t� nzn1kڰ.u&�����d����[\�^��;p�6wF��׫G`�8�GN�M�<��.�mɺ���n�t�.{ﯺ���K��[��Ǟf:�Y꣫�]�&��{ei�%#e�#,�%P�����Yz���+��!�Н'�r9���K�1�˜�f���ft����%w����(eܵ��|��5��%��.I�E��:6w�=T8w)Y=}�^�R�����Ou��_��ϴ��~][���𞠳5��j�m��j(��Ә�Ӥ��-^��`�ump��\-�����6#÷rG�i��-���`���B	D��9��*�
;��w�;Jmm��l<�[!�L�ڵ�u��j�It\�0�ʏ8�+�~�$:������[j�{�z"m�����C�A*#�Y��Spb��U�nGXh��\�,aʨ���%A�Dhn�h���9���{�ۀquY�ZM�`�:�t3��w&�2�om%���y9��%#�Ɍtg��Ѵ�N�{X���H϶�v�Õ�]ɳID��ȭ���ވG��q�m!qs�]���Vv��EM�z�?�˧�l�u�sFu��s8fs7d�Eu�|�}X����m�H>��r�0�;WZh��>G�>uʘ�;��R"o2�}���*u�vR�����y�$���O��]�J�[	�$#N(�9j�PAw��]Rm�Ȩׯ<·{�@E�7DY�Wp����͌0ؐ���Lh��-����;�4ͳ�	3��y�����n^凈����A�^]�p����(�{[��s�rSg[��q3�Yw�:�/~�O�T�X)��*�p�=W�'����
��ڼ��d��ǔ�>��s��P?PĽZO,��D��7�	��]��k���[/٪+\\�,ei5)ڱx�[:S���l�-\Lb����Ϲ���V�����Jh�v�n�c�흆pw�3+��)��W��}��;u$h���IN��<�=���{ή*���T"�Pù#Ĳ #4����[���S���K"���g;s�͆B��1#JT��5VZ�����3UN:����e\�Zy�t��潀R�t��b��L�ucT}/y����C�ڵv��*z�nY|m�wT�Iռ���n���|l���Wnc�"��ٵ.{�rE��<�7����u>�C����܊|�nC!-���3��i�\�k4���
HWid���V}��I{/ʵ���V"��5��[��H6�ά"�-D�3*`&D��T=���ܹ_s8*���Prj��gt�әM]���!�z1N�b㕯.r�}�6h��l���H$EW��h���j۫{e+�竫[�ش�=�N�N��oUe�ɎF-H�R{�Ųv��r�~�{6��]Z�3�s1��*c��}oW_o��P�Ww�����q�Ӂ�#���b_$�zJj�^����^�J�6��Vfϝ�P�^w��ѓ��uu��:�j���/5�j�$l�h��Gm���=t�{��d^{��z��n������}WY��[s�j�Lz v��<���q�d��8�	�c�����D��A���{���;L
�;Β��o�1y��:mc�繣n�"7�O�y��e�Kb�m]�9��r�K����8�R 4���T�+Ie�e�D��8:���p�yA��5����l�uʆ�L��b�o�o��d�"6�Zq�U'�/�֘�h�g_@Gd�v��la��r�h��5�(�bP"ehx���Z��t���������=I>�X�9Z��TM�;%d>����{��{6^7n5k;���*�}�X̓�́�˗�j��Xв����*$X9�5�Ḅ.y�}��eک�8+S���� 1{���}+`�f��������}x5�e������R�T��yo�䚖v��~��f�Ey��2�|K�+�`��J�B\{V��vmsm���9�{�C;ꅤ��(��If�!\�l�.��2mu<b��ۄ�w}{������{L�1ػ�t�ϵ����]Ϝ�X�2$m��q�����]r�T�����plN�f��Ὦ���:����J��;���f��
e_��r^f�ߍ��1�r,Q@��{[t�f��*?a��>�V�3��3V�F���7{�9�n�֩b��i �ö��F']�炡Ck]�����ְ8�����e�<W[��uc��m�u�k�����㍇�Z�K�c�F��\��,�Y���ⳬ��E-ǋ���t4��l59����H�Bkcy8���Z��c�lۋ��u���<����v-��=�;\vr{/+Y��m�㿓Y�9���wBF��{
�v�+�Uֲsu�޹�z���]�Ǆ�][�Rl�|w�|xv~���YJ���u+ōV��r��ɭ���;��ިؠ�sַ	���7=��M�o7U\J�b��^}"�ye�Ku�ҏ�,��:��ݵb�5�r�a�~�9�v_5*���Dr��ޠ��wY�q�]K�*�f�; 6��z����;C0]	[�i-̘�������1�����i���:���"9�L��`���4pg]�Ee	� 1�z���ٹ��-ݫ���������+�z%�Z�Q�.2��n �%�5��
��wu����$m^�;63*��˱�3 ��pY��.�7ҶV:�t.MQܓ�n.��j:�q��Q�T����e]���whRE+�����_@,=	�9�k��f�:�ܓ��k��e�ը넡[��UK*�����z۽�b�#Y7˽��7{<e:;�q/�aS�-�8a�.np`z�rP�v%}�ى���}�&<����S�vV�#���+��sG+K5���Q��F��}Aݬ�Y��B�q�d�2�;�i��[�����5�9j޲E`en����Y����X�o����x�������s�4���dُ����Ќ���mF��^��pw�%8���]~���]Y%����L�2��y7�UUh�ٲ(!!�" �Q%���$|\�Uܼ*��;���c�$���heLa��̍�<044��G�Sڨ���[���m�a�V�0�dqCF�5�2�K˅��,��n��S�
���\Rwl��ײ�C��V2����C�ٲ`��p9�>8����S��](f�W������f{9��+ݺڭf�GU�1�z�E�ޛ��g��g��~���]�fJ�9��жT��(����V�ĝ��~ͮ�c���5�	����e�!�U�:gz��//�5�B��x+{�iޙ]�ڮuЫVr)��0v�r�A����CiC(~�mL('��J�&�������{����1ʪ��J��~��\9�m�dj2/�b�'F4ǵ�%��Y*��j9uDŷ�U���TX�`�Jgī�ec[ho��!���\� ��rCvm���N1��M	E�h+��ju����[d�+�l����T�����k����l>["�($uъs�]�����u�L��At��r���\řz���K;�!�j�u�_]�������b�.��Q2ݶ�k�&("rD{sxҗ�
v�Si��!�jt���[Ը\7|$�K:+�Xk��!��؊��e�۾��f�Q����s
���R���cW�u4��� /l������k���P��P����Û8�M来��(Q�������"`�t�g������8|�@j��k���6��+��ȷ)v5F�:����G�˙��/Z��~�}钕�P�f�&�}�����q�3O2�y�[�&a�r������G3�zfbNwӴ�,lC`KW��m�C�.�*���:#�V;냥g�/����Q�he�U'zl�Z�y����D�n�������A�����\�<�out5t�g��H$���&�F��r����su��W���;���h�t����u���9Q=xz��/���JW��EI%IQ�/��e%�}�vK���52�8�n-9Rm�[�-�N���[س��&t���g���{��� ��[zɷ`�����5G�P�\P�m"w+#U�3����\��6�+R(X�FaJ��ۖ_U������훞��OP�XE�=�f��2��5�5߹���B�(ʋ)����M^}$ZQ
���~�o#⁴�6���}���X_�M��#=�3�(I�:��F����=Y�z��qi|v�D�0�������Q�"Y-�X�Fb�˶#V�

��b�ڤ�����(�}L�߮�h L�J
8�p��������åd7��8��;�Ȥm}���q����[��ّ dm�`�`�>K��C�uM�1۰sA�;Tkq�6�,`�i@��
4�ae��&�禯��߉���Bq-^6~�XN��[�
x��|�b���~������=6ֺ"O��=��̬Os_۪�fȃ�9�0���KF8�L���#~�fZ�}���X1��ҹX����'S$�+TF��L4(�,�Q���qZv�$���0Q;��w��ºf���l;��tnox�j�3�h�u�P �0H�R
#Õld����#M�e�Y�vw�+_0mz�a�����HxR�[z��:��p�Z�W�8���o�#�b�e��I/�:l��in�����W�(�Ү��X��)�g��W�zhV�A�.!b�'=�4+��q ���^7���]�wQ������;�l/���$fa�7��1��N��`�����2еa��qD��M�M����pk�"V޺�Qy��.�W��%
�eR�ܱ�u��<|��=�`<:�"��"�ƶ��u膝|����&tC�\��Қ���m�3�>��F�:x���LUґ	��t�D���^9�}��劉�<P�/6�*x{Xm`룱i��s Y{�l�eӫi���x�D�mkG��JO�:�h"1�N���ު�r9��e"̑�f��a{T"��[^�8����_'����XV�����v��VXHꑖ�.�	"8��8�	m����ˬ��O�9(�Ѽ?l1�ާ�s�����ŕrM_Qdߏ���t�K�x�|��5Y~6�~�ϼ=M�����M@�ؽL=��RB�I�����d? �@�9��T4�N�z��<�>{�t4�B�/���]�7��3O��
�"�"N$.�Ǧ��#�8p����׺<#�̑FdmH�,���Q'��L�:a,x���s%��w ��w�ʧ�c��W�=�iC�
��dV�{6D^��R��g�%ybz����.��,�a����|������C��cl�ҭi4��A�mN��ʯN�V���������36P�E���uU�z���`�+#�5X+Mbԉ����1��o<��%�Vf!Y����:�ˢy����U#ᢈT��l!�i-�����4f}c�R���۠�n�c\�(Q��6�H�"7��v�=N{k �g���E����pv�AI�n�q���ڞ�c��cۇ�G���ї�'mtm;n��Jl�l\�ܦ�/\gV���ݹێC���玠��zݚ0]�`�SX�u��c`�n�O{>v�����4r��fO7<��z˳\J�8�㣀���<w�a�>g�<nW-WeK�P���ry�͋��쳰۷���ƻ���tf8�tR]q��%�m]q�iE������_)��%�v�Z�T�8d�8�P@���}����I���'���*��ҳ޿�u�����ځ�LkC���W���9�t��L48��G����]���#�`��"��� ��2IvF�1�dC�g8����Ӌ|}"<���#��+��#��4�S���6"�g�qp���+Ӏ������i,p�٧�!�X;@�M��_A?H᱇�#�����g_����n�Y�B�!�o@���h3�I���͛5>����P�����p��By#����ܖp��8�5D,4h�D������2�0�fI7��S�k�OL��G7t���R��$�ȃ�޵W!���,�T\Vxݳ|��W ��k����dU�=��G娵fH/��%� q�XZ���i�}r�Y�M:sV�$ut�a/�}��Ud�b��qb�$�XW��G?*�_qazj
d���H�D��댌������=�C%;L�n�(H��n.�u��@]m�ƹ{>ј1ƞ�]��n����8���bc���y�{�u�lw����(�X�ԢD�g��R�(��\F�������V�"��q�e�0N:nn�@���w�i�����0��N�I,��U�?���~qk�p��{����[���-U;�$�Lm��X��'[j��F���t��2�E���=�x�ɜkN�ǖ�\Z]60���
�����z�X���>�N:�6t�J�(Q@�)�;w�44��=~��N���x��x�0�	%112 ����i}�!"Zc����;:>���M�+�"��u&,��gB�ّc-���-FjD_���}�w���>�|?a��RWP�EV��KE�[dWV*��	駏wF�y���Yr�?y�Y��I��i�s���f��3`>�tW̳G9	e�+�3�E�]��s�٤!>H��H�W;u��x�ģp�!@�\�;��ڸ~Q
=%_b��:t����h��%�+n��xK�xgtW��IÒ��>�`�Qu�`�����my�Ȭ̈:B��,�h#^�<ǝc¼��Vm!���bQ݅�O1���Y�=�7=�z��q����!�G��'ng���<��j쵿<Y�dqp�y��_�d��n�0fo�0����8t���篞�&�4���u�:h�ܚ�i
(�ٹ��0r��	��vB����I���PHLppp��!:سR=�W�����>���[�H��Qө<��T�D3�?'U�4�$ih��{2/޸�+�)P�AK:�~����0�#���j�Y~�*K�����ޕg
���X�oi?�VgU�:Ή�;��0����Ƒ�81�z�6op#7�6q�i��f59r�ஙA�Z7�l�q%h�:��������x~�r�>�@���3F0��{��O�l237�x��5U�VKYa�k�<;&���Ż��;y�A�R�=޳c�e �?^*�/}�ҎR�[7��cW:��#L�9����c7ӰF��M+\|V%��c�3���e�YU��Zܖͯ/p��8A4ex�dU�4ק�Z~M9Ƿ/c�\�-��I��0��G����$�D�q�o|hg/��҈���f�I|��{x��3���rjʆY3���.��s����M�Ҹ:70q�S��r��h�S��8W��-�^���6֩݋���4/���p�v�I҉���ݒ	ԭ+_ij�>��򼹧�����Q����௳��r��J�K�c�=�P)bnCvt�;��!f��r���v��0��kN��#������V�����Z�scd'�$I]$�G<�>��nG��7D�U��!E����݌�$)��$�'>�W���H�3��_�{J�p|l ţ�?��T�j�cy�d�����Ϗ�(�uzl]�zd��#���������XxxD2��K��@�P���ȼ8C1�q�|ϡ������h��~��#�;���n�{��4�R�b����B�iD�V�}]�Og���*��<7^s�gwFJ'�^8�9̫wl?��b�\�X�e�Cd9���9J�ɝҲ"�`�ֈ�|�ZG�K���h i���JR�D)�P�g�y�N5��/�4x(֨'���]�����sU|טg�w���h]�p���KN��#�Y�ZGG�>w��O��){�����'>%��#�_���J������Q�D�]���oV��#�㋶�E����]��qR��DțOSמ����m"N�F�=糎'ЧO����Ux�8,{��"�S�>2(������V��Y�T8�:��G�ے��i���B��ң��⏽���]Kۡ�� �iߢ��-6D�,�������.qYQ�*�葄*��^��(`d�ç��m�B�"&d��&pt�%vD�Nl�������F���,��0�Ƭ�b�qߋ�^. �y~廳^^#���E�!��y�����5=�ƽ�[�AI�1�l�-j'��#�:�O�ێ~�s|hx�������-W�:�+U�CI�1g�~١�D!IQ����h�{�M7��g^�N�����>BW�C`Ĥ-RI�7^M4o�],�ڬǾs0�Dx�K�T�>�a*FU��U�9�Z�1+(R�_��E}���E���˰���r��#��K]�w��vO����v�S\#yW��|8���V]ܕ󽚨>Iʢ)�7�ӳ,H2����to�-�G��ح{�=ۊB^l��^j����&HWJ7ElZQ�uv�L���%�����]��q��mn��m;l]�e�һ9���s뢓�;�ҙ����6b�W0v�Aݭ��k<�i��m����so�w*Ga(����ey��s�Nwg����d��H]�˄�n����cR5�d�Ny�[���w%���s.�j4�Q���<͐]�:l��;��t{5�!�Q�<�e�)��/="E�K��m�j�g�����>�D{m��nL�Wl��D�T�֘�٤{Vj����������4G��ȫ'T�H���}X+��ܤ(��LR���H��������݅��?"O0��|�<G6�"7Q4B8yՇ�c���aDO��9NCb��F����[�E��]�����"*������x��볶�>:~��`�/qؖ�ل�<Q��'��dV�	"O����C!z{<��h:I��`fXD���$����!	���~*�����7}�X`�e�h�Ogo���0�"�j���]����Uߍ��^@�Gi" n��]5=�'�{ٌk���~l���I,q�2hq���Y	�,����YӇ��Iq�{8D#K$�8w���B)<@ڒ[\<��wk���X���ăt��]H牉7
�NEb�|�����L��
�ƈ�D�a�ϵ�o���<s��W�hY}� ����8~�#����Q����Q�h�L��{����M�D�ʌ��;��]n�eu�s't�[�碸�^5�ReH�n9p9��T���2[?.�8��W�n�H��dE�Fj���>���$�B]H��z{��9铯<Sb��޲4�p0�����z��:�t:�dx�s?G ϡ`Q�T�ٿ���[:�o��r��g�� I��Pͫ��C���>nn��{rJ�e�-Jt��ق"���Ջ��S�0��'*�t:l.˭ܚ�/�Eʀ��[�e�q�iƕ���(�2�e�vm@��H��
Oߜ�&j�#�'O�Ea�ܷS�<4��ߡ>$��9�	LFc�@��(H� W)�d/~��|�<$h��B�	�;�ӱ�����B[��bT�~�EW`�!^��G�
}CL|���b������դ+y�3���6�E����(����=���|Q��ȡǈ��"���E5
"L�h�%�p�'y}�H�f�(!�q��*�OOm24�g������ZN$L��0��H,CO>��}�Q���>�:�������$�av!Uu}F�M"+��4	ӆ���D�(�&�ّo:	DRD�C�/Dy؈9"������ړ��M��]����W������s�Q�g&#�:ev8}r7~~�mC)I&;`aI:��� �GB��V{�z��Ն�'e!;~�7P���3�I��~��ie���aF�-�!�S�C���ֱ�܁F��H�Qk��F ��4�G��z=Sv-�������~�laIY̿f;�ir\�_2���^
�D�Hw"}#i[~�C���-����<Q���{AA�ʕ��i�cORQ�,�=U�>���Y&͍b��_:=�j=Q��蜻���t��t����佗��mE@|Π�^�m����r)eWv�9щ��N	Vt[�;�B��w�6)���h`�<HE}��Va�'8��]V~��;h1Č�F�t8A}g�Θ��q��'����X�*=��uc��EJ�hQ�<��(9�p�$�tn}'�f-�@�dJ낥*�2��+�-��f�N=#�w�cJƨ�,��n�8���zq���F�ۿ<7c��FL��U������7��"1KB��o���MD����4X��e,4a~V�6��r���>�V��D��kB ��q��Ψ�`k�����I2��������vN��a�bq$�i�!��=����I��G�Ş�	^Р�}fΟ��'�[���:T�$i�l����(�^~�0j��rox|�����d2I'>����;*8�^�^EX�|�Y䔦S��x"&;��%$@�x+��$������D�mb�6}��|����+a�&Ï{�Y�!�F�Lp���\�&����8���6r�迸�<B�"�ԏ{�ݎ?I˱�.rC>�a$��c�xp4�4W��O�s�n���q")!+;���P�:K(�V.'ƫ�����Q���N�qfvv���_Y�$��'y�vFsu��"!B,q7�ğo�(i<(��OY���ѹ�Vj�k,��yy[��[ӓ>�\0��{N�r��]A����y놊X������Ve��A�l,�L Պ�~���6�1�gm��R$�DX��C��mD���\���L F�"�*�OӐGF9�!byj��,����#�Z�U��@�z�P��4|t��s��gO�hH�[k1L=cY]+ᱧ�QC��r�9�<7��=v�b5�������6Ϲ�q��ƍu���R�m�������l��y�#����(3d$H4Q=u�E�u
8gT$��>�6�d=+3~��8�(os&�E�ڂ���"/����lt����٥ֈ6����;��h�u)�ԟ@)Np�&cZ�OV衧�9��}�t=��2(���Mt�&����8E߯Bj|�F�s6G�~kK.�`���G-R�f,}{�~�(I�g���ǙB�f��W�j�|���p�F��e|��r,Xi=�@���{��k�����A�B��=���P(��n�:������]� �BPv�E_�ߣ,�A	?h0h���Pvjz��$�͑쾸�GH�(Y<�`����������P&����~�ߎv��'#M�n}Ǎ��T��J�싲u"A��n>�T����^�m�(��$�Ezfk�A�^h���g�kbR|"����xa�8����Dʴ�&��D
�a����
�����E�R.Vr[+0f����,��X���-E�i��,���˟Yݷ@͗z(d.����B6(K޷X���>{tr���{R��W�-wi�M��̫��)h���S}wŇHVm�2�T!F�X�P;V��Z�M��֛(�������m�J��cջ�K8z��-����fH5�u	�hG�����B���Vً�<@1�}lS}]�k��5�[3�ۊ�L�	Z���X!�~OE�N�#�`���(���Km9J�L[:I�����	%����xp�E�CuL���r>R��;���

���M��iՏMq���əΦ�^b��ӯ3^@K�x!7���8&�*(�%r����v��GfZٲ��4t^Ǯ�le�uKh��9%u���&���dV&��������W�^�`U<d�R,n� ��5��XYw�uam�[���*`u}c+ ��>�W
�����Bl�RؓK��Q=y���[m�\�l��������T��BF7^.J����{��,蝭�>�0�)���R�4ݦ��]�{QQu�t$�����rF�Y��Q��]y�Af�oAB�r�t��7���h]ڽ��!ckò��9��8q��0 ���J5�_@.񹂕uIl���dǎl����8��G����n����r^��6>9w�?=ͼ�kr��D�k+��WI�Jv���z<˷��f��vZ�S,�ݿ�2��ԒH䉶�I�#
Y$�Aؐ�-��5�� ]c��)����=]��\^� Z�U����+ƌ�cNA�4��b8��Ji.�C����{(2�m���yS��y7kb�#l�zB�s���0�9yܱ>E�u�y��-Z��=vl�7柹ݟ��\n��m��)(�7]/s��������+�є�������\	����y�#9�.v��CBr�7l��<���ޝI���q�&㣪�&+�l�l7nɽ�nv��P����Y��4�j��7oar�0u�css='�c�s쁉��\�}�����e�x�;p�y��ּ`�(�:���q�����9;up���nz�����wX�V�Ύ�s�X�R�n��<���tI����Y�<�&�[�/nӗ���'ph�qurr���uK�Ɛ���:8״��v�-��ۇps��!�/m�ە�{���o7
ʧ��nVn�.��䜼>�x�a�컅[�u	�7i�]�m�&�\)��]En� ݝ�q�g�on���f3�9��;yۛ�W|���$���G�79lA�3��p`�`��t�M��mgqm;s�b���n��p���cs�CBao:ֵ/����{\�n'm�+]ǃ@������ݸ{�����#�	���n��p��[q�ڜt�$�k����X��8��v��kH�l�5�Y���K�t9<�ٸ���qy|rF݊uq�����SvwڶDy���:���u���ۋ��3Ձ0m���]vJ����S{��5���v����Gj�������[�6U�uF�q��0v�Af��\j�tٮ�
�n�כ�Nh��>N÷B㮀g�3F�5�X���N���痂��6��S7<�-��\�۴GS��s����R�:��#r����=Q�\F;S���v2�<��k���q]l�a�X0�8�4v6l��b���N�}���v�Mv�o[5lu��{<I��q�%�v0������ˬ:�lc���}a�����\=��`����]��f���7��%����v�6�� n;cs�l�6ԡ���+��֗�ѫ+���jٶ�i�tf7�z�x�xȝu�ɳ��Ѱ���ufѷ.�М�����v�K��v����$���-N���eQUG���u��6���Pv�z7AƓr�Z�:�c�8Q(s�g��I\en@_kp�4���Wm����@��6�kD�oEݷ\����8��i9:6��8�խ��.â)�;�1��6p'jT������88!�F��Ӹ��۠8�� J��p��3pԥZw=I�,/.�r�_63β���������@�'n�~w��G�(�{���C�1���9*�*Ϸ��xN�.{p���L��yA%�{"�����R'��#�P�!HP)�`i�Ϭ���G�l��m�jFNq[�*��S?8Tm�c���~Æ��ǯ��Vy|�}&0Æ��nzb���ctc��=�A�d.7�x"�N�E�\��C�������Gk=�B�f���I�~ȡ���6N䀹������<nG��h����!`�L�3~�Й	�Π��C�"��I�L@��8�iY��S��D+j�IDe�{��6�$����P���VI�,�E���E����'� �3��Sx)�����L��b?~�ϧ�B���,�,����k����8�~����Y�&ɍ��^��4�?g=?.��y�Ӻ���=@�8A��h��M��UH2��bx�}��?�TL�Bm+�x�le�V9�9��;�9:�&b��9��v��Sbۇb�a�g�߽���?x��:�7�1O�P�ga���E|e�"e26QY���9�_M��x21�I�M�0�5�>�di�n"5'�7�	l(�)aj��Y��R�&��������^��������,f�	~>�v;�ʁ��}XP�������gn�F]��2��s��i��Ԡ���J�a�OX���y�JO�ؽ��r{�"8T�<葵]�bb�˓�ߠ�衤�G��!���n1v�#�����AOORd;�����8#FG#��Ič��U@� ��ܖ0���`������W�5i��VԜ����=�:~�a�ť��Hy+���-C6}���i�g�x�W�([U�Uź�s:&U�=��<]1��.-W���q��3v<:P���C���Zl��ۦ{�=4�a�����584��駖bԺ��X��}_��l�B��K*��ڶ��qñ|��`�X��L��6w���>���/z�+^��ua,!�	����1L�8�Dp��=���+�Ǡ�0�nfl_X!� r�Ϩ���ݏX��,�d��F�m�n��t�nW.�x�̏��ڳs����wF��W�E�l4ZG��sҾ�M��Q���ْ���^k�����(YJM�r���2�^��.��*qqt� �0�M�cm���qг�L�yݎH��lH����
�Y�9"C��_������IU(��v�qD�(i�p�RdY]�#�1lPt�"(�Dj�"���vF�kս���!E��H8�M>}!.�M�(a�U�44����|da��Q��
��&!�����̇�.ה����T\ڝ]ӯ�Z��ƅ��Bh�G�_^��p���L���|v"��Ք��:�W�e��h�#��w,=�c�����EG��ae��G��_K�^�~4�$��
��|\iA#�.���Zp�1W�nT�f_���O���������(�_,H��ՙ:B�*��-5N�{��'͟H�j>wu��g_\5{ԅ�͹�$BҾZ� =b�8�ET�ʜ��V���w�5��	�[�2�@|#.���=w�V5m#�:~�5϶�d�`�!�<_K��c�"F��e�D_{\fC� �߭K)A��4/ZV[N�l�͞��mt��[��=�E��wna-v�=�,ۉ�lv]�*����K���Z�߽�C�4YS F��^���6����AZ��W�VO���/�p��A%�$��H���W�i����O���+>G\�iqrp�Ӗ����ZG%N�>L��p��PZ��F��U��]�`ᣄ��C����sVwP�������<j}߯O�R�kED�X����� ��7�C�6��_a8�ޛ�v`��0X]�^=Dd����h�����I�p$����"���C5y~�~��.��PB�J9j��oM^���]	�[��W��gN}e���x�(�s׹7d�����2Ȑ{�$���
�H�}}#�_�~�a�̴�e]�*��o��2�7��ޔw�\�9_�ÂT��wge��`gT��imJ������ǮȬ��Y�mU��fX���3�R��Ƽq����5D�X��>�1�.!����n,�N�ԥ��$R^�}����Rq!|��,*�1�y���M�)��1
H¥ŔϮ�8D�?Y�n��KP$XA��$FTW��}�N/T����4����9(�_�w�,���^\�Fx.'66;:�wg���d�flT��r7���19<4�3�t�l�1��ۇ>�Z��!gH����V���0l���܎�{�Y����p�'���w_�cW�=�ԍ���Ql��9)�_iq��W�s�wE;�v=�Cy"m
&��i�ٞ����G�^,�L�=��f�ƟJ@�E�>�5i���`ʤ�}�����o�V��*-d%i:���\>�C�簦 ���� �_��a��K���;��?,AｎlcH��������b���4)A#R6�(����&"q����|$��ĝ�ؠ;����+�����/�����i�v�n:��<p�t����Vkԋb�~͈J��Th�o�mh�]��~>�)~��Y$0�\CF�U�_���8��#0�8W�����7U��u�CQ��4�h�^�z_׈+H�(��$���_�X~�a�+vb�
�A��1�K�pfϾ˼�[w�ht�i�a3a�[�R�a��C8b��e�9��Ҙ�nxj���d�}�Y�^��6�� �e�j��RM�yn\�d�h�`y%H"ݴ�㋎�/9�#S�C�7\M��Gkn-��x�+��{n�n��C���&1�e�ۙ��7m�N�=.^1����i���J�dN1r���n��)�ݱ������_$�v]�'k��3�+��<��xg.��Sl�ي�`GA��]�UF.�VnGp�g���8��kss����8�,%y�!�qڮ:ݑԍ���1���N��m���^��}�}�I��.�NN�gY�7f�9x-�.v��z*��<]��[%�c�����H���d{�F�o���:x�8a=�>�̋�F D�-q�$Yu~�Vwr�1���ǋ a��8��4x�N(�1�4C9ފ���^r��B��4� �4��-\ɞ�zv�-.�\�?7���u�7zv+o@�d�őGr�D���^��t��D�on����X���^�o�� ������#�R��rBً��5�~�Z�G+��`��l�=P�p�X�y�j��Sy�d�٩���D6E����j$�Т!�F�sүP�8F�J%f`�<d'ϠP�M����|l�WTO��O��%ey�zN|��{JR!����y�^�M��$Yհ1{�5�HX�
�H⁽��#̺���Auw�c���)�#������D�҉)�G�F<���;���vD����Ez��-s8����M}]�~8Qya^{�8��å�b���_2&���mϛo.���7���z�S��Y�}u���5��۞���i{s�zB�\L\�#��z���v5�m���[ō�~�I��'�U���F�9k�,HQDϟ�P<{4t�O/.QS��yu��(n�g�����:~�>�4�$��B)9�I���r~��; �[u�^��9	jeiF�/v�E��+K�r�\��F�ʟ�n��.��8�Ի|f��ś���*���JpՊҮ�h7|�c6�܊v�d�cCq؃1U�Hb�b���2C2|Ͻ���@��n)(��1[�aT����ǹ��=`���W����1�Z�o�|~���<KV3���`�	E��)@�-�����zE�5/�󿬉?F��V���ņ~�w~�����hL����|r[�����`u�|�����VOR"���x�h_��O�)!�����4,���D���^�c}�zܗ�ęUΚ<��-�ϥ/[�u��6l�N��"�h�x�'Х�I/b��e0��˛� 釱$�x<F��~-Td*�D���/5�Z�Mն./��9d�;k��4�U@v�DxZ;^�����5�|�cެ8��X�#������ä���}�Ͻ�m>��6��>mE7b��:�ۡ$c�5`ʰ�$�����q
�S�ɻg��M��L����sq����R�,�/��
ı#�)�U(�"��诟!ؾ�,�~>�ą�U������0�<D^{���Nv��(:WMe�;�8�,8!�D�8�3�:�7(*H�!N+���$�Y���n&|u������ʭx<ԑg�3Dv��V��W̌�Z������<F�{��zN�xڽhc�[H�5�e(@dL�16,�H�T���Da�}�(sOz���a�^���!����8~����[�}5L\��2\��q՚syP]9�;��rs�^_��\wk��EkK�Γ�"%r���Hn+��]��O��"�%�^��D�؄4�:Ei�h���G�Z�O	0��e���ˁ �S%�0A*�����R#�d-�{��f���E�{���9�+�n�dg�48�g��{��)*��'{�Vz~��#���E�xW����j2�9%:ZT`#:�Fu{)м$V
p���Q����:���݌!�B�+~���^�#2�24��������e(���9"LK���v� 2�]k�c�K�v�8�۪:�{ �KCj�q;m�oT���^&�i�/3�l�w�߽���x�M!�ۏџ2(�s��o(Dj^���vp�aCү��zP���?�k���-X��{~�ksK:!ָ��1�;�8|�N.@�%89���E��0���UGa�<a�3���α�����A�����C�@�	�0�'���B�oih�}u�;�b}��}�<��,ߑ&����8޶�f2�p�N��) Α������"������n(q�$��وs�^�tzy}Ѓgo����!Y���p�m���:~��M+��D�+�ڡY�l�l����ͮ��OC���||"�(��qf���S��Bh#�Y��3��C���<��̻�vJ��3,��CI�oWZ����u��1 r���{�e��ز��[v>�w�C �&�����0��}��\�-Z��0�}�{�����ߠcGӉV�N���Cu��e��j����c��n�
$���Q<NT�#��:=\hUll�˞?A��H�J�b�!b�9~b�U��7HC胸,���>Z���g�F�ѧ�<�l��<=X��� *�;l�m'/PQ�ܻPl��uDMZӌ�e�;-��^���\��D5�`��P�䄑z�������}���JuKC����z�#{DH��yw�D{�<A�s�E[�lB�E�D{���rD�-�e7��a�!dk�/{>�O��7뉽5�
$��ƛ#%��4��?Y���}�:XF�g���h��_Z�{�~��l�<BMu�g�?"����l�\��:l�5,����t9�DP�_#P#���B�[�Gr��UE���!�ݦ���,Ӽ������틬��O�6Wdq��	������3�3"�?;H�y���pJcF0��w迴�G�P���~W����e�u�A�ʿ;p�?sR0���3�X4��ؠ�ѧc�H��O�;����%W檟Z�V��0揺.��5��� �B9�tANՑP� t�{�@�3�=n�y
!�.�<> ˼1�n��#L6	�_�����'0� �[L埆�w���X����A8��P�P�*Όo��|��ȹ��H
���Zժ߳;���&���B�',z�������4�s��k��|���р�Irk��M/)���8V[c�N���<�z�э�y!1�s�1���_���}0��f�<�<qq�Lu[i��k�m�T���kZ�]�n-����M���a��p�7k%<b:z6wm#�mۙ�M��0��ɭml�r���%�nؙ�+э��h(\�1��\;v�`�V킊M2��#��,v�N#��F�����',vb�l�9f��\�8�R��܎:���Wl�"���l1��ͭٺ�5v9�f۳t�k{h��@�R��#���ƒ��~�d�;��up���4О�{&:��h��qLH��c2�R:��"YY��5-s_Y��Ȼh!�e�!4�q�����s�+��Ԏk��o
���=ho�9]W�9�3��Z�=��Fȳ"mGlG�1B�e5�}��Bs��VF�|�������3rg>�?rc�w|�Eem�e����CH���9Yd�`g�B��ܲ��HY���١�4�eVA=��Ӝ?p��=rW��#��8��OW�W�5}����"w3����;m��f��x����=��mD秙��cq�gW�a@���'S���}����Z��z�G����x�"�cH�RҰ�g�ÈewY'�/C��e��+
$�W��j8�2ʐ�1&��ђyo!�pm��o�y)"�F����p�{E�!���<�F>�fE�j �Z�����G�ҏܾ���"�=��+,��x���<������<`/7k�gI���J{o%�1��Z�↝���g�nBj�4�N�L����?<���4��,��dP�4��[H�#�}|+�j���~o�f��y��;*�B�.�RX&f<Gg�����#�o�Yw{�bh>r�-�� �L̖t�y�qY���fJ2(Tοr�5+DTbE�5���u8���Q���}�d��j�����4�6�--QU����k2nd1��/�m1Mvۄ�{��c$O�k�a�Z���=u�;�"��E�!߯b�F��[��}�+/G���0fD�l�* ��k��$��u?{��47�Ri�y}e�.�u�"
:H�5~�i�\8U��֡��gHX�C��<��Ԉ;�n%��H���}`����X��S��5λ#�]uߔڪ��s�O�E���'�B��C�Ϣ�儓H�5}i1�B��G-<5��sA���z��5���`�DC�n�_�m��h�	A7�h��"�<3����ӄajD�)К��E���W��6Q�@ٲ��E`'W��VG��"������GKݱ�ΰ%����d�J2?R����&�rzwa{3Λ�nۏk#֮�ƍ�[�`��Ё6`l��ф?ZN�$�D����?w��L!"��=�K4;ǰo�Ζ-|����uݕ~ϽyM����j�ʭ�Y�Ry:Q�O5���e% h(�����R���>>�0LX���w+D5�p@j��k�ưUЀQ$;�z({<���(�Q�t{���FT��9[b�����?g��Q����p�8��DLI�M�w��}z��֑Q6��p�Ń��@��;6���g.�c������ԣ9=�&R�grw�X�j�b�a�����*��{>�"�|�)�"*Z���ќӷ�9|)�e�3d�����z�"{�8��5���ق�c�u��� -d�쌜f�Gl�2��w{ogTW:��A�kt����n��oJ<�_H���QN�֫kg*n�9a\zɩ}7�:����M�I��7�JaY}Rv��9ѭ}8��N��6T=�;ݺ�V*�$�,QvT�]^Ѯ����`�;]�9Y{Ug�^]��%�	G�h�DV���Yi��n�R��C�d���=�$�k�\�h��ٹ�u=��j�`|��wl�:��b��FkEm�9N��'-�IP�9�&jI��87 �:.Ԕ.���kb��`��^�)\OVe:ʾٸ���p���SN
� ��v�(u�S��l���~��5gws6������3�9�$�*�ץ���y�9��e��dC�ڒ{�R;# ��nn�6*ܲ9�!Jb�U�.܃;�d�:]�u�6q�;���+;Xt<Y�.n���r��x�A;Ҹ�"���p}�;�%�٧��Z�(�wo���7sx"V��v�v���Þ:4(��cc�ou	�1���J>=�jt�z~�¸�5���-������GR�����n�m��Von��^[����+��Թ����Crgڝ=٤Pu�a5i�{�����ZU�ߦ+�O�S�ŝ�=B�š���FV��G�Y�/��b�I2��w5X��(�!�_ő�^��p�H6�tRh�}�s�aF�s�S�[���9�+��Ǽ��#Kμ��đ'!���_�v����4�Aq?!�������u�oR�=�Y��T����ǌb�#���R�%�BjI�#(+#"����珲�:R*�$�A���Zɣ��f΋W���o
$�F/��J��2HѨEO�N��-?c顨W���)������!�qG;U������
����Z���4n�n:��b��ɇ�wA�m�3+@�!�H{�{�,�,���T4�lI~��eʯ���,�$�Q���
�j?{L���^�1hU)hg=�����>�&?��kܟ�Q8�jQ�E<r�E����%dk�tԑ�ɱ��Ř�|IR"��A�r2�f��E
C�,*3���CnpM!�j���l���t���Ӂ��m�8����a}!85������r��sZ�a���Z]r�����Ί�:A4E��\��T�'}�>0�A�5x,/P���!��~��]�X�� ��S�Ƴ��������Ĝt4�a��Ͻܺ�a�\}�o�J$�gH�ȯt��}Fkc������CIiI����*��� �y[�;��\�n�s��9-��8���<�xr��u�o-n��k�㲩j�Z��L���|F,�g)��lP���a���o��>�
 �$F����a�f{�	�=5�4�8��W�3L�m�^��F�$#����윰��@�!r�=��D�:Q�Lu,��q޼����Q��hD -׆^��Lt�rA����65+	,s&���F��_�l��c��$��My�ٳ�\�����D��@�d�����/�K"���<�l�
#d|�Da$1�-�#t�tm���Z'��<�����H�%8[��T�7}�3��~�z�+	ծ����U�0p$gY��FI~�\#�ekd2��{9j��8ZD�B#�>�_n�q����G��D����0���̐D�E�(a�f�'���DX�z�/H�(���h�V�A��^�=�OG�Vx�=TD��=��E!�,rx�m�:v�/�k��x�\VPh��l��[��c\e@\��}�����_��p�7�ܶ�>H��"4 ����_��h�0��\r��P�~�A�!g6�36ڜu�P>����icq��p8(�����+n��UZ2׵�EE5�u!o'��2~�tQ��۟H�V{�ߟ���Y�
����/��f��ȣD2;�C��TȘ�\��u*�����X���/�V�bs��xwf�b�j�So\�d%W�\�GZ��D�5�g�=0fܩ�n��8��ő�[|��N]�7DB�ѩ]-�����;�iwA��Ʋu�t�wg�Rl9F�9^2�*m���7V����Yd�X��a��l#�הዮ���듞q�`���ѣ�.�6�OV�v�SɫY�}�lS��m��ְ��ͤ�6�j�F�i���]w)��]����D��G�]�マwb6�6��wX݆��lx�g��]�[�Ne�@0������,R�sOX��v�ŜT�M�ݙ�:�l�I��j۲.�cZS.�FvF��;�9���g��,�7\r�~dp���_�<H����
��DY�����_o(��u�����Z��}+�)�_���SD�l��vE#���fN��A��^�� ��BU	-���O�Zl��;�ݦ��K[O�OM=�ĕ�`2u�<T6z>��j�(�{���ei��_:~�L��Q�K��z���d~�����A$�RU]��F#�2Db~~5�8�Fj�0�/{�j���o�a�t`�ه ��<`�9�r(W���p�!��q�}�oN(�At�����o����#2D�E����Nj<j�����}�7#���~���O�����_
åp������b�,�U#����rq鵝��oU~�hx	�]|h�x����S�I)_i�� ��B�^�{��$�!��}����O\����E�i��2E�!�K4���a7ԋ5=�J�DXУ�"��{�Qw���m3�HQ�.��q;�>l�״��V�rM�̇@��'��=�A,&J��˒ӞL+�����<`繏�ΓOc?-P���b�f��g��ݛZkgܨg<�<���ݩsJ��(�[��z�e{DUTp�}`�q~1>(�8k�:�#�@��nӥH����c�*n�׷&�y��b���T��˥Qu���sTo�Z�9�v�ne��P7�
|��R�a^�U�B����Hxt���S뒷�3��7��2�2�"��.��*9�A�ZE纯�#=���?A�߰a�N߸���z_�a�R���-�@q�AD��?B���h|v�0��Aﶢ����k+���	fkv����zlг�Id�"����5'Hf��$VD���'l��)�u�N:��� �|j�?*�A�D���G��}"u^5�t�G�����(l���=�׾	;�z���g�]��"x��;%��������'jGb�#�m����%�f���;K�n(����6�+l՚��uY�N$I{�ȱZ��6��0��}��w%#�!dXG��  ����<���m�I�������-�hiQճ�]\����غ(�����S6�L$���?��~�J��?���x( �������b���M�,���m�]����@�����,��E�vῴ�ڈ"	������~D��i%��S���<������to��\gv�0�#Z�6�$���c��q�B_\]�''=1A�"��l��ߖ����]�[��t�(���s��,nJ��il���u�ɷ�{ ^���<�TP��$���7ύ�Z�$`�՜�Y�Nь�=����T��+��Kۢ�=����'�l=0oY�����ӕ�p4�;8���9'Ş����>#�CR�T�ffȢ+���^��H��Rt�x|q�Dt�eP��Z��??7rc^g��"ي�s��+��F�wuW�m+4F�8Y�_�v:$�G�"F�:��Z��|G�̜��{F�/_۸�(�'�ǯ5S���^����!ISN�jvןq�T~���\�U�7g�D�>�A�t�á9+]���W�U���;�#H�:d��p����8��qVo�D�<B����a�]��=Io,@��C~g���D�Lt&����8�7O��[bcj�7hk���<��Gcn�GFJ���b�Mq����/o�Pe�J��h*P��=��'hW�
��G�{����[.vv�+Skl�E�q����#��}Q@�G����,uBX7*�RJkO�k�=5���4�P���c�:�G�g ��K5��W��8��F��o�E����x���NJ_�٪Ӹ�Y�'�⣜/*��m}�c�^�H�l�mǃ���� ��p`>|hX,�?l�6}�O�ύ��cT�8�~�M�zs��{��.
�[�����E44�U�J$������1�"h�gl߽�&�,���"�E�G>#G	�oz=��:~�:�P�g�����$�J{'���P�. �!�KB��=�W���@��=ݖ�.���Q�c�X3�hڗM\��[͕o:ki'O]��c����&��\f�	�j˽s�x�oy��U�φ�5_�kO�~������:[",2W���O'����:�Tf�DBO�P���?Ĳ`Q�U��yJ�%�ڀ���
�fH���ƽ���$��
H����n�R۸<h�<i�����ɉ{u�ⲽz۳;]���gv��/B�g��n��Fp݅��:�ټ9���3���:�Xc��t�B�!S?I=�I��u=����?~4OF6��/9�Y�x�%�ΐg�E~��`�g}�C����&?�dV nK%�^6�5g��ue�_�}�d�dC��G����ͥ�P�������h�u��C�"իMZ����Y�J>�]����=�H^�g�]�-��@�D	8s�i�TY�C��B�<�A�"y
�A����y�4Q�Ճ�T+dYU�#٬P�^#q
�HK%;�U��9�@�9�s������|c�JRյ��CliM����L�����&q�V4�Ö��a�����P=H6��&C��tqW��)p�E�-Mk>h�~��c'���^#N�2͢����m��RGJ�M�#��eOj��V���elD�%6c��J_w�V�<����h�CN$7ֽb��+�ހ��p����*?D]�(��*?֨_���\��P�/�.��V)��6k�*�+:��"�����̷̭N��;�x%A���G*o%#%̓�]�A����TQQ�;yu�>ƞhSq��Cn�s������۱��;@�������LW�֟K��s�dېCu��n�8x�l��;�W'g�����T��t�i��`�l��^[=\�u�rkk�H<g8)��{j*��'�*ˎ����w	���n��n�b�fte��0�i�H��p�
��i�\9�pi9��ӧn��'�8�j:n��:Dy=3��V�4��1�M`�Cc\�Hn�����-L5��B� �Ɯ�߉��9<��=���ӆA']�/>�n��0>��?mȁ�����p~���}K�|��rF�?����ҫY'Uq�b<���%���V,�@����u�~x(g�S:�<5U�_i�}/U}���(�R��{������i�3�H�m��؃�g�>}���A��1�'i�x�ؐ$�>p�4GOH�$sջ��Ӏل(YT�U{�*�l�Y���\9��dS��|���D�O�����}�`��Q��Yd��r''���*�#
���\�ʱ�w���f$b=*C���P�i�ȳ���˴,�~��C����^t��]^��~�,�/�*��jM��<�����{��FC�D�J@SpW	����,��ק��F��k{�o�1��ֈ�N��c���Խ���7�G�l����/��gsΊ\#L�0�"�/,�H�W5_}�@��>�-M�J�"H�EG\�gk����`�:Q�k�\�Q��ٻYܵR9` �d��^������9����"�?CD�_O��8������B����s^�aQu~E�3/W�}h!�H�ӗ�ZFj���>��"~�_>H�3�'��)�������_�W��mN e��[F�X�c�1�%�)���p�����]<�<��E��&�KJ��(�����13geNR�o��q)��6��XA�͊���ay���ʖF`����9f�G�^��q 	�>�����D!B��l-D�L���mz��3�J�`�}|�����'��a�T�Ն�(�l��7[�Hx����.�@D�\�䈂��T�ƙ5~����+���XGT��BI1cNU �u6p_!�����i�U$����?_�"�i4l�p����cőGH�5n�/>���V��O�	]�p�t��4\%�����5��3k���P|�4��b�8� �о��}\��r�N�s��Z��9�o$Eb��"�|�#� 28񣣼��̃�ՠ�`���y��
���,&YP�bi��ۋj��z9��F.��5��ݎ�V|��]E'#����TB*	%��?�F߉���g�� ��\Ly.��V���K����q��5�H#^Cu
1���Vqk�{̂�!494�^����%��,��Zo�9�F��\�6�F?g�<Z�Vo�����z��AQ�gW�}ooi�D9t���{Y��EJc���h{=|uQ_�J��y��Mϡ�)��u�-�y�@A󲭭�[{u����V��l�(���	�����awz�#L<����[�D�b�ng*�ҷ\9&ǳr�i��Vg0=�t��� Z}��Mf�����t��`]���U�l��]z�*\|l���&!r�e}��ۥ��="��t�M���$b%$��;���^�*���~��$����e�$V��{�衆�6���9#�F�G�W�@�Ry#|"�j�0�|Ȏ{Ƣ�dN�"�5�A�ǢL�Ҍ�N8(i��FH��<��=
���B2{=p�Ic�Y�<���:\}e?^L}��:� r~�<+#��{&���{�@e��NS�c�����ͦK�@�A��d$kv-۶:Gq�6�W5��wL���
+�t֬�]mr�jm�XRGߴ�R���q�ᳩlh�(�N�����C���f-"9��
��D}����Dj�D�N�W�g l/��?:��Z�%'�(�REcة�qB͔{���(����F&�3��GEz(g/��?V �/�B��k�20��ƽ+�$	=�����WC�~�桊 �
�+ez�Hv�v��3��C�fH����{��Wdw:i�d`��~���$�y"b�6�8�C_JC<���٭�����!�y�7��UcqRIlŋ����]>�x���8����۪�G�Qdzw�4;�Ɠ�zl�t����z�cP���v����A/��v�tA�e��J���oi;Ju��O$��]�4uy1w&�a�uj}y���aB�۠��黲GK4�v����3��`x�#Ѷ���g��ZKcRR�_w�������䏼�U��4���u
0U����3y���lՐ�&H)$h���ɻ���y�$I�=���F�@#R�l��k�	ʵJӷ�6~�ŨX,�>,��<νѨ�&z�C�ur�B�%�҉��l����$	8r#x�f��"O�� �F���g$-�m�ˉ���\~�Az�ج{������gd���0��j��_L��K!�܎
 �2	&C�@d��F��7iG��d�|�㱆�%=T�d�� u(Ȃ�k�iC�Ahaz�W�M3#�|�ӂ�}�dU���Z�� �_z���y'Ã4Y�FϬ�PE���U��mu�Po��5�ǝ�Z8��)XA2`�{}���27�������v��$ׂ�Cg��g��ҷ �^��?��-g�A�#t�CQ�B�>e���n'	�@����(�ڗ�W7�΂��d�#A�mi~�񯣉A)�20�5���C�dC&�f=RU{��t���#�{�����?��qUT��#*���,�6�V4'0=��_q�貉1n$�պ�`���/����o2����X�P�$"���(���5t���(�H�6D�>F���:d�����Jf�bY{9t��re�f�y�(�cR셤[��p9Jp�tY����ҡ��:�D�np���Sm����NKՐn��P�+k@�O�R�(���vlY�aqF>�rH5M�5Yxb�8��9�����:�5�Wr�f��w���=<ضr+�[�9����q7b��ԙz켫��jbъh\z���ڝ*vwE.S��g�vI��l�p�3{�wS�E:��L�|3��-�Ac�	[%�Ô*,Sv�Z֖��O_Y�5���_$�2���7g,��-�f���h{wq�J��7���jA]���2q󕥋�p��2n'�1�C�^�&|v��:z�Y��h����u�Ԓ�f_h�\m��V���'	����jO��/e�=�S�Ul9/�c]�F���vD�S��fC�wVb�J�]���|w�z��/O����rƷU��Ȇ�X�7\o\|�oOs�Q{Q[���d�{�]<�1n����c�oSvU�tk�}�R�'��.�{�`�}��2gړ�"���|�^;W�T9��S>�E)V��:��
���{�Z-�\��uُ0�}�U0͚�ٶ�"�"���=d���*Թ�q�)��})7[Gtp�J������;~�4�m\ޏ5fJ��F������h��s_V-��'6���'V�ZՎD��w��m�޹W���ӂi����J�vN�G_޼�{e���i�ӷ�ǘ�OK4&v��V.J�
�F+�z۫�����5&��8�?`��yZ�:�F�j�MM*ʨ�ڛ������때t)g���D�Z�\�Ê��%�-��6�5++�
i*R��V��kK��Y\�.F�k8�s���Qj���tl��v�#��^��8v9����=
v�0���<�n�`����ێ�m�\���K�cǌv���<,3����y�sݞ�u�vܻ����k�d׳ͽ9��ek׎x������ϗ�mv��y�6�P�M�k�]���L%�ɶ���j���dq��)����������ns�Ǚ�=���'f��zwd��Ʋ��X��jn;-�F�g�M����i�&Yf�۪x�2t�v�(ݛv{�q4��4Gbf��=c�����pg�M]=��z�Ź�.]l���m�1�[��y7k9��#��l��kԹQw:L9.Y�R��:�zꠞw]@�:��_>A &@{>0�n��zێ5����8:����ų�0����Ŷͭ�v�v��ۋcY��#и��F�<�;3�{p�2d��&1Yz�U�^݁�wK:Ѳ��ݻv���F���j�i�u�8:״�f�]�C��6��vyŭb3�3p]�ˎԘ�<�n�/A���y�;.Р�ɚ�M�E=<j�]�q�\+@�`��H5D��y��g��.��9x9st�N�&G[)-�;�^�r��A���nՒ;�V�4�N�^ї̺��Up覓0�6���%��9-��1δ&��9���G<��f�wWU�d!�;6����ݨ��lcl�����J�;9�/6��-grF"��]u����<S׬Y�]]k�,�;=kv���cG5)�nzW��kr�v���D��ۻp�<8�>�������A'k���\�y���&3۩'vǛ�i�tt�A؈bz��*�[v]�OV��N��Xk�Wqmσ%�¶�7��7�m���ڷ0��콸�Ny�I۝���i�t���1<۶�k����=�qr;m);S�n�P허0:���]��Y��]�ؑkR�;Hpg]�\��Q��n��z�v�ɝ��6�݆I��it����z;�jdj�9�v����@�¨������ݽoc=��f�4��;77H��p�n�y�)Αy7:�w�^�n��u�拸ꝥL9�`�;a����g���c��mK�a�m�/]%�M�=VH4��ͦ��sU��G9�n:mu���q�AV����l�3���힨��Go9t�l\
��΢�G�׵`�u��͝�vz��n]g��c���)����u�m�8��=���h�h^����8���pPb�gUq��#�h�qI��F��v��cG8�Y�t]�6`�k�1w�z��T�uqf��ފ/��دOb�O�#��ȻV1#�9|5�4�~�+���dXO�1HpJ��T3C-��E�W�}�y�N�H�x�sJ��6����x���>�D�	7��p��+J6u�0��V���iڕ���n*�hx��x�k���\��h��W��'�ɏ�n���<�n,q$e��G�E��ن��BHlc����w�̡�`^;��֣K;H2<x��ۚ�H�Eڂ(Ø8��M��"v�8�����]h��u�S�����C�q���'�H�&��}�(j��H���@����c�(�@���)y��zbj;�����H���ڄ�d{O��E�bH�!�4zh���X��{=�v4�.|QC6}=3�rrP��E�$Y����&�g�.Aq"��\�.j�ha�Y�����Do�(�H�(�����l����ܼYx��:{f�qY�tYƹכJm�[��9�WѺ��热�G�Q0�>��ȡN�ڲ��LmNt��%�1�Nc��2��$;����Q�43��"�t�����Y'�W��Fp�W&��U���/���X9DYoVuW�i�O����vN%u�}윱$����^9WOj��[�75�2���X�����h��+��9g6�X�7vn�#��v�[�#@��x<0�~9>����g�laGI"�j����P�1��$��w��ZF�2��~���ս#O�f�������7#�Q��x��D'z<�+�=�i"8�5hS��E�����ͫ�&��4\�2n��_v#��k�g�L����O�l�w���5��ґ1�G���φؓ�zt�,��bk|+K!dq��jOoʇ��HZ]*M���1W�s�����rԚ�zv����k�a�R���U��/��e3#)�jH����h���>�<��ĳ[��L*o�=�����48�Y�H��K�ؠ�Ԣ4�E$L��V�Y��-��P\���G��sa{[��ȑ��^&�#��Ɗ�T��n}�j|��X�&T��͝;�h6W��W��Mj���Kl����*����qL�<�	ԷS"G�{��f1_B�Yd�D�R}o==Uֹй�{��u�^�!��*��#;�CG�1	�ہXPC$	8r�gxGHgH�ظ��T��<��&�-r�Z3~W�c��h���򼪘��A
��2�ק�����g��᝛�{\/tp�dK�~�} e��C�
0x�: I�w���9��!}W?i�X��K�`��������S1{UCR��{�b֋�x��Tuz0����s��E��f�erڸsn?�l��L�$�v���zi�~�s�E�}ax�p���N}�ܾf-iw=���V;eU�[}bo�8��[9�)�V	��*�<B���z�\�{*+�}f��,�ǦL0�HdBb2u#E{�>��8���%ۜ~4�:�v�~��Y��J�e���W�qAM+1숙��3�Rh�?g)�P�@��	U�;��5]��Pt��F���w
m2-�	��E��U0�*2>�0���_6MK�Û����G-5B���v9���b��w�+]�Ă�`�=t[����d�LA*�q�A�D�ZCH�����_n�I����b���Ey}F�m}�qGu�����w��an�a�ګ�l�W��~@�y�3�y���fB"b8��P��p�py#�y1X(s���W1�)�!�BQ���VD��pύ�]�:�j1��;�sE}�EZ�wa�CҒ�����c�9`�QjGb�#�.D��aD*�{��a�Y������¬�ޟ����f6��%1g�|�O<�,�4�C�6�q��*�^��E���E{Ԣ1di&Bn+�K�6t���9��>�f�|��<s�θ�?Q9|�t��s��_<p(��T\���Xx� }�|��f����զ�y��P���o���Y�Z���Y����]�&�0.#��*�݋[{Οv�Qѷɢ	�K��T�/w��^����ä�:_$�I|AcQ�Ia��N�tȉ�g�)�{x�Y�Cw�[��w컸�S��U��ῴ1׋Ċ��U�k�R�BRZ�r>~�ջ��0w�l#�h�s�{��[f�����6�g!�7g�cx�z��h��<ju�|kh��-��}�䭑GI�����-HRDG��.���P�Zx�Cê>Ӈ���B��/��mq�L�}���ν������C�$�o�����pE����;��Ϣc���x�mO�ҏ���+�Iw﬿�em{J_G�:d��x�ΆA �h#�~B�٢�<hީ<Q������^��ҙ[ב��G��5��<}��o��[A0���ӵ���;��Ѡ˔��?Y�Ȥߢ��}2OUu_;w�D0G8>�XK_+�#�a��U��3��j^V~S~Dz4�JTnCqPÅF�N�<4�*��E}��2�� Y${�(g$E��΀�ߕhY�A�&{O��}�c��\t���d���)���!0BfD�1(���"���BȄ��}���1΁G
������Y�򿵭9hF��qi	v���5��F�=��5�x���E����wOr�#��"�5z�j`-5a���R�����l)�:���˪}�E��PN��Xq��ɋ�P;�<�B�^T9֒ȭ)ۙ�eڒ�A��1t��f��A��L���m�ڭ���t�ø&�����ɻtФb(��R�:�Ol[�lǕm��r�	����OO��qqq�rG�����.m��Q.��Op#uݭ�����.�u�������[S��ʻ�ɍxϫ��鶈�G�Sj-����u�ݳ�����N۴mk�7@:g��;M�Gڳ><��& �Aq�㭝��wOF�IM9^��'Mq�iZvy
�N�EHZ�����:O"M|�сk��?H�Q#O�TNc�8�F�$�؁W�tP�4HY�:sϨ�> �:6>�f�T2��8G@�/�(Jb6�m�Sr��t���eטD^��*�H�}�%��ؿj>`���Ro}�b�^�DzS��S`�{��_Ki�S�2\��W��S�iBC��Ř:Q����D$�����>"��W��V��3�6�?>B��ゆ�e�>��Y;�o���'�牻zE����Ͼ�viv>S�.��"�l6�����=����־������F��ԗ��*�o<�a�yq}r������]D�B��9J�		��V����!������L8�-�T-�(a�`�
&�!b��}�w"�a�ʞ<tv��i��^��A��y Y���߻M
W��9M#F�$O�ő����;�6��u�{�4*�<�e��,�ӳۑ���苎���[Z^Zv���7���Y��C	r#r8Z�{�4�l�B��Y��F8��h�$��,�������V,�B5#%�6fof�S�`���w���MO�M�{׵����(#ĝ"	�X�e���
[�k~}�omu���i�0��u�<�W6#�d�*Pdеd��3n�e��z�V1�:��c��G����q(*�}�����c�p����<�����W��-k%p��q�~��=n��l��di�,�=9�7{*!MS����^3�fx�^���X1����"q�⿺{���� �%��fz���.<�&}�$+������C���Ϩ��H&򯠲iU):�ܨG�>�����#ۛ���D�q���7��iL�RQ&g,�!����
��7��W�4�(���Z����Ea�V��Œt���׏���4�!�o��r��	�n���-<^�2U�,����%�d��Jgx*��kO����:Т)tQ&OQ�'A>�P�5X�A	:��2��������� V��Y�K��U�h�G�Z+�C����]��~�Y�aHc*��8�*+<��w���9��iG=X�5�����gt*'�	��NzE��D�{�>�x��c�Y�BU5�7���#��FR�q�����fOM��(�}$a�����m�������i���o��Ƣ��3"�,p��9�q�qsc&�G�禙֣t�auXdu/�-�Q��ڡ��ָFD��C��>�jF�\!�ߝq��r�?{�F�H���*����]��R0�Te�2AxO�FE�}�����t}����#�~�q�Q{����f,W���}��+)�|����H�W�<�&^el�sjPw�;��P��<μ�;��l�t�Á_�]�a��-L��bUJ�|'A�u��뭸ٯOR6i���9OH�w=)����=��!s(y��%ue
q_�5g�|�.�!���Is��C|�Ԝ"O�|jr_�Ѳ�i��0x�Q �7�8��p#�'z���5��ސ�{�n���[N�lƇ|���I,u8��T/PF/R"��{=4�C�]�����Mǽ��8�����5}D�~p ����T1�Y�0ܠF/�>�g��0'����C'�Ɯz�%<8E��u;�.
5����v�ɗ���.m�e8"�;�ѱrXF��=;Ul6٧��w�`�=���p��6G�֯g�M}���?+(.���UX;�Ϩt�o�<v׌�׈�w���<�w21��e�v�%�XXܶ�m��S؇�yH�[�샪=�ƫ��z{���@��@Ϳ�	��PSH�~��}�A�d,U�2#X�1wG����1z��s�M𣽼�M�،�R�&�4,��G��*Р}��T,�^/��]>����y0y�_�jĐU���y��~��Y��U�R�b�9Q���{��Ć�I��p]� �>!��-�R�yXK�Dϯb�dY�tA�F��?����K,�7K�蠎�0t�D���~=s��/]�4�J";;Y�o,�ͮ��  :'��QN�M��k�nXer�U��y��^��/�yC�vm��s�l�ꡇ�G�Vt��w��ai���4��}��օ��u���#�4w�ן��'����W�k��=�v��(ht݋�������n���zK��x��/�D��6o��D)�������!��6��e���9�m��r��!����\�ز�D�灹����ߛ�9YG��+�#)"AԅC�{?A�Z�6C��x��̜&˥�б�D��뷋�}�B�D�B�my?q�PH���������0�%ʬ�CK��q��*S�9�W�=���R��y!��"�?s�/��)��aw��Y�eV��D���MJ��W���������*!-9ŌOOLidY^��t�TE����D�o҂��4&m�埵!ܿR���0��Q'���CҸ���3}�t��)$M�"m�cI���p{������ѯ�a�S���詅Y~�_���0���X��?YD�:�c��}=�������Rt����@i!���*jH�K:.�¯ԯlO��}��!	_V�
�]��J9]22�P��ғ�A6����ݕk�;H"6Cc�����ɤ���e���>w�L6*`-��OR�2��}y�Ote*��T�H�hWk�5���������縑��5��ef����
�Z�|i�r�$���5�RIk�����-sw&.L&rQ��,vG�݆�sK>�fs�u�8���/ly۰�n{;�s����НkMf��[y�Ӯ8==�m#���q���g�뇝�z�W����֛s]�mq�v^pq�X6'�v��!���V���
�pF�z����j�p�U��v���j6��:}�\ ���i݌am¦wа��u�f��FWLc�G)�A�w#����ν5�]�:꼼���m7L �t����u���'�"�^��T,�Q6��A�4��v��9	<d��E�eM���:yt"$�ډض4�]�$*�#sո�nƞ+�>֍h���˶�ٌ��F���U�N�8ի(��Kޚ�Mǲ�";�� #�C�:�P��O�L��p��P���:nd��7��n*91��f1NupwE��:�pp�hF@a-��N6�N�}��a7�g��m ��D��ث����ǥ���Z�/4�ؾO���ϸ�!����z�+H�2���M�7{��.�iڃ�ꖭ�5�t!��y�J:423�oE��ŔC(��z�q]�Wȣ�H&����h�ك���q���"j��"���I�G�_p��[��K$�n"[((���q�*�Z\A�C�_�X��'�C"zc�5:H�lx�ˬ�d��4�I�f�N���1���6����OP��U����r�a�w�6B��|�m$��d���]���(N�N����g�94m�#��N�y�a���l�ׇ-�2f�������>��Q�������Ҍ�t
:F{/�C��x.$�V�c�E��|x����3���:CM���ui���G��ċ�s��p���&�rJ��Q��a��li��5��Y��G�TX�܃u�½�]b�Zja�l����r����<���J#d�G�:��kx���&m��eN��ԏj�`����+}����͑D�gH�o�P�_!9�	�ȯ?v�@���C���C��4�!�̎�fG�JB�e�������,V��yo��C�Jҍ$Z�!~�`�9�<ࣦC��uj���L��}4+>2p�2c��8T�8G���-"�q��o���j��г���?h��.Ut\FH}��v��uP����h��g�L�4,�͓�f���Qמ��a��k�����6W�����Fߞ�\z�%�MGs:�OטrY�(D�"$&���0p�l�(�6�7]屢8s����	9Պ�����Gܧ�P�b�ܾ���#g�2k}�k�"�D���֪��Ebj�+�.N�o��$6�O���A��r�dE��c��=������k��.�u��S����d82F��)!���V~�P�=�^���D�C�������}��(�Ѕ����6�n�=��� ���=��6_/�ts�e�m!����9��#1��E�/	��h_S@���p��jԀu�5l��ț�M#���Zq��O~>Hk�\�҄
���&�EO��5��F�椃�lp��7�8�YEK-�Z�ٯ����^EՂ0ߟ�P�A�<!��DY�PVW���ya�4|3�G�b<�0��QK�rdt��Cr�шsV�1n�Qlʤ�G�̭	��E\�dsI�����7cwA��q+���)�e��vs�Z��x�y����s�[���
���7Z��/-P�����k����A�-@����L`�Z@"��P�(��������5Y;�o��`�{�c-���d��)�\�ǫ;!ht6�hrX�Gp�����|����ɡ����dg�6m��c4V<�;�
0i���|~�1fWv��띜���E�pm�+vt���M��y��n�t1��d���/��f�ڹ�:����J9j���S�	��y^:�k7;�H/�9Z�X\��4C3���̂�eC���לD�|ʵ}5sd������{�Gj4��N4]3|5��m��{������@J�'\�r��G	��
~�k��ns�\*N��u�2�qt��a�͗W���O�����rVQ��N��z��=��;:��'nB����Y��2�f����u!��Zj�f1�oh7a�o-[ۗ*��4=�;hen�Tn�ݙ��U��:�Ƕ�bD�1/��nr�ݪ��nd�D�/Q�f7���vfY�]������x���o#kj��dNF�|'�2�eՋ�8`�$���^�ƶz�a�)-�g�ݾݖ;���Yq�r�Efi�-��(���ۂ��w��q^��Ԏ®&�N�u%v�����M�rݚ�n����b�&���XM��b����4'澛C�ޘ��=7d3��<b�L8a�i�HӐ���Ƒ��e��e����3/«E��W���St����ڒqu�ݟMeY��?�j��lV�Aq^+,�+��������y�C��0�G���cl6d1����}��d3�kWQ��g�w㗯�����X�\�u��k�(��Бï y�uPToA�2�xYk���N$A�4h��^���yz��9�Q��Aq������rG�ZW^^e۞z���wm����I�f����,���H��Ϊ���g��~�B�鍈�Yf��wz'6�7,ϊV�IY1�!��y1"e�כ�g���"-v�$D	^��{��ݍ��[��^���F��c��np[~��p�T*�q��;�/��lY���u�,I!�Ч1_.��޽��kb��}e��4���.c��<5�*�R6;�"��[��w��V`8,�',�L1���?C�&w{:f��W��z+���p[w�Z�Ǖs<���e+��{g۾S�к7Q��7]���*����(�K�.W������Mtm�CA{36�e�:�Dv�˩���y���T�uu�%��_3p�s*D���$�۞�5ǹe�W\쯨L�-�W�+Ȟ�A�L����gi�S��Yrw��G�u��z}�M��>���c�l�f���%�u��N��-ؕ�1��S�b��)�̂����E	grq�Gt�u�,��n�>�[u3��32�r��y��#1^z�sC�gEAJ,cްEE� �u�x\�	�����ce9����[���p���\��M]qo#��8��(^t�K��.���TOβ��0���Æ�fe���N�m]{P֍d/F��C�܆�Onw�|j�74���B�8��R�.و�C1��R2c��%s�2o����{[SNv92�u7C#�-\i"z�,�6q�쉶/X�mJ�z7$K;�Q)�#h�m�s2��)[W)�W{��uNru:�hm^����Lu�vܽ����\/�CL�!A6��;cu�����>`��a>���/��+\�5%i�8.��(��N��s5;�N��y��%���lR�@��F�Oa�Eʭs��j�^Ak���켹y�[g�,��qv���ݲi�,F��>�����"bK�x�x��(O�^���q6ώFs�]��m��nc;K�YG����%��8ݝ=�wWN{[�(��sq�,n���k�ͻq�bb������S ��s�ۏm�KK�cV��>F��mp�`�wN�0v��Rm^˽��6�K1�)��u˹�ZN��!Ǎ�']ek��.ۇ�Yν�����V뛆����0A��K�7��u{"�\o���@L_,��ӓ���*���	4f�N���9����3(�@����rfk�����Q�A����9�w=����Wy�I��{�}T���v�o�֙�kb��2��'$F�e�y����A��=˽7LǗ�Q�^=W����NlQ��{���.UcT2�qm����yf�0�e�Z�'�{���n��ƛ��M��@���K���:�O�g,z�2�6v;Y�s��2�`^�0LL�l�iȹms:��8q�ɬΨ9A�n�]��5�m��������y^P���:���Ρ5Sy'	�b%|U�\\�v�&v�KvιCA��Ҟ��74��.��Ąs���Z$RZ�B�Y��Qy�-�^H��Q#��;�3#J\���*�b���.w��n`B�.�l���ЌQ�I����Y������nf�PA�\
e��q;�(l֫�:m�7B����a�z*�;A���	s��,�s�sYZ��6��J��ܺ�3�u��ㅥOh�͚�IX"��W��u��e1֒�[0&ci Ӈ�s�u�ܫ^���ܯ���[�s�����L��!C��-��h�1�_^�����W�yMm�-�5���9�;�*]�yM����ȃzd���.ղD��w��
59�����4a���k�H��W�;wY9o������j��;]�ۀ��Լ�e_m���o�¿;Ц������#�s3���Fت��ҹ|80��X�[]��g>6�8woF{��m�ڍk-���m"��s{
�{��<�b�;�O3Y�j���/�{�WkB7���;c2��v��A���,���`Ĥy��Y�b���ʃ�����w**��#.�=�����)���zafV.�C�����v�r�0�O�8IJ�n,�8j�n,�ʑ���O��W�k�^�����_���m�E*�k�Cs���,��R҉�<ѭ��c�b�bȕp��6�����{�6pp�yj��^V@��HZ�˹"v*zy��:��-����$��#��!�>s��GW��V}��Uig�e؎ڗ/,�����2qZt7b��[{��Z�o�z�]��%J؆JQBQ�z�w�}�����_p��M�&d�Q����JL���xy��1����ֿ����#h�ٹ:xk5�nӗ��*�Gku�gh��kcѹ�zk�W'lT�L�12xj����ʵy*�,ַ<2�o;C�u%EgN�Λ�Y9;877zlV��.B'�C�\��ڻ�-./��X�B㭹gO�lCX��2���9�0���Ҝ���l��뎕��,/�(MH�Q�}�F�V�יw�6�}��a��km./^7�d����rc�|��[b�>�[Q�dq5rNi+�M�΄ڷ�����G�/hG�";s&�R�w��qk��T��2�t;m����p\hN8�Cb�+�C.���OV�Z��j��Z}^N h��ާf�\�Y�j@:��EAi.�5s���e�^h6.����(�NC�Ʌ�9�ss2,Ұ��Σ�_p��p_ϟ/x%��a�����䙑1�ήw����gw��CoW���jZ�B �����q��{Xs�B�웏<�xm��.ܘ,쑮��b-ȴ(��n/�:Ѷ�ۦK��Lj{���m�#���vb�Y��xWB�8�My��U1B؊�Yl�<�Tt;š�����|��f�/�z�:��_�E��Y����	��]��(/7]k�d�E[�#b�&��G��j���Lɦ��d�t�%�l��^d��K��f]Wz���=�y�}�1�a��	�E���7;t�V�6q��x�V��ɝ���J����W��H����7��������.��4s��֜q�`��p�ŉGk޴���Y#�S�BZ�n��qy<�5�.dЇn�;ޚ��2Q�y�>�0Y�:c�����.=�dܬbٻ��A�p�f]�'{wra���B��QN���̦-�Vs��t�N�?R�6�;	۶j�2����χa� ���Q�H�t�u��gwn{3�V��H[�ܖ��2�ݒn�2�7شI�n�ړ[7]�ح"�/�����^"�nE��z���֔@�C6�{�m狐�iOH���OOT����d��vt=�|�fMs��x��
.�{F�Q��]�-<n^��>��D�˱�@5��,sc��훃I��\��=���qv�_lgR�&8�'j{/sǄ�ݬQA�Cq3	L����_��1r�������\,9N��a�.g�":�'}�C&S\�<Q=���$��H����V�ٶo�h��j�]�^��|�zhR�MC�����x����l��>�(�g>���D�[3o���Y�gOn���p(n��\�!��m�/(q��<���vj�(`d�S xZ�y:^��۵��$���ֳ�.�n#\e�Y���e[�sZd�&�i�'\�]�s��ȻL��j3��0�l-{8zhfT3w+�*�TZ8猐o�4�F��B�=��Ą��k<�|qk��������⒦�@�xqlݵ�^�k���֎��<tmiw]5�f�+����d�#�3����j�8��d��҆le,����5��"��G���.�Ŏ�p�5l������Z��!h��A�&�§9��Y�����7��Q�{ֆ҄��6�ی��!�P�G��-��˼(+��ɛ���S@�s^����'�xw]�oz����X�W��7�)�.�W�<��y"R�.�Z�Pw9�:�;۬3"D)"&�F��{Gp���o�aY�N��f�M��#�[�reAso�Ԏݵoug>�X��G��s0l�`T-�'Y�;��J�E�:��ˣ�����Ssy<R��󽭺��'6���!�%t�\��
RyW����hv{0M�a�{�����<��Xj߹h�tj��=����o,J�x]�����oލݚ���+!r�Fy�&1ۘ���×v�@��E.���v���{4Ӓ"\p�!m���3�{a[��e
����bo�nY6/l�W�
�:�CT|`�V9���%��8�b��*TɋÙd]���z؝��a��7��q疞��hV̩��oͼَ
�~�U�j��-�Tx5f�}T���$dyf��_I�^�{G���2D��Њ�+�z��	&����ۥ.��)	���α�����������]���g:�H��k7������4�{Pu�u�{'���aE�cس�=� �"��sY,���n����uܶ#���O2k�ck�z/.��������֞C��%9�6�wˣ\����u��N����p��2_{˵�85�`�\p���e�=�x�ib� �:cW-�^�?����#�o'��n��Y]G]_eB��g�
�\u�W*V��qxT��\<7k�\����Mfчʺ�W�\h���<����V׽w�Sس�y �U"���@h�c�Z�B�7g��8��ѳ���NZB�d�*�2+#�������,�|�Yț�?	����t�6�J����.��PK�&3a�z �]�D4LQ��f	 ��+w��(읝�Kwtf���)(��1ϯk�z^��nv�f}/�7��6�k!�6�E$�����)�n�om�E��a��!��3o�:貱��(�;�u�98iV.�I%u�tw�
�܌��٢�eZ.�Gl�7q��a�v��r�j�/NVgp�:�*Mc�w8���jCH�d�>�����K�<�N��P�Hr��Th�N��^ח���X��e�yf;�&�.�_��)�V߳O��v��y���l*�
���o�o��q��"u ��������R��v.)���JRX��?s�yOI�{�t��8/hg{�D�ۜ��=�e��+�=��x{ͬ��(,uЊp/���d��f^�b�;���/�fj;��p>��4.���n0U����-��"��x" =\������Fݶ�������S���1MEw�+=38����������a��05���`�&�K]c�2 �2ap��M�s�Jݢ8rŻmm�ӧ9K+E>�r�8L�VmҬ1B���K[}o�6��i�SʻC�Y8���1p��jFb�c�9�;�ͼ�v,�9���t�;���,K�L�g2J�Ƞl����nca!���m���ߕ���5�
������3�I2�Q�����K,�����X��	��+���Ѓv�ʶ=�uY��X�E>
�e�R�Z������	��Z2�»�%b}�<���H�ϱ��j9}clӲ闦8�+�+�dr�����v��qZ��/��J���3q��͎�h��J�Cݾ�1�bl��j�^H��qUi|�e�ȳ���0�g�,������Zz:�[Ŧu>�'���Է�NUA�)��0�_hw�k$��6�۔ic�h�v���ByH��ɢ�3�۠:=Y�4��E�Θ��e��r�IɁ���gr�yx���J��W���[��v�Q��ۗo`!oRk��Ž���Pee��T4�]L��A0��m���h�\F�әUzحi�\��M
f�,���3��w�]�z�5�9V��NbDb�ٷfr�P]y��X��abئ����,�>�˽�XI��6�o}�/(30J�Ts Y���M�m��S�oJQP�ae�ɈR/TZq�f�n(j����*�cN`���ҡ\�^)�d��;Fn��G��g�ŻM2�vV�fj7���L��,�rZh(�����&�s��1=��9�U -�|X�N�źuh�]��eμ�1���/1j۬G1��+���Cr�
��P�q����v�Z1G֫�o���6�*�4rZw���2Gx]�a�7n�꙳C�k.CH�/3C֎�����H��P�K/skJ�be���I$X*���Jb�lH6�@i0�*���f�c;cAJ9���s���4�iI�Tee[�f�n�
:�B��컧��&v��C���Guqٹuqۮ�z�|U�r]�����!A�j-��ыs[�X�"�/e��ǯL=��v��=��z����m��㴻"��̻���OnP���ۃ��NnN�F7h��4��;����]�0H�ݧ�x���m]�&�r�Adǎ�W�t鉻��4gnmv\�Ƹp�ǒ�W#=p��V�*:�R�2�f�k���i]�lנƺ�w=r��h^�ێ[F�3�烷�+p)�[p�7��G\A��E�g���k5s�{x�v�;���Ӯ�wӰ�����n�1��g��r�;@��=��l�C��s�z#c���A'�X�g�s�=���<댡���/;7m�k��Ra�c��S��H��ce�y�	�g=�ԃ��x�]�&�.;g�n�v��ݗ<1Ɋlv:oZ�����;GZ�t<���3FӇ�8�[�m��b�!yU�0`�㰱[v���ֲ�I�t�qQ��v�W=c�v��B��&,��4=v ��\�ڌ<�����lf�G˺N�:0�q�`�{z�]pݜ!��[[�jvM���İvsr^C;[9i�6y�(WnS�i�t6��<[�pv�]�v�N;P3�k��\Y���RH�n���½)X��#[{Xd�Z���<<ֱ#��g�۬M�Igg9��f;n�.�6����۸�^����Il;�M=�vB�8��<[#۶'UӜ6�:ݲn�D��m19��	���^M�&��-��c�l�S�q:8y��aűi�n@��oc��ӦSq;���v�b�7Wls�mZ\��=���c��w^��'Y����:Eg�����GO�g��nۓ��;=u���4�8����׶#Hښ��=�$����f(�8G=�<M�z�G=�����C��x=�8��c��s�`zpMne�#�	�۱��m����p+q�ks�6�����c�;��s�-���Vi��b�أ���+T���ݶ�T�;<%�=mM�ب;sv#u��K<k����;�����ͤc�|n�[����uG;A��\�p��R��Ʋ�p�՚���O7��l&��x�ך�\(ގ�!����kkl�gWl��#r�V��e�ƻ[��!��潃;(�qc�Ϯ�tc����a��ɶ#<�P������!����ĩ�3����/(\�v���`,�ϭ���m�}ٸ�}\�����l��,c�':���m��c�`��.��^�}����V���kٌ��ڊ{ث�]�ʻ:��
b�d��itn�>��`2H���rs8�>��������jZ����N�����4l�.�vDNi�=���H].ۑt5`Q
��9l���Ɂ}�kog�oW�������x�M��r���v��G%��"�a��c�C��#�^[$S��;c"7\/hN|�s����"ule6�.��u{9����S�R�*�z��8��B���3��ţ��\�����r,�$�Q1�/��@��o"���қ���Se�ǼE1���\΅Ӱ/����j ^s��w;8�<�VՇN�I���U��E��呵�l��W��N�~�t��d���""�K}���%z��[��7�ajy�����%j�̯i �z�����.���B��]�^p((:Ϝ$Q}j��[�V���Tu��s�h�o���Y}�q.���V����$�����Ǻ^p!wWQ�z�:c�٤��KHK{ҥ�#+ж0���0��5���v]墷M�	��o��;U�w�+�r5#�)��Z�7��	ss�^�rQ��z)��;UbV��|���/���7����n��I��H��
$�#3��jlU)����rW9M�y�Xǵ}�hi�|'a~��2�d}���P,g�<55��>�XHHF����;�~��mLY--�~ϰ�jׯ/��]Oy�e�	�/n�Š��9-W�o#�2��3��u�ꖷ$����7J0�%�Ӆ��L�l�u�Sۧ�9(ñss�8�q0�+��4]+����ݢ���d�`7�M�od�W$����Qd��"���g���{�4���K!k��ױ׎p�17;�Y�.>l�	���G#����:���8d���8g�ݶըc���)��-�|j�/���<�ou	z���m��A.�B�AVZ�>
�'-cw6����E3t2��
��tv�ݗ�6,m=�y�{��0=۫Ȇj���Bb��:a���h�Nw���o�����ɓR�%0����9�;%�p��U�\��L:�K՝�+b�q��e�)��}�#)̝�Yݷ��>�/\p��0�p6���(�[��W�6f.R��<�-��k(��,�afTR�ѼSRFMLg��Y	��!(*��?�[`��7l���n�;���y��⁫�7#�v4]�Z�*bC� ���K�̴�����f�}�[��y;�j�܅��ވ�ۊ�9C`!���8Bf3#*@\
CQ�q��w��g���Mv6�^��k�{2��l�ma���y ���MY{�j
z�m�"��2H���rg�ۺ���}��L��B2%cqMl�7��U��29��8�뾺Ǚj�*�y���%0�RS2ci7-Nm�w%Hy��s�T���!�-Kq�� ������F%t�+�RJ��!�f�j���̲��f��w;�겚�|\.�=���	Y��t�Z���}�e��ϐٔ3x	�=����yc���r��VVYd��k{�C���KP�M�t�[üq_rܰ�i���yt�D�y9�X�m���*!Ʒ͟iZIT��:��i��JF݇�jluў���h6�_����E����]��ܑ��1Zwܫ��3+@�n��3��Ҹ\A��p��	��f~������1;���t�Bx��`��S|�a�����)mb�=�v���d*Uֈ4��;t���-^���8Tꂗ=�p^X����
j �2pw3%��ܫ�Q�''C�B6�isL����3[}��O^�@#i|�U��\b��bP��3AP��1c4�d��;ao�̱y�b��^ϗg��3;Θ�oqˬ�N9����[�Z�n�0	w�6eY˵A�'O�v\�=�Z
��vi�6f+�[����˿z1%ܙW��,g�P�w���ܮ�ˠ��
��v5\�v��wM�.+46��(9C.�sZmfC�ɕ�֗"%u����]or�ê���3�]�o�_���$��������(�ٍ�����v���m�^�u�E��7�^^�ٹ<��	8��m�a�VH�yݬ�v8���vy]R\f��ǧt����g����wQ��:9���o=�l8�����tVю;m�Q�U�5u�n:��y�$����4�nɧOVn^y*�vyҦ��`;k��b7W���lۣ���/=�0�F}I��~�����tdOQ�b۝e���n���Iw[��Nj�<:��n^&�w]�{/=�D�ѧ�c=P"�U����~u5N��2��nm��C'�c�=°.n�*M�|��q��[�.� ��h�"Ϭ��9u7��;0��{��vXt*w��L,��r�vVS�x'2�C1u�F�%���q%H2%	)JÆ�-��o��
f���}=<�Eaʛ=@����wbɕ:_�y:<W���p�P���ZrY��Y�ú�����ȇV������ձ�����븾��&С�1��dZ�Ȫ�5`�2iggsP�q�R��KǓ.����fM%��NCn����R���ܹu�_vu�{�rt2����6T�=��<Ƕ�C�n��&֚�|#ۧ�U�b7]nr肄�O�ꔕ;*��{�"����M��d�]�c!X9S��.VV7�_a�q~۽58����d�e�r��)!�ʧ�y}���32vӦWd��%�-�arsO���Wo���uP�!�qs�NYv�+�1��8�mnʼ�j2!��YoC�Q�W
Kn���Y)�7r�vw�q4ۭ���Wu�A�O�(��v�d��*$���M�=��f�qM�{��x,[@Wép������R�:�.�i��]Q$P9m�%rqb�|���gs=X��18"R3���Cj��q/�U�Q����.hӾչ���`��[IS0�,��Ii�^w٧��h�-�V}OK[v!��D�{VW��{Q��k�%�H���L�]�{1ɩ�d+-���E�p�q�n4%�gw7&[���%��q��i�{=B��DH�m�����Kd�o�ߵ���M�O�]c���ni�;����^f�����mf�z �W�Nǳ}.�
9wwxE�l]�e�M�ſ{{����i����8�Q�$�Y��Mm��o�5VV�o@�#f�ּ*0�+�dI�1	|��l�~��ގ�v��y����T�~�Hn����N��G����Z`��Lm�}�Nb�3�r��}2rpF��հ��e��ֵ��t%��z��V�v�\�9E�}a�Z�o��Z����[�	ݍ�b-2� �A�ի��;��R�<�`=���zk��� ��oo ��Ŋ��mS��v���K;qvC��HxS%�i|[I��:��p)�[�x�`˨������3�n�R>�XF׆߂x�r��q��`�k:�tQ�٢i p�c�7Vhy���Q�I$�:tE�.��D�\lݳ����'kWi-F�p�]�ߟ�fT�֞+fwW"�m���MGXT����/2]��Y�)~��Ω���cdL��Q)7���{Yf�@�����С��bV��ܫ�;��7�l�Nm-l�2�O:�s���g��V�I(�>��xf��ae���=��i�{��a��ñ�}t��-� ܮ.nZ�����c�*,�}]���t
f���dr�:�3�����kb��z]\�1g��B���^v���!��{�K�zS/���֙vG�^[*��*j���{�`�ʼ��V�<����JS�j��{cx�2�[�}pd\=Q�
X��5�)"q�Kq�w*�s��S�2vv�0�lk���d��ʁ�4�k��e�I6�yǵ�e�����ڿV8;-�04�(&1��un�<����͟ �ې�'\�.#���U���PZ㲜�ީ���˳J]�.]�݈Q�M���Xz¦�֭f7�ytk���nΠ���wGϲ� 9"D���2*T�>q���E�co����ɺ�;�Dy b%ޚ�S����_hn�������2Ԑ�	�3�zi���ypR�t�n�9�;�F`��r⹸�7��~l���4
�/0��`��1c�\�׋�	'�.T�u�~Ge����l��5�����	;�w��v,vj=q!p��i�/���|�S�R�:��@���q[۴�kת�T�꘡nzFwzPܱ���|h�����o㠼uv��g/I��0��bYgz�]��:���H���x {\P��j��ze�d���X�(��n�c�Δ�slo;v�X�.7;�ln��7d-g�����9�����c�������uֱ�fy�b�=n,��Xヘy�ɹV��}Ms��Uyg���yw2+�p=ۅ��ܫ� ێٜ�+�N�1˩؂�ݸ��|����jݺ��O��8u���moL����^�gv�:�tn]q���0id8G��9Ɵ��w��ܫ��h���aNI�nr(��n5qqɸ%�:�y(d��Ձ[u��䷎�Tsl���B�.E�yѣ�zC9�a*e��<�X�����s��ɥ�ot�ܠ�|���npꁱ1H\R<��`���6�Y*���l����5��Ӟ��n��bq�Ϟ���I����<lt
LA-�䎄�v�^���s����h�1:�ʸ�Zj��:r�+1��ھ��ԳY�s�o�U���IH`)"�N�Q��ѱ��A�Mmݶ���7"�'�<YWݶ�t��F���bs!t}-�Ks�gN�U�)Oҙe��1�|s�ox���XwB��u�����f�H�����=�֨�n��=MF��2���[�%cmxJh�$��<��ݭ�{k�	g�Ǒ�ݶ(���uu"��ה6q%�m �r��]N�r�K�vn���s|e�]efT�VM�)[Dvb��εO�u��r�|L�[,e�ϲrWՉ猅`ς�����[��l�ٱ=���F�0+���n鳝u��)��]��;�V[��x�)�Z<�þW:���s�ِͬf��5��Ŭg��5�����ok���]�a �l�����~�=�e�v�f)&T�x���"�c���^z�Y�oy｢6�<��>�-�,0�C+냲S[�4�kb��:w���b�׎1�},Oj-M��<6W|���V�{�t"�l�[�w���)�P)#�����C�91�\oΞ�����+Y��i	}�/��O:�SA/q\!��W�hx/�'�Ź��U�ok��v�'����O3�X�;sT��^�vm'Q�����}�;��7�uɓÕ��^�٬���y���ڃ����p��{�*�C����%�C{��F
��18!�.�y'z�io�l��xjz�OvX�]39t:��m�v�j�K���.1���<���<�r�6L��7M�yᎥf��rS��^��]~@���8�=���Y}�\%�\���ߺ�
�@��M���W/���5G�jn�]�mw4��b�Z�|��Xo�'H�=�q�E�nf��:��߮%H���Cu����6)�B������c:��U�11h%�1����F�-��Y�����z,ޡ��ڻ�����(<)�v�v�#]6�s�"�\���*��.襵�vbĀ�\>(�f�1^wwLe��_v&�������]��1�AM1�[�i]a�c�짜��_$ҽCvL�؄o:nýB��c�V�sE�V\��5vFV�.��]�}rɾO,9�Ͳ{��c6u�3WV`�EX"�ǐO�ཌྷʉC�ʃ��)\ɖ�A�F==0Zdծ�F�pS�Y�b�^�|6s�N���ko�5�lMŬn���')�`Yy�9�m1aM3���"�fԺ��|��#�zq��Xy�`�/�-�Cˑ��%�*r�Z�<u�v~�[�H���\��ݭsX�R�h������d�1����(p�i	��,�73I훜��f� 4���ز�>�%G �nܽ��0�ԗ�,!L&sxs�A�1ؘ�I��Ǜ-�EGLNc�o2����*�Yݔ�v�b�}�e="��x;Y�
�f��;�.�|J�Y� �9�f��_n�'���4��.�p�f6_K�&������b����Ȱ��a;|vހ�s��D�Ż����7*�fXV�ۗݫ�'Y+<V��l��>R������Y�m�ܲeݖ��-�KRzsM����晼��ܙ0��9��1�.A�����j'eC�iw8����q��w0o��mCqxp���a�k�UTV}�w�4^�T1pH��f`xF`�����)���㠖{ޮ�gS?pܶ�X]��z-��C$��Ru��M�*�se�&G>�v3�g'0s���:��rT�k�3^-����%ϊ
��f1[���驟���nu/f��[V�d�ڸ�E�ekB%���W{��5՗r�m����4�H�q�!H�J�3'�lC���gjG$��c�[�2�z���~��>���*��v�>u��'n�rg�$��5#ۼ�}l���y0�ە����i&8�m,G�vc����]͑�M5�tn�2[-��k'^��'03�@�3]�m�d�Ӷ��e�3i꣥��m�QN�."�hL�CU�=�J�]8GI�X"�����ޚ���]9��ڗ|�.Ti��-�e�o�f��7yLξ|;4{����[s�,���F�DD����o��F̹3�˞���v���ur���F�kg]��V�uaܬƪ]N�8�|�s�8d�7�g�C��oG��s͋nTΉ��u�Sm�P��υ`�2"����e]�ͭ�����e8e]F�L�Q;u�3%���KTVUN��0@�ʵB>���~�#b�(�9!|[!�����Y���]�n9£#XZ�{fvum�\�/ʎ���:��� �Nz�
ToPށ+T�����&d�!DL2n�p�1T�c�����ڼ�%�{|���4*�8=*)�K�����;�����nP�E([7��&�=]
^�|����R"����c���]�+��e�x7є__G+ݒa����Lc�"��u�Y%��.uy�GP��sW`��j�N�Ys�1������SY�߳1����<�7�S���fW	�T���z�%ra�����L�:�+m�׊����g7���ЛsR�Wj����Z�r�b���o��t����ӹ<��p]�8�PI�F��fI�(lsb��'��:��&���pm�[O\y�&7�Bڹ"1�\4z�gq����=��ֳ;jÌ�V�F����qĔvi�m˷b�l�9�:�m�n��6�2��cěQ;����(i��`P��������雮�����ۀo5ýc��uC>9n:6�n�I�ӛ[�p�wE*�i��;yي��R�j-N��V��f�=u�Kv���u�k\�{mc$�����p��R;�眯-�U�wO3݋��v[�����
��K7}}��3Y���oOq��{�kq��	e(]�x��?�h^��k��7o�X�Y� �E;%X�5�����MJ�����ʆ�h��(; ��ʽ ��_8d����M�����
�7���OZ�hq��rx�<��y[���l�����f��'TD��KT�אޜ����um>�z�mN����}�Xqӏ��Ҧ7P�P̧�c�w������67��n����loc���}S��!�������T;F��m�*�G�6+�<u�h�^� x�ˡۍ�޹YcƢ���bj7Tb�ônm���<#�rm�l�ͺ�%�n�[��Mj��#��N�G^\��x���V=y��EtQ��NYU����V6�[b��}��'8�m��n�F�m�&�Rٗ����Q�~��o��	�ůXv��	R�z�y� m8��� ����I�V�X�S�v���\z��[���X�u�<�Yb^Yz�kf�wM5��/��5���b�xSf�m�ӑ$Ԏ�C�Ju�챎����;�#��*��}p^�ٽQ%��� ��f�Ѷ���x?L�*qR�HKy�;K���k�}�C��f��COY=.,Ee��̖�!~�)B���O/fn,�^�n��Q9B�]���	�ׅ���#�K)6˨)M�vc"�6��ֳ������rx�'��!�O���c,�`��4�K�rGU=��.� �=q�.�nǫvs^�u�Ɋ(�RY󱺚"�e�^��.v��jjn#u�A���>K�/*n&�$�O�9��ˎvə���Ia�Be@��w������q��{7׮�5��xW=$�q��)���^X�_�I�r�3������ȰX���VY��d���\U�ᵲ3�O�����%w.uF�3u+��:�NS��&�őV:�K�&`�C�l�S7%���s���*��;���H����b��H~?)WK9 5�2[�W��hr�}J�^���Ży�Es��1&F���0)m���}���=�QKY�s�:z��{-�K3w��Vٮ���}/s�I935��^�>���=P��ߘ9F@fI+����O�8e�.�E<� r��um��"����Y3n�w�{'���[n��߯��;�-�[9��#I��ֻ��r�p���Üכ��W��#�N��ѹg=�� �e�g:���)��\���!����'ܽ��ʼ��O_F-���g:|�p+Ϟ3Y�B�%u
����l�oe��s"��;��JZ�l�Xض��d��]NR��w�s��{~ݫjE^�p=��b�w
�u"+�i�Y-��Wr]��S�+�m�3��K�z�8Ib�ƯZ}/m1�u4�KE��6o�W���y��b�D��|�޾.���ݡt�v���n��J��U���f�o����s4R�'w�ǩ��%�>[�����q�#�K�,�rl�9�l|���{Oa:+�S�z����+�����[��jhD�h��i]�ݾ��
�D�v�X}x3�7yRQ�tu��z�<sPw��x�B���RVQ݇]s���h�R�.Ttn�[qsU�9ǊY�'�(2��m���e�����>�fwW��/Gf۵mU�ٱ��M����-k���j[���?L�ӝ�N��[8�h>~�hY�h��OsWR/�]�0��>��̂�n"+����S��\�0�`u9�Z�f�n9j�a��(�=������\�v��n�H�zy��%F����EBї����a9Y��bba�G�A}`�e
qmK��"�w���9�r�w�3��Z�P��=����d��%%�\�y"v�.����tn�<�伜�9-I͈�	�9�&�1���f3�®K*�۶3D�0\j�Q��q�3�(�i��T
B�eX��]mƋ���o#,�����N
�w|�wMr�Һ�c��Z��^+N�ۗP��#Kr�dm=.���m͊�T,��U��9W�Y���8�h�$��ggMK�L�o�j,{v �`��C�m�mPV值�CcV��Oh�v�պ��n3��g�ݎvͮ��Z	�ol�,L7�h��麷Y0䋳n��>;��X�\t�f��om������|q�<l3�h���k#�z�.W�հ=kQr�닋'o>֒�8�qw,myuN�N��}��}��oki��8:���3������6���%�'1głK�׋&�o^+*���Ql�@�볍ی�V1����
�r��Xv����f�r.�hNGY�=��a�@*����2�޿N��Kh�O���O9�x�r��&�{�'ݐs5�۽����vэA�-��������o��T8���e�&ک�St'wW��]�n65UN
!W�ns�A�pD��e���/
22O��c��5��.���sNH�7�Y������2a\���^�o�S�-�y�+hekC1-�Ƽ��a�D��ף���W�{]�����\��l������N�L��l���'/gbo�K��%V��!��HB��Q�`��8*;�����2r�N��eI�x�_B�O6���1\�|�u�q�r�|����[z�z&����<��m�֛���l��ݹ�G��A���Gn�B*ed�ٞ�o޶a�|����~~�n#R�4u����]]�S9w}g��31q��K���F��I�̑�.��ވ?}���}~u���
	�Y,���S�ɔ��*�Z��>�eǩ�[2��8�S˕�v���)�\�v�U���mr�2G�g�3�O-�;�Mp�:���j+L�;�f���d�N�}�2Z12V[Y-���&<�� [���z�f����f�ѯ�B��9u�w�z68v�ZO_x9#h��%�a-Ǜ��+Q4<߸�y�T�p����̧��7�כۡ}:�{{���G�f�+5��-^3#l���lv��Kc�0�2����9���Ý��7��{�ڬ����{m�d�f{e�,��~��S���h}��r�~�ksp/nU��N9n�+���p/Z�4�mu�C��q'WҺ�z��LH�^D�.n3M�	�͛�M��Y��������{:��b��Q��^ٍǫ�ܼ�*�al"��J�]�U̘����pLb�.W7V����[�N&6�̹d:ٹ���Ȭ�K"a=��K`�'-��eE����\�9E�Yr���d�b�_8��s���9�Ɂ��v�I����(g"�R�jݝY�#W�-�Ջ�eB���OgU���^�Z*����Ewo�N0�����9��s��»�;�V����B�Z�"��JI�8�8*�9���<��z,fS�����/w��[�W��iV��.F=R�;.O=�NћE|� DDI�� �̶���7���qO��S,���^v�����:׳cF��U����>��ٴ(VP��X�Q��d5��6K���^فDe=qpU�LG@�\������0�( 2(�GM�����U��S�ƭ��[���.oc�����1�f3%<÷��!� �=;e��(�r0ٱy�o��}�[~�d�60���e��lQNA��6��9M��v59������ݨt�}���%�g�&H�����I׏�Z�����F*V�V��=�w/�������e��tl�~{���;>�c衍}��c6��G�n�a[m}�VT�7%��8��"&�w^���{�\��6���v��uEA����8I���*+���Yǯ�%��w�S�c�D1�3��Hӌ^��37�޺��D��;�U���4H�^�aQKۇ�IHeSCv�= ����A?�rk�d��:�خ���(.�kI�[��(��F�<���ҔY�J�S�p�<1f�Ǜ��x�����Ρ�m�QM'I��ö��cM�g��5�n;s���7j/g���3!���H&&	p��kw��f��j���qj�Y��۞��k'��_E��]�́X��od!H�Jff��m"��07�˩�v6Z��:���f��Jb�MD��s_v�ұ����3�����zTi6�R�iG&d��1��z3�4U�B�۝��ۖ2y����B��:^r���1�T��Z;���ɾo�����"dt���-����N\���]Μ�94ܼɋ!9Bz�����n�0���9G�����p>��R���q6b
0K��[��+��[���M�2�=|�*���mOmln��������3ܳȽ���IW�__�i��'g��$u�n�Ǫ�R�:KokE�����+y^+�`�p٩[�.=��E�qD���3�;����q�Rt���o��wC޻Z���_=5���m��/e�ی9u����ֳW/!�,�*_k}��f�ƛ�ʊ��6'��ewu��������b9G�3WǷ�>F�iH���w����ĳB��Wӊ4�!z&\����whH4%ź�̅i;YGN�3eÃ�-�5�W�7�.�4�#}(��e�kw4��z�5�,ݢH�sr|�WRy]����նg^�ٯ�l�=�]|�Gc���{P�Qrf���/H%�Ś�s�+ql�t�I��������O;a�f*F���2:�PnA+o7^ˣ8�T�[��ͬ�G�:�ŋA���e���&�'W.͹݊�ȫJ���<�k�4X�(e��!�J�[�F�5q���ڡP7)� \���VA,fnE�;�wX��+r��F:�I���f�g:G�XZ�/,s�cv	�T�M�Ǘ0�y%GC����������ʓ��ҧkK����ʠ�t��Eh!j|�Ӆ���E����Ʉ<y]��T3��h���I��}xn^�/��+U�i����ﯞr�����ֻ����i��vV-+��5���[��|;Y����VLw�����u⒛�|�n�YGzQ�]#�����dj�Yz��Tz�tɵk����D�*������z����.��`+*�+� Y,���[+#.�, "<;�g;C�}�E���$^��؉�
������6�t�5m2W�m"�n��'�+�0�:�T�2i�p���wgѠ�]eHN)x���q����q�og.��tp�#w;�ߕu���N�fm&�"ۣ�����ݜ��㶻=�F����-�����Y�u�����8z��#��nښv�ex��uu��;��9��띵�1p�<��;��Ne��s�b��;a�^Nޑ�[����:���tq[H=v�j1���f���f�T�.w|��X�vݩi�Ȇ5��n�7!��彥���}��^5ɻ2<�=��u;n�+���@h�����f�Lh8���]�Y����mvs���Ol`��D�3����q8�4��
��2i�Avz��e��ad��Ԝ�����v��1����DA����T�\���[�.�\R��9#�vŲuEk���H��.�Nˎ.���t��6ǎ�W؎�(��4�2���ݛ]�y�m�s���n���#Ve������e*�δnn�\h^��OK�hx8�nuؗQßh��r�c��J=0�݆L1�n���\�ێ�J��v��=��+[���=;��FI��mB�6�vpV�9.7f�룊�W+֗���.Z���׌�mt�A/�ґ%<�*�{7A�wX{rlu�����ݗ�Q��
2�֡۸�=%�"r��.yMQ#ۺ�sF��xlc��NIM�xw]j���o)\8�r@�ϕ874��&v����[[Gn���y��v�]T�W���B��Z�q��k�m튷�י�eL�c	!{=�;�m.����������;EY9��������]\�����=��ʷ��7vN��*�q:p=���9�u�]��;��]\��[�^�f��v�����Ǟ��.�Z�$\���Mv�M����_|Qw�cD�$m<q��g=<��\��Q�u���s�j]&y�T�NU�n��9�u���˭������nsv��;�9��J���cY�PNBb}�xs�n��l�g���SGUu�ۮ���[�v������N-�nۑ���s��vV�-us�q���D� �=c��\�uΞ�rM���7T��kv�"�ٍ�=һS\��2]�7V�N汗�����9:�٣��쉯ay�/������*�U�[;R��.�YLێn֋c⽾���Imy�㰏C4��m 7cn�S����t�7n�����u�6��y�N��:��,�W]Ë#��O�$��$jD㽺�ϻ�9ڹ=y_Qʲ���B��(�ۑζ�8��3�U��i��\�Y�끗D)>QĢn�>��V����	�^q>3^�O��ߝm�[���G��&�s��1��H�V(�����o��v�V�UR�k΁v!)�P��\$dљK�^��Þ8D>��f�z:��K�\�m��e����������Z�+v�(�Mv��ݘ�7U����¶���um?I�~�����R�<�=x��E�fg9�p���K��.����eG���Y�z4�UTi�v����J��m��NP�C=㲝K�P+�-���c�7!��mFn����X@�($�d�!��ݔ�lnW���*o[k�a��qq�u���睸�&�BF��'5�i�r�5�Y���^�莅u/dv]�1�˙��	�v6^b0/L����6.!��r��J[5�r��+��lp��+s ��D{;�Z�z,�"�U�]*����g�%�l>�:����y�"�v:�d�b����33X7�6��()�����)�♧�⡺q�)슉i��d�W^Q���pVκ>��f�G�k��1T�P��� ����>k�����DD�3Q�2A�K�ۀ*72�=��\�nzW�R\�s�氞ʧ�|hXD+�%���/E-��
|�P��)��b.ދ���t��&�~���E��S��������*��mu�Di&�F�u�Vμ^ݷ��=H��C��w��K7��WQMӗ�׳�X�=ޛ�\�T:���W��H��������RW.���qqW'V���h����&���W��eN�%/���_7�=K���@�Q[
�1Zh�w��T����w��#���֯>��o�����<J�S����_!�<�XIQEuJ��{G��'[��J�Ƨ	vF���}�)]v���B�T̹{��p{VRP���eE6��D����P-��&I9�+)S��n$Zʏ�kq�v�9"�]M�����a�sÏ�*bPh����&��2.y�+_u��Գ4��Xs%�N+���N��G��������_��M[:DKw=�b�r'9�c�����7P�Wc.��L��'�{�|���By�<�#X�uL��>�J˱�-x��u�]�
���Q�A6@��5�ldH�C(�de9_k`#7���k2	�v��r�i׻9����������ɛ}��I��#k�/���
w��:QXn3��pP�[-Z�g]�k��2�����6̛���T��5���|������pvLKssC1�7�M��抧�gO��\�c�:-tb���i}[K��j9�\��f.���P�S/���o;�sÇ���,�'��ꏅѯ^H�:�}����,gh���n���6E[��@�E��j��D��$B9	q�X��
v�9��T�#�:�X1^:R�'�43e奍��v��ӿzj&)�����L��v�J�%����}�!�u����N�v�8TE5�bprw+3�܉�p�BcE�/2����:)���XosA�e̔D�7 ��wf����b��78B�M��ǽ{�n��W�j�//EǼ�Rh8\�0�0�������鼙�]�&���d�� p89n�]�]>sap���X��R��8��nj�"9�j�jsg"��;F��#,[-����\�)�1�܌���$`-w�-�y	Gph�Ӆ]W�îL�n�vid����RIg��9>E.�o�30�wq��s��_Z�F���3z/F1���!T��јˇA��� {y;��8H�M��JL����WS�2b���C+���ٌ�F�8�t�Ov(fC���2~���3T�tX�v޻�L�ro�.�n�i�$q��m�ƣ���mvQ�v2]+;�^ͥ�3����h��Wk�+���Ķ�޷��諤
��|�a����>)��BI}���d���|�U�⃭�4:;��FQR6↟�����Z5��F���'��_���/2���8�,ܜȮ� �]λu�(��\�,��5���N��.��~Ҝ��������R�O=�|jY��?F��j��n9���5��ˁCVem�ZvT��1,tܘ,qgu�5�:�¥BÁ�-*�gG3�Q��9/4豮���8�@�A�p��� r$v�C��k;����u�u�ϻ<Ѻ���jy���uexq2���Ј�u���Z��sJ�ȔF�Խ��՞x�����;m��������76���/cɷ��;q��;��u���Vہ�l��6w��\�j����vH�y����?o���3s��Y�=K�B{:<!�V�ιΛ�ñ�#�z+<�9�u�Ď���[s���z�J�xۇZ�é�p���F��Nb����mu<U�=-�!��F4�M���xs-����sӱ�qe���v�f�&���0�\L������&�la١h��T��J�i�4)�e�k�Z��׮z����zD��DY�u��k���Di��6�p6*XXZ��"~�گ
U��5'�z�h�gZ
B���&	n.�֎g D�Wy/"����J�!%^E��O$�Wtލ$����Y]>=g���5��gu[�o����H���ffi3�Y磕�1�B�������ESn7o6ڌ��8f�W�j���\��d���kn���/]}�lX�;3�����r+�q֭�����3#'��#�#`���z���N�k����	hmیdX~�"�	�<���\m���n|�T����Z�u�i���P�F�:�E�J��F��N ��Qp��j0�iP4Eg�E�h���oH�ڛv�؞	5��y�<��e��w�9'���Y��}��N�}G��r?�)$FJ��(��B"����#4����=��t�\8rۗ��;�hܚwm���X��i�˷�+k(p��[�����%mtw�Yζ�]��Û{��q�a��b9(����t݂�9gv���<k0�����k[���>���Kl#�2Y&/zl0��ܞ�t��ᦦi�mgs��om����v�v��d���{���u���P�r܆�3�h�q�������qu�^��(N���k !���_ݘ��"���P��_*õ�Q�:�Yn#"��/"��s�}�ڊ�t����D���v���g1��h˜��X4�cuJe�{E�o)�H=qH��6t{F/f�r�J=��+�wI��(l��w3�����rP�Uړ��ɨ����bR-7Ӹ,��P�]+�9((���2OO�r�ɹ�;!F́�����AG-��rh�2�vqi�f��,c�s9�꫇�2�����v3��Xui���rM�C��Bb�s�þ�����(ې�;�e8F�	!�U�2E2�e¨�޼�����w���O�I�U-��&��D��� �j�o!��wݎ��ü2w˦�W&�,�9&<W�mn�.�9j�/NX˻it&�pE"N	$�.����z4|�4�E^Q4~���d��TyR�'$�	���M:����G�s�X�z�e��UX; ��fe*�b�N�f�>؞���?NH��ehcGdD]c��x�nQ��e�F����כ�H؞R��RR֨�	�@K�W���T�Z�_F���:ۧ���<f2�3�2�g�PT"�Lf3�/ݷ�����3�yY��
FgL�7��}K�2�Ӳ�zh%ֱ�l�[aD�%I[:o{״`k�!X�gb�]HLz�Y���*��b���{U�Ӄ�w�n`Λtc흮�X������Ah ��16�M�����P2���MӚ�Nmh��;&���{<���ڈ�h��NPf��?�T�8�MYTɾ�7-���S��E��j)�9��Ef�Y.�\%���7c�b���1��K5�/�>���!{�.g+�@w�rP�\UD�B�����Fm���ώvF.�\���k* �^KW�p��x4�D�A�ꅳA�1ɳ�٧����ʌU���Ź�f�yH���_Ʃݧ�����19�zv��F���3q��J�/��6*X���3vI���ø��c��>.�צ�n��b"r:盋`7Q��"�Y�T��w��Z=��\c�2�g��~Ӳ˵}�P�U�F��?c4=�t�ȫ3-1Bn�OS����ux��nH��;�y��r��0a��I���}E�[�݇Y�NUvvV��������Bq'�p➇�s'"ڒ7�����x�5#��Fbq_�6?�z<��e��n��\��q���y��1��26)���юY�2���
yO��$-��BَC����9/��#9�^��ڝ�ɨ�OC]���ȩ��t����}n�p]�����s�څ�4���0�LpA���Fm�H"%�����c7CcU��Ӯ� �ݗl��n�[���=�QK�F��E,gp�>�F��2�+�ɱ�T��fw)̓�*M"�r�֢�,.�;�ưNɩ�&�ʰu�b�-�cCŲ����-$p:�]:� ���XH�,�\�����c���1��1e�M�����h�s�rn=<s���σ�L6{Křq�����Q��vN��3m��1�<~����4�6����[�v	���,��]v�m�˞ݵk1հ�����B̠m�dn��85(8���-�� �6Ζ�ۜ�Z8��&�^��G�]�ܝ��ڽ]��l໩�5>Imv�§Y���سȼjYa'ay�랎y���<B1)��l�]�<lq�w]��̝��'��D:�Rp��C�0�.�]g(+�ԨblQ	�F��ݮ����G
�UN����'�S�8Hҵt*}���� }�#��@�c����qE1$
���,���A뎨˜Q�ھ�whw�����yc���w��k���rqyU�U�Ý���䯦��l�da�Ӆ@��h�ϑ���d��Y�����#��N�޽�.�Tv���}��X�u��J�Xl��u40jx�P�B�d8�1(���妖;�1f���ս�ʞw���s vC���a3�\�0���߯+C�,�L0��,�03MS\m��2#�	���d�Uw��cG!b����H���sA�DadTTs��Y"&c!V�c<'+�)��H�f)��[]{���q���Z�m�mψ�Վ4-�Yp�	O>��~ϝ�g<���[s�Ԝ�ݛn�\�H�"������]���s��z�72�,{ub��w��|o���_K�<7��~푱����#��18��RK�;�K��V����_�%�x�.�yqr�UB�d�/z��]ܨ๻�d�����Z���A����
Jz0[��J�쥬�Z�Y�yٜ�6����K��V�dQFԽnQ�?F͐�*+ R�©�sʚϵ[x㺶�Ke��҂Ƶ��<ܶ ������__ː�!]�q[���#H�&~M3|�Ϡ�="�y�E=���f���LO$=ot�*��Η�Qi���J}
p`�qY�_t��e�{܋��k��]w�,;R��E���WV2昄A�R;��7�U�q!���푴c|�����+���O������fbR�~ά[i�bVf��RpD,��\�	��YS�y�փ�0�����9��hK�]�Úx�P� �������9w!��v3�I1�G&�
ʹ� ����k��N����z�p�5͎]�L����o�1���۪d;�q��[�}<)ez�>�#,�+�{�e��+WS���o/���v77��>��\�6��r���>��Jiq���8���kE��#Ś�B�A��콯.$!>�����uiH5�u�7��+`6�O��j��?c��^D�k�&s�˸���	1$EI���]Pa(o�g
����od�~����|�����cb��[���f�¹�׹��X��;4C�mv��2��d���ו��0u����W
���F�__�[�Vc�k,�T�e�o�x
9�;�ѽ/L�WL}9��l��T��W{��k�E9/�ego!�Q1ų�;v�;z�Ջ{�j�߮j���r��Ս�0�Ӝw��)}���$�Eá"�o���{ۓs�� �XDF��#@������ֈn�z�h5�3/_z�d�e���
/��
��e�6{:�h}6n���͏�nl��z�N۴0.���̬�Pf;-�.ٽŭ!ɲ֗�Թ�83{���hP{��O*_4�l{z�w{�.���J�Y!TU]j�!�����Wj͝f8�͚v��	���rі�X�ҭ��sl�S�N#af{�<3m�>����)��xI�3�{2�4�5e�ͬF������}�WM��8V@{2]ޜ�x۹�F�͆A�z�9Yi�b���X7��� G�Y�+9�o�rú5�����"B��2��\�A���v﹐#��3qW���R٢�����=�O�mc5�NB6�	��Z�������1Ӝ�M�ӕ��\ui�?�MQ��"ٵW�U��*U\����w�X���]t�U��Ҍ�1��lΩ�����gA\(���x��enLŝ��wd��c�;���Rm��ftmCEL	M��aK�n�}���ԱE5˥t������h��W[�[�l�Sz�;�Cy���k�Ħmk��.�>���#
�r�ݬs�V����ߴs_��e�>�y	��^�X��>��7ڋBy�3�q7q@c���VqWg�<���fzo�]����'��P���U��/X�zc{|~���[�W՗8oԘّ�.=��*�9�>rH��%�GmV�c�����w఍cϜpO<�U���Y�c�ڦ�=�Gr2G��]ׯ���L{�g]*��eF���^uV�<Q��t;�xm�*`�:]�s{��or5H6��hb��0\[��e��Hmg�q>]g���ݥnl�خ��J6���a�Cv|Ť���o2U}���^^5b���u���/�:E����W����L�J���'�g��~���TDm���TA�b��BRp���qg�vF#8�TX��c�6%�aœ���`�'{��`��`�����;�zE�+�Ϟ�>��\���]�R'm!��� 0�
�"��~������كN.�{o���,���]?QP��{���[�}���7C�^����v�X��H<���$`��� 2M�������¯��EC�u&6s�+ڈ�b���Hnޙ��>��*ۆ�X���/�E�k? D1si���)��7A�u�ɐ��Z�u�{Q�����Y̎�\cM��uC%�$�96�����`^]�pQ�ŻK4����s�7��+�6C#1}w�[�G$p�f�Xy��F�B>O�,[ʏ�B>�a�p�>�2�h�>��1�O�L��\�[����$E��n�;��p3*�.:�\yL���J�fNֲ�Ҥ(��A�Rrt]�E���:��{�9����6�a���0�)$j���t��9�L���*��)#���x��F��ϹH�"�=�Q��D.�a��r8j��p{��� H{B�9��>�2�H@؍�[��̯��.h|�o��ʹ�3nY~\g�.Mh��`9S���|�.F�*6����s�Wd�O��B�|î��:���Y�V���(p��!R@�i0L�{�Ew��tȷX����� ���}c�ڱB����޼����Wh�麂gq���l
h(5��^��u��[�jg�!e����Y^������J����'}uQ�rB�)�`|���d�;�Y0��i�>���F�s�����[W��(����*z>OμO������*��x��Ww����|���U�-�{����1��Jé�3��^I0�"E ��P�8�p�E�n�]o��� CQ�k�Ai�U�ᓼ���M�G+��$6"�2��Z�I��c��7����{�:^Kژ�q�ٛW23q̅V?t��q�37Fݚ�{)YF�g�!�m��T�]�c�ǭ�h֝��l����tB��F^Y^ӼF�+��RM�ې�=��4�=�]�9��0=m���v�t<X8-���G��ݪÃ�;c�=j7bal���_8���;�u���/(7��p�ݐr��#���]�u�@�1�����tu������mq��ń;s��v�����J�	MFd���Z����^a<YN.Ӭ�b�U횱�8��n� ��v\��.�HB.C�A�	���P��e����N����c��?��\@b���w���4>>L��T=��o�}]W�Cj�j���|��=8�a�Lrw�����������mmTg��+"u^�qKތ�D7�r����SA5<��>����H�ƅy8{�����GDh��b
�������{����b�#�ܦb���t���3����B��^���
����H������J�/�a�
[�C���^"In	"H�������}�|{��G<�(g�i��B�����ʫm��%����J��Y&م��h��z�N���V��O�q�?���q��5$f@����/��2�:���m�;��qnB�y�U�Hz���5C@��
C��Z��o��g�:������1O�r�������e��r� ���lV^��t'm��|�� LA��yU�Wn�9ƛ6�{[;���WK�A,��~�ou����?!���_�*ňج�����٣>���O�r�cζ╵�q�1�i����v'
�H������kw>��$
Bar4�G!��o�h��ڜ������W��.v�M�3�E�0N�Y��޸��շ���7�3���7,i89��z���Z�]1�8�̔��ٜPWqo�uX�qq��ޝ�C���_l�u�P�Rϻ����)L|�b��T��4(�l�W�]����_�k���Q%I�b2'���`qw+��۱�Nφ(��<��G��b�S�J�m
=Z�%k����U�(����ށ�~Y�z6��[H�HK.C��/���
���.?�'���
��ϯ�CWy�Cޝ�_.����/�@ޒ���yK���j�s�
n������?������TM��p��)&�w~�־�e]�D��"�,�ꀂ����Quފ�L!�O����������&��ѫ� �"����03�����$y�\��PE�e�y��-�{��{g�/i�]��;��xݞ췠fn�{t6۲��
�SZ�e��߬���>���q�9�@2,����TW�3�#?d�
��W_�Q���4�����k�_P}��0��032����zO�jj�[k�Y%�^x�����nB��"pWr���<�#-��t��L�_�M��=}�]b}9��Ta|���Z��7����sOƪ�ő-��K8�?Bǣi��i��%�j��o���{�s� s���	�U�|`w~?2#��;��b5��w!����L}���q^����ii�6���1���Z�ozP��Bi�Q�xT-���`����4�`��6���aC�z����U��t<u�?>��Do�_��v��Γ6�{>|��S2�L#aD�p���g�	�9_zo��q�U�3������DJ�zX���6�<��]Q
�W�+OtC��1=8�-򣕓w���z{��R�>�����[	U���I^������.|���yޚ�毟Zp���W��</��r,��`O+���/~s��p+v�s�(F3W�s9uo�Mt����	%9�W��;�����y��e���Q�������-�cR�U����,���9S�7~w~��ݕ��~���������OӞ^��X':"��K��R){�k�F�O);��30��@��e��޸�|~G9t�����~k��IUhCtv��ޚ�h���(I-{��63�x��k��'A�����Lꮔq}O]�uUO��-�-^��b���CEӅ%빅H�ANK~b�m)��'�?*�Gm���ڭpᵙ�EQ������Dr���ߟ����+�+�R��~���D[x3�6r�{�kW�oSޛ���D�>qKD��B�:%AS1����o���ة��ݠMom���dt
����:��̸�Wͺ��z}��}��}�J_q5˝o��V�hs��У�;Viㆴ�0o"�iB
��2��Y�$�y�P��&��,+���"P�V�ep�Ԗ���r��,i"�$�-�K��k���A�p���ow*�<�/t��T�(q�p�z~�b���_w/����U�q�vm����kxs6}�_?{gi��0�B�#��/D+7�P��?X�|U�.������^Ư\��m��r�=w%��qv�r��9u�c�����Z09ĕ9�4w����V@('��'��}#���v`��/��������}O�+`k�:���",��O�\��Vnu!�ܾ�.�:|�*)S+������^�b��QUk�8�^ͬu�߁xI�y��?cC�@I�x��<���G�=p���!�4���K�,���5&w�*�k2��f%�q�r�Y(
����okso���������δ���Gþ��kuC=��3E���{�xzi������#��Ț̟�Y|u�ԍ-��/��l@AB�r8*N�#m�kޓ�Y:'5�l`mn"A"��L�/d�������^��v&�dQm$�ˉ��a�2���u@�����`^�nD"p0ː�b2�ƒ�C�F������g��Fs1ÂE<�QF���P��ҟ!r����2� �VE�0~��z+!����B��}���3D���"�9C�2v�^�"��[5�љ;a[�M����`���㱼�jċøu�!���nẾ��)�s)�o�"nDN6��e�h�	�K���K��e�m�u�q۷[�N��'�*{0K�Mgl�ѱX�>��糸�,��l]ɬ�=p i6p>nM��<[�����݂�ǝ�6�z�Sɻs�=8z��'���V�Q��t��n�ؖ�{��E ��1�m�m]&J�5��yu�	���λ�	��{\��v���n7�~���{��t�&n\�P[��죸�_AK����ɩ��x�5���k�v�5�Srg�p��z;3����0-�\�
�_�~������#�sԹ�nY~�����b�=��[��V{��س@4�i���|��]Kꋷ3�Y���x���������ij:����.��G���.E@`hf!F���p�����s"-H%�}�;\@fU:�)�m���5K��sl�$��Nf����$��(]��t�������>�n����<���9�9nG`�7��;h"��@�4rI���:x�羏[��O����Gv�$���{گ��*�ԇ�{٣����l8�5�*�~M2�M�l9#��8x@���/��K��+�{ �/��y�}�����A?o!����W������n���ɸ�V
�w�����B��7 I��(#܌�I#���jG�~�0�~��đ��(��no��P��q4�H���u^���47��HG�~�b���$���r��[�?Oz�x����P��6��;Z�ݜ�\���������ؚ�Asn��u:ʘ��*vRH9[��%��G�{�� Di>��_������,���?���ң4�׶X��2�&co�?o�_���*'�zWù	��×�d@�9\j���V������K�����c��mTx�z�`�^�ym+��t}Z[�tE���O�ݾ+��[v-0v�2�f6ȼ����X��]]�mrA��c��rbKEm�⢻7�"�D?������׃:��Z�O��}��򯌅��DY5d�Y�z+�,��[��&ml/����Oܝ��|\�$"d(�������̀��(������>��Ֆ��uPRW�~Gۊ�F�}��S���%od|�~�T�y���96�o�>��|[���sѕ�)IL�Ϻ� �����'�hy }����}de�a������������)-�a���C8�u��#Ω��m�C�lޗ�e��#�9ᘀ�|P���l���*���>[i�߻ǥ�Mˇ�!���}dc�6��mf著�Aг�4>J��z��20�2@���~�^8���M��X~��^�Xx��n�r�~���gss{t�U��8�q���hv$��Uqs�lbv��H��5�1r1�SG�y�u|4�$����W�z����~�(�|������.� ��)�O�=�Rt����m}��W����k��K��s�Ϡ�%�9
�:�D��{X��ܝ�����!�>�}�A����ۮh~~���w�uW�4�5|����_���C��.{�쯽��6GÚ+r�5Q��Iڿ���\?|E�|. �������}5A�!��ǂ�6���k=7�6�}��\wMT�j<�HAc\9V���s;�f���?GegVL���tA,Ym�B��f���J���xS£ޭٷט�M�7#nM�/W�Y��>��o��	~�3 g�o'���Z�i�@��iz�֊1ϔ�����"���g!�y�Ӟ�"�?Mt�P|@�!�,�?{E�_I q�V!������@Yt�?@�XVu\��k�n��k�����EƮ���SBPb3��`p�"� 5�?��j���߽`YoG���0��f݅w=�{j����J�H3�z; K����8@�!������_{�y�����Zilr�[ebų��'���vn�n�vě)�\��М;AOBv�B�$\8����w�C�� ,���Nz]��+:��1 =��U�:������^��E,7�����h}��,�7kފ��G����p]�S��j�]E���u���D���k�k#?_MY���ό�ѝ�,�7�/�奈��Fs·�Gר U=�}�=(P�?
?��?}��U�՝�'����i�	$���Y�N�����ޟ/�����r.� #ጯ���?g
�a��oW�� yOy���k��K8#����>��7����V��>���I#�b
�禀�O�:�����?^�#�J��Bۑ��4��Pd���;����HN>�����y3��@r����L��O���0��;� �wڍi���
,��� 3��k�ek�����W���!��q�le%�S���h��.����R�[�Ն6yV2�;�8���5��65lx���]t���}� ͮ����P�� i�u 0����nI)�dR�7��=�}iq���ﾓ�̏i����8o�~ ����_�������C����@�>�_g��]?E������@a�
#�d���_~� �@���>�)���3Y�F�6y7Y�x�^��tb�ŋ)�qs�}s�x�mh�uu��ka�<�v]0�8�e��|��a p 
�����=���$}�F�8/�+�}���qk����N/��0bG�*Oy��]E�}Rƿ)ssX��<��N������~���?�b�_W�?��\���׃����vY��d���rG�G��4��_�<�w�5�?����g���� ������W�.p����_�����gX���̽��.����jA��v�{�U��ﲲ���~5���ė�~�M�~V�]�$��V����5q|~��
��U{ξudg�8Q�Xǿ,�֊Q�	��l�}�பo�N�� Y��?� �����li!�6���g�0���C"A&�1�?d{�X�?0��g&��hY�=}){��*�t/�K��>�E���^;5��r됝��x���B���^F�17�G�f�b# �ɫ�զ~��&~>�]rѝ:����AA�˺��{�:�:�w&�C����lm��J@��HJ� ~*R�)�J@�R�?U)~��T"�IU*R� v�H5)RH���)�R�:Ԥ�)�J@�R�;Ԥ�)z���1AY&SY��� exY�pP��3'� b�|rT   �  � ;�#B� ( 
�  @  � M�  jDJ5�@ ��O�                                      |�      � }��v�Ǎ�=juy�x�F+��ot�o=����f[x ��g���E�{�Zޝ�w���vQ<�+�wa�� =�[,�˽�[�绽�B�d�V�+Iw�����k���x �j��^g�������y��
��֦�� .�&�8{��y��Ii��7��7�w��z���Y�Z�E���        =t��;��]�R�Z��G�yۥkDp ���Ƿ�����6�{�n򈇞��N׀ ��F�s^�WZo7vj�eil���Mo9��5�������� �W-�F��x�.�м�{ۦ�;��M{�[� ��{�-绯W��*ov����۸i�Z�B���iC�         ޕ��w���i�˩{y�[��m���H� ��kn�wY
y�sxo]���=m{7yk��K=< �w��x�$u����*е6��k�l�y�l�.���lѫYz� �lPkZ�ɽ,�o]��)�;�3m��;�����Mǀ ���Z��뷫�sb��Qw�����nK2��ݭ��E+-)�P���(ǀ        ��֚4q;��;,Y���x���A��o,Q^ح^w� �(5Ů����E��m�΃���m��y��ٵ�� #���Z�&�{kE7sZ���֍RMݚ/8�ֶ=΋�/ei< ���جq��UݳM��Yvm�6Gl�7e4W���nlV��� �zm��8�d�S68�٦�6��gh���5�׭T��:�J�
���        �����r��.�4S�n�حnX�M��yw�v�٢�� �h�C����b����:�yb��Z����s�lSf�� q�Q{5�7����l/-�I7���՝;��Z�B��м�G�(W�g� �)�(���s��V�� zhQr�Q޷C�hU(Q緀 ��B���a� ��4.XAA����� �"�� J�@ ?bb��P������4�!�Ob�Ri������P�   2hJ�1 <�����m���7���gn�s�c��m��n�uۮ7�m�z�*��ף}t��WjU=�W�U� ��*�\��|��է����m9�|q�M�s�]@I��+'Wc��瀊��{�81��U�#MX�m�Y3��ma�f��r��ͼ"'j�K��Yxǎ0K��w��34�b�1ߌ\5��Z��#h�_tt���۸�#���mo��Q��]�e`xvc�+n6�i{��s�v`��]�ۀ��.��h�Fv�9'�vnW5:��ť���/ ��3� CҞ�vV�=���C��&�_������Ls[wP�9���l�i���2A�ݹD�Yܻ7�o�+~������v�{�D��b�޽0C�(�s�{^���ᛐ��e����;����]�mN����vhoq̸����& ]�=���1�y5�,	��!�{����Y�ӹ��3�uM�n�tm�q�-n��wP������J���52�s�to-���k@�{���rn�i�zq���	Ǖ&����.�&�8�,�_,[U�~WN�9�]���/z�����3�*��c�!���k���voi�*S��L�L�s�x����qgefT5�w��C�s%�J��%�ڎ��F�ǡ�I�Ћ/V�H9a��u0�E��T�(@Н��ꆳ�d���%鴧��*I�xt�E��9fLW7��os��h�P6�[�Mg���}4���k[Ĕ�Ÿ���cl��bE�gj��L�������W5۽��חl\[����9�vt}�en�Z9)C6�H\�ͳw�
����}xƴ���psá]Q&�܍�鸺3��0-���2n��0�P5��l���W_�[\5��ݠѷCm�qm�;ۺq���=&�X`��#XCQ�������_jN�tF>��= ^�^��LC �Lrٺ&���ؐ��90�w��
T��3R�P�#L���g�@2��Q[J��_��Y���D�T�M��}�a���'�6�T�Y�FȲH��zs��smt�W
{p�0ڲ�_��Y_%o8"��6��M�<�Z�v%���d6��ӟN�0%3�xR�M����.s���-=�L �Ħ����:�sy5-��;A�9��{�ђq��+�̪zE�Q�m�=�y��f��]�LCAB����x�V����i�}������Zo08��Q�q�#P��Κ7 ܪ�-ֶ~#w[��z@�Ks7K���v��9�Էb�k#�F60I���αW���
{��٫�o��n�[���ة���L�u!FT¯.E�.w�ۥ����D���
�Y�9=~~�UB�νU�F����mpk�n��J4[���u��O(�da���?>a��(�c˖<�3��l͘s��{j���3�.�'(г ��&��p��0�Ga��8�d�FU$[Ǿ�;NG}�Q��۱�㓉�*JaKpwj��>:t�A˔Q�MI��+���V��8gp5l�h�;�eO
�pD���
ŏ���Y0pyZ��Δ�Fp<��=��w6%�9 ;�n��؅[�'܈�Kr���:f7ps����۶˅�	���/�6l��%���w���@�Wf�o" �v�����v���i5��Of�Ǣ��ŷH�ֶ����HMbvA����{vGϙ;�����&=!��e���F���c�Vԍ���֡}{�ĳ��Ñ���Y�s�=7�'4-�h@ᩜ�2�6�����\}�y��1ۇL��mG���%�5t6��^uE�qc��44��U��<��sAz���K��&��F=)�[�xY�Ф9D�n."�q���tkr��U���h�2ecNj-
��D��se�Q53�@*H�x`���͑�j���go:f�^�t[v�B:�ifZs��r�<��Zuo@�\�c}������PLBsá�S4iEod�^����@9�;�if._�w�:�4���k�맦�xF�Q-��3�(d�j�*9�t��M��Y�͞�C�͝�uET�j\�x�q=�v�KyI���pN�a���\g<�w*�J��&RQ2�5,4pR�@�-��WN-B�����H��5��:�X�9vO�~���P��[=�ޖN�����ߖ
y#��x�jr���J��l��S�nO8��1Vm.��F���zu��x���TO]��O��JX��_gr��G/Wb4��#�ҵ�Yv�A�6��vjx^R���9��o��ќ=#ϡ�޷R@f2�kY�p˦��}U�#h�r����՛���W������+�]0b
�"��vj�M��{��vh��^��Ф�i5�/�:<�;��3�T���ܞ扳��٬�m� +�V@�b� ԗd;��ޡKQ.ک�]Ѯ+-���	�Z��a\�`��[K��K��1�if�xbx�~Nëa��b㴮)J-;�[�M̈t N�i��T>��3���SIVJ���Ft��P囓;��;l�cPA�j�Շ�廁��V*����%�zU@*@sq!�zn\pE�1�p�I2��k/*K�a����{�ވ��t��»�/M��*�`?q�6����j�����k�γ*K�f�+�d�׆���F!����6�tӵ�݈�yJ���p���W#�V�4M=��� 4�K��GWm#*QP�Ӭ�v���kݛ��Ȩ���i
��7Pb�K�T�������x��Ke�,tH2��"�N�L��1�r���~Zڍ�q�2��L�ǓI�)�]bȱ�����^����6�d����䜊Wx�Lvn3vM7tͼ�:J��~��]/P0�M�95l�����	��}�����9�2n0� :���ofo-�
1�u��?(���.B����e����,�&���qԒ:@o.#�).�5SvY�`�f�%�m\���6:�ǜ�D@��sg&�u'�z��9��L>%�����tf�9��\ǩ#cc�ͱ� &]ʺ.s��/=p��T���M��r��	`�T�7�4GI::ҽ���csH�D?2p��A�� � *>]v�m�����}���zNz1��+9 B��H�f��r^�ro$�&�c�qh���w��X��n��@�&;��Y,�dAq��k�y�gv�'�u��:$��s�	�e� ��s|�;�q�&�:x5:�wN���!7x�v�s����^��^��o.�7�m��N'c8�ta��`�쏊�Śͻ"���]=7:),��dOF�6+�oiq����ٹ+�{n%�өgIŧ޷Qjjw5w�ŴZ,뒃��";���
91�m�f�cJ]��a��_f��]{�xu�s�
X��.��
�g� ����3D)���+���_
l� �Q��X;�5�!�{%ݍc��Ldn��u�{5�9�!�8��2��X�gd�'#\5o%
�e�.\�ק47�oeu	���2�;�E#<�}u\F������ Ik*W{s�$ˉL�5��)5'�-75I͢�����'A�Ϭ��9���cѣ�$�8�PPE,Sٝ7��{z������i���xݗ��]ݫC�ef�:�+#η
.�4��vsv'ԡ��Z�ݍ�8��y����T��w��Xۛ�X��Tx����v�D5'۝���1��3B�]ۼ�tɺuQ�ٽ��:���xp����B;l�"�Y%c�}�D~@^}�p&���Gt��\o�{������R��ۚw	�	Q��9i�.�C����U\��&<��ns�G\XI�P$�����"�H|�Jt�6�*������D�16��%��>GP\�&{�H4��ݎ[K�7�O��fM�ʰ�7zsƃ�F�	g�e��ª�U�;�x2a�d�^�#x�Pl�p�r+�7˘�X7)s"�����S��nD0�����Cε���A�7pyg/����=�9e���M�Q�M{�!�Uw9%���;��`לӲ�rf��q�r]ܵ�z]{O��is��!��CR6����ġ�2/m{�l�7yq/.����}n�Ʒ4[{�t�S��T��8b�l�l�_���{8�Y�ü{,7���l��M��%��;�[���.M]dm�Y�d�3f�	E�7�r�5��j�4��=�?=i��X���W�׫.{�K�Ӱe���{��UFu6h�2d�1��u��ӛ���Q�U8'�J���&����ɝ��\��ڸX�����U����\&����X���{�	����%�S���_�Ь����R���n#��P�����M����gK���g\���f�\�?í �*F���@4>mW���z������eL��xC�F��֡��Bѹ���I����'f�"�Jq�<�Qk�B�4�p�6���;Oc��\�c3�����=�w���)�H֨Ut��2�ܺS�r��+�mF2��F�K3�Ki�3�"֋wC5oQE�-�7��ӡ��5�2^�[������4�4L	��'d��+I��M�=6�������|��Oݥ^5'5��:��4;���et\b�E�wf��pPГ�E��q�78�r�6�G��me�����"k՗#��Q��ƨYN��_�Bܸ4��ٻ�6�#$�'c`� �;_W��Dѝ��p|Q�4��a�hR�0V�$Кq�{1U�n��fֲ���B���"�b�(3d\w ۽�ʞ6�!B�v,�^<����ǌ͓��dȪ��9�~�8����a�F�"v1hC8.�٠S���Sr~�h�f�xv��Δ����ó�DjNu��_-ؘ�s�.��`uz;�JI��%����с��a�9Q���2��\0�"�2��*�C�[�)�b��S0\�L6�^ڣY�mS�jf�����'���7�o 72@��ѹ�T�%V�������U�^^�pv�I�(��I��<O}�G0T��/5���3�Ď�����j1��㨍U�Nf��C,K�����1�)_�&"o����0��,�5s��ʪhy{�;�ӷ�y=�'2Z��ђ�������黗���<��r��D��C�h�ǋ������h*
�i���;5wn�b��ͅ�S�l��w���%�;y���K��.�G{�m{^�d#��f$i����G��y�-$U��ì외�I�$djv�0o.��f��s�X
[�Y�f�2�(��w7��k;wm�'u�_ɳ���M�exb�z2�8�q@��7j�j)�t�V�:�NM�����S��`��r�t΀�,7�ܺ���Q�!Y��0:w*�����Ӓ(c��mr� �V� A� ������Wb���ELl�������]L��`���B8��Q�x{�4�X\�:�Ò`֠��w���1w>�&��@H�ē��W̿��;4Y�!�t#vU^��1Ր���{�Cz�gw� lQ5�5��o�Z+0�:4Rc|5��	=��X����_�����7������I���j*:�@5��qO�vz�I���頺�V9Q�{��#����t����a�`��f=��Y���x��%$��t~%�fWWn�F ���H�`wR�=+9����7{��LȨ�ܹ�ì�O%�FcS�8�ʙ���{gw����l�%��I�E�#5�<�������rb�n������b�z�FY�|��/�h����_��o0�c�����*�#����wl�۝ȞxA�3'8�E�ē#80۝��:ʸI%r}��va����=���8l��n�M�"=�d��m�Ǉ��<�׆�UWe_7nÃCp�2!]8k"Q�'��,������R�i�������צ)���v��OC29�ū6�P��C��l�;WZ4l�^��{������� �I�`� nt#�D��)V9�]���ə�J{�E�:S��y�:L������܃\9+<�>~��϶m���u�@3���7�:�=���~O��G��wwPf�#�4-d���c�yI���e���-�q/:��vn���u��ms��qq�$��p��H����(�1�Ċ�V�Ǣ��yՁ���Q���D[���h�.*vN^��iX3{M:v��+-�dZףz�$Z7���I�]��������n�:��i��~cP�	�v��5��4�6x�Z^m���N�4D���78Ď�3k`= ��˭%�1eڶ��o�����VS:J% B����V�t,��M�A����F�-�G�B����-n�Q�ng��H�����f9��OǆuW��2�[-x)ѡjʐy���!:tf�#�&��r]��q(ڔ]�Y��:� �˯&�O����ܤJq�k��Ϩ��Q���4���s@����.l;��w���&�c	�/$Ǽ�)�D�78Ը-�Gv����`y&Nw�a��Cʧ��ٮHvI�������u�;-z�G��s���d�_Q������_+Ɲ�7s�X���D�A����d5��EX�ۀ棨�Ŝ��{��7�+�\��O�J��A�t��]��B���Et:S�4u��:����	�ص�tj�.=��f4W�rtz��!(-��e���]S23���F��¨r�|����r4���:�-�4>yO\ӥǊ�jj2ק�F��R"�9Fw@3����\�S4G�r�jl�Q���r��q����c{�u�1��ѫNx�"����V1��{4������������࿜{�xs��2�1��]��;��[���7n�1÷uݳ��b}�N�nu�-]p�:��oRI�Olǝf����i̥�A����3�v��<����ۍ�ِܝ��t �N��%bLpnʘ�JA{��z�G[d��� ��,;���i�M�,(Գ�y�T��7�q���`ݝ �XL{�1��·�X]�Y�I��*ɣ�� ���&�9
RTtt�pm���f�
C��=we�ŗ���p�.�Zp�G|O=��~?���O$�ڍMu!/*ur�()�\��)YeCb��r��j��u@ �>v���JS��ݨ	vW��l��UUJ����@]M�w�������Z�ڪ���U��Z��&ڸs�+�uU�vF���U\�J�u)<�m�y&K�}���P
�R�ljOpQ�UO\k���n�A�me�^�WJή��,���-�	����L��Jm����e�;�]e� �8˴�F�:��Շ�C[��u����&�nV��]�����
�ي��ێ�^܅v��9Ϙ؎xx���ۇ[S=s�@�ݞ�f�ݺ��a�^�	r��!���9��9g��R��Ku�=�;9M]�ծ^֝�1i�k�w��]���=��ݍ�s`PݸĜq����=��hǒ��է���9e�Sv݌���v�EV���m��zGT�)���Ͷᓶ��|6;*�se�K����GOAq���zL�Gt���l��{&��m�N�2�=�h���7�q���q�unǎw\�Η[sG�<����mҝ��&ݺ���;���m|O_-�j�q\��F��<X��;��������ݑ+m�cnCth�\����. �q��㌞S������\$��,�[���m)+:���m<� ��k��Nq'lS�}K��n������QvHܶ��������(���C+)uظ:{�XݸK����Q��Ju����=�xT�k�W�4얁ѻv��xqn|�n9`s�S�W���m����D����{v�v�ڲVӑ��'n[��zn�g[�Ggr=g;g�x����ymW�uyx�GGK�k�9�9ɞ؊����-��)�]v[��l�3'X3p=��6���Շ��n2/���M&����lt���b�U��ٝy�͙;�{Q�b�T��ۘ�7��s��^�g��v[��7l�0Z:�v���}���=���x]��vA���R�t��������"������7G[e�]#�ٴps��h�b&a݉3ƺzz������v��h9�������-�b���Ӟ��q�ϾM}��㄂7=�����u9�-#��j���kض��d2��^M�=]�������7Y�۵�y7Iݜ,cc>������ݎn����ci�Dnr�g�6�n}.����Ǳ�-�!E����R�lY�(�9��	]ְ�FbMѹ���v1�n1�U^���m�arh�B!J���p�O��lE&��������s%Ʒn�[Y燞{��7uǈ��Ȗ�������z�r�O.�7@��km��!��=mҧs�v콧��j�R�l��ҝ��^8;^�u�t]WZ����r�Y�<��ë^r���Ѯ��~���m�uR�N����<�$��֝�/���s���ǘץ��W�/[qV9yx����[tg�x}�#���Ϭ�]!��V;d�ێ۫�������-��%$���Z�l��ݜ��VY��]��un���͸�]d-�쑻�{]��N�u�s�lGKƖ@��Gtq�j�x[Ջ���ۏ���{G:�&��:D�k�`�xr�X���f���4���q�ޔ���m��������3�sv�V�öȕ��1=fwOˈlLy��K9��M���6�x�v�m��l�n_#��7o�|�<}���hŢ�����p�6�hܘ#�=eGn:ol
�/s�gd�V��!�����r�u���mׇW]q�o7!t����cn^�n1�^]&����w6݄�ܲ���_ip��k]p�lvyv.��lrXx��������rtsӹ�tl����F6�nU];v���Ămt�06�k<R	�vn;8�^��۱�<I�Ǭ��j�3l�yk=�!4.�nݬ������s�	�:3rF��f�2�-�E����gnk�m��>�s,�.zs��'s����� 6�:S�]��9c�����C1��.; �&֬�"6����Yh�X�^n�]a�"��ы�L��Sv�8u��N֪��8የH��#�Y�����v랳[`�g�7]�]�='�+rc
^�]X��uF���8b�v计���_}�v��cT�Y�s�c�2z#]mڗ��r��k;�؁���Vz�%��#��8���(q���l��t[2c[lȧn�x�w[�������\t>{��9���E���+}�����kUT�N����ֹ�S���]��9�~�����sӡS����,
rގ'f��p��y;;�[z�Éż�I8���5g�1����c���z������v�������\&���'��uHE[�!�ۥ��Ss���Lb�#R��n���^��L��X�<b�щn�uv:���Ɠ���,o�.:�[v�nλit˳�xܷF'Znc�F�ܾj�j��n�rQۤ��&��i6����[s�u2S�ɬ�=���OMd緫aن\n^1�^C�t��r[>����ݻy�k����uv3����S�u���qRm��9������m��tە�ș�݈ۘ��.�l�N�vWv����-�lq��r�ӌu]������vm�qn�v���5����&�+e�N�k����xF��Ƶö�W��o3��.�Kf9�͍��۰=� Ŷ9�ϣ���&^v�ǹ=��M�v��Ŵ�^�]���@9�7m˸x��CqP�7m�V��k�Xŗ�[�7bnd:W8뷶�l�m�r�x�ڶ}1����a�����S�W�]��=!��u��gE����|v8N��A�{#��Ǝ{g|��=�Ks����e���a8�!�gf� ^�=+ȶ�uq�%/=un]��1���� ��ƴ��z01�s��:��K�Xݷ��N��S�<�&�5����m�l�i���-e'Wn���]��5�U�^ӻ#�Z�ݞ�n�u�nz�9�g]�s���pe۶�uRT޽��;��ez��ۍvçt��f܂z��񳁪����۷Hkvv�3�!���ͮ6�݅�:�Sq�6;3n�J�n��K�����4��IsWe�=B�9�wH#�Vr=��Rrmn�y�mt�Q���yd�Yȅ�� &��{�1&WvႇR]����N�zqðv`�ӷ��ۋ`Gj�q����Ńe �{G�tz����n��x��n��
x�֔��c��G\�s�a9�%�����р���mV�{'=j9�sq�0c�x5�#�2�M�x*m�5���d��wB�f<䛯v�x�=�\��E;ͫwm�cwl�cY=' k�n�p��:��(�_Fj.�i�:�c���;�k/&�n�y�s�|XM�8�;v2�N�s���*������>ܼH�=��q�"7 ݥ�(���7n6��k�A����c���6�sa^ܳ���Ӟ;c"ct�z���=�����NN�u�`���n�+���F(������1�7�7nN�O�b�c�7OV(�!��q�tl�{E��Q���]�㑎u�nn5Ȣ�`��yؒ��9nnA��ap8���z�F�M���^+Gkpm��7k�@j]裎��#k���ݛ�������}�/��5�N]�Е;��۴v��m�]��kb��q�>z���ָ5����.�v]����g���GX�n���;Q�-3��&��y�V]�{Iؼ}�;k��v¸V'n�"v2�g�s0v�`��x.z�1��ls帎A�u�c>h�۞��=v�[xq�yc[���)*ٕL�[��k�b8���x��l@s��ݮ���9)vv���ˊ���c�wo,�l������D&7;�-��v|än;�/��,s�Z]�1�s���r����ݮ.z���혘���x�5���krf�u���1�NrNtj�ܹ��
nx;�0m���z3oRD��r�	�<������lu��tLd��]pثۄϧo ��]��0l�a��/�֎յ�7W=�<��4�7�ۆ�gr˸�6�o	�k����v�ݷrcf9�@�NK����������F����!0g�=]T����{����n�۵���qC������i�f��M�t=���99^l`�� L?���7|��a�CY��Ok���=g�cߊ���콽�qC\�T+X��ض%n]p[v��q<A�۵�����+����`s��la1��N�K�笴m<m!�,�;�H����X-���^c2!q<��m��̭ۭ�����)�Z狞�^vm����vpn����sp�J��x�m�z���fn.yb���N����z��z1c� h�a��M� :;jvk�:�8F6��׷��kbδ�u]&�z�V)5,�;oi�n�`/-��IÓ��;rv�;�{lv�8wbJ��k[\8��p	�Q�Y�x�K'.�d��\����STh��7=��	t����m÷��Wp[�a�mn�s9ĳA�ˣ�ۨ�S��p �7������Y~[O"�7z��ϭ�ے6ƓG="�<q�g�s���S &�vz���q,a7E���뒰��r�ٴR��8۰<��ٮ����M��&���Ze���ַ>˨�buxGh9xۮ��9:�'�B(�O\qp�<�m���m�<e��K��B�e�2l��o3�9�[vW�ps�p�.Ƹӌ���'dc�����naQ����X�ݘK��Xݶ�öL�m�j���-���;X�*j�Lf�읆��x\]���1p��h�v's=��"m�]DbJ]+Z
��Y��v�-�ۃ��k��9�l<��ͽg�x��oF1���G[<1�'mj��ƹ��_V+fB�8g���d�ط9s秃n�z.�Us�=��1��N��R���r"�c�o!�F���Xx�FU�F\�c��#n2�kn8���]qė^���Yn^����q�!�;0&v��^{��h�u�g�tq��pOn���v��Hv�oct�w2�r��[u��9v:M�{u۫t�@2ӄx�pNNѲ=�WDj��S��5�����1�uqkmٶ9����+�ܗ���ף��,\�%���ms��7]���-�풧u<m���ٮ�j��y�v�t�'�[ɮ�)V˷�����u�5��Xݣ\�$LW#�Z��&�u^�'&�ݞn�PكK��Mn7#:0���vã��]�/gm�n>�u��\��'!�h���^�U?�j��U�UO���^)^y�N���m��m��dq�lX�v�;n*Jc�jhUs{d�z������Ǉ����6�ں�6�+�0����݌�z|�g��1q9r@���vޚ�ʹ��<��\9�J�s�Y����m��
+����t�,�:�ڐ���ll��6�۞ѣ^�;�j����q�]�`�>6W�q��k���W"<����qqu��PN��.���+;��{cu�n�pz9�N��ێW�Mv����s9�
y������k�Κ۞��qr[���=��ph�A�!�f�P�I�\L��mz3��=\�n��d�V�Y�p�'������������n�������Y��>��a�W&G����>!���v��p�:w���S����0VV��c���ٸ���c�y8:��:���Ƒl��K��]سcG�U�Z��^A�[��#u�Kw\�S�tn���[�FӢ��Ys�`��{`��Ls���,�<%o#\l:����h���{8㑛ۗ�e�P�e�n��3��H���M���g�Mt��q][�vv�����/U�U��q��V����9y]pv�n:�b�.��]��������xN�k]t�v��y���oG6ݞ��l�x�6�lSt1������:� -�v��*b����x��:�n�(s���]K�F�S9�|9�E�s��\WeGAgrt���;��N�x��<��q6pS��5�m85Ŧv�8[�v�"[��ӳ�q�u{s�`�<-�Y��nb#�s�ݡ�U��n���Ov�<8���V�M�9K] �ɴ!{7�C����\!�Z��Y��<n=#v�F�səI�����Mt3�3�8�[L&�M֦�GE�L�.f�v m����t�l���&�K�ۮx'F@㋃mY{8�sgYM=ە�mZ�;	]��kv7)n[�s������m!��\�@ݨ���]n+���^Z08��<Y�������m�=/W��{N�8���5ݍНDK�ǋ��X�݈;A��s�۞_n�u)˭����-�2%�����-I*� ��"* EQ?��nyzm^��\��c�g�m��O#FY��LN�;�\;ps�n�F;�a�T�yC���.�+�k@mݚ՞���ޝ:R���]�n��cְ�G;�b���ײ�N�V�v��s����He�N��Ü&�1��X��d�^v{[Rh�k&H�ύn�S�7	�ض+-��xe{G�u�N;v9l�pcC�d��}���N읞C��܂��^����0�]�>2n�Ʌ��{r��rWc�� ���~��>~ǝ���R��Ѽq�_k�>F#���^�.��O�-�e�����S��U],-`�^k<�
�U�E��cҽ ��������?`���1-{�׉���f�Y�7.�����Ee� s�u[�>U��T`y0�gWT�TA\�i�E���r"������0�����roX�a�����#�	U`--��T{�О�T6������ߦu��{Z�\׼�0^�yhP]�5V�є�\s��Jю�޺Ne�:���3!�(�M��v��}ʸ���ާ���g)y�EV��Q�%m�b�>�p�5��4�;]���nyM����Y�v`�;\n�v��e�����U۴�����c�,>��Łt�}Fa��M`��*q��W51�5^i�6{��Q�2C97 ���0�HU5e���h��d-�GY�,�}8p���e�ߦ:/nY�8������xx��\���4)˳�����j�M	�2q��BX
m��P\��7bٸ{�����1�Cv$�D�)�|�_
_՛[+2mw��ɑI-�!G �o.�k޵SvGd��O�}n,Ш�B{���	,!�^�U���ki��%�I�n�$�(�qb���� ևJ��m��h�9�����ϼ��#M�X�Zr}��Y�ߜ��2��d,L�(�(��N����v~gi����/�x�P����ǁ��b�bӚ�u{�oƳ��Æ-��K��od�?U��	�`;P+ �e�Ĭqa�xܯmhm��ۭ�Tu�x�8�Y 	#��7$�0�BF*&���^�!��ܱWݒ��S]R��1k���˨۽g���۟V��l�ѭJ��f��D�0�%92�M�3Lv+ۘ��h�x���/#1[��.�G5nд�ϙ����k���B2Z�u��}Б-Zr��hJH��}�M/Ϧ���w7�.�=���y�CA<"��|���=k��^Ƣ���n�1���w�+���*�Xp�Ʒx�Ȃ#�\��ʷy�L�+:��׆rո/�����X2��U�c���#$')̄�r�,���+
�v w���Ią�0��=�.m"TX��1Y#&�j������v��2�jג��JIA�AbXM��h�Gr싮5��iL!�;��d;l
n�u�T3��i.\��E�J�s�ϭ����VDG$tE�vGJ��]9r۟;��^K]���v`��˨��1[�|�sQ�u7P�b 5�I�^H�~�nk�3�/��Ot�������[�ܱ
w6}Aޓ�*�x�![KFd1,��cvd�ޥ��/�)ضgɐ����A��Ҏ=���Xb�wY����wp}
�����zwm��V�ve�,	��P���͔�{����j����#��/�q�u�^k�1������V#�a����R���vj
���_���]��5�ϔ��ܛ�7�}����]!{�nm��t��QT���Ε}x{���@k�d+s�5x���Ǟ	=g���%�횰x��]����e�ҠިI�������s0=�[��5���A5k+����]�(7a�TF��#	-�H�z�c����g�Ǚ��=���X�ˁ�r+��F���Z[e�r�Qi�m��<�q�r=y�:�7�������s\�ŲP@	
�߳y�U�)�����쳹6���_�e���s#+Y�ѱ�<�5w=��i�(T6RKw��1��u�k�̼��<��/s�7k�ҡW�>�e!P8eO�e�����Cx�7ͦ�7���b�� ލ=��ϸ(Y�^Sv76�vW����NX���<8X�i�wwa���С��IE		�������d��+���\������1x>���c�U�l1��B��x�wG�iF�T��Ո�I��he�b���x_���Qrk7mm���d-l ��s����/g��l��p}��%ncc��p��3����~ �b�,�&��G�P͑�)�����Yl��cI��I,�-�R��eD��ʞ�4��?ޛ��8; x�qͲy�NJ|�Y�Z��9y�f�	�Qg�n��ܽ�τq{%Okc��뱽�vw�Jrk���=-�Z�=���tp���0r�Ͳ��*�M�쩳T��k�c��/F��Y���J��0�/8�p�V��z�D�_�x�wb�7\��=�5u���d��Ӟ��O5���x���M���d�e12v���nJ��5����7���Co>��q��z�u�.Jm�^��܊+Vw�Lv�٭�&$^S�FǇ���![������z�נ󱊐���x.ؾ���g�2�C���,�gmg�����o��bN�K5�6Woc��O����Py��ɍy߾�=�HnT��G-��$yCn7H����bVnԌ�BaHa6ܟ=����{W�/%�]�������Ǵ�C�owR�)�e]�\싻1w7� >D)BIH.qyk��[���1�����b�/�p���zP�;p��G�}�i�ħ�6���r#9��Y�z�X6J���V!����2+�����5q]��.so�wN����qe��d���)m����xl��p��r����n�x��
�m��j;5�k'�0AW�뮁h!y���Tɘ뮢2�E��>�Ͱ�4����C�ç�]���{�+�Q�;��<[?L�$��n��7
�)�1[�ݻ��q_�/3r�b֚�\d7<Ff���X͛yf�o�	����\��1�6v�/�^�FD���{�#�#s�l���?@m�F^5{�f����Ӿ�f?���3�|�_d���0
	�$�7/YѢ�]���s��.��n�JhUH����u��W;��o�>����2��ٿ�hZH�h�|��L�|��ϕ~��A��Ȫ�;(fR̉��Ԏ"5r���8ci�'U��3)HRT�D��&%�X����ث�Z���b�v���e0�ה�J���m�m����\�� ğx�#�Sd0�FS&������v�#�޺ˊ�a�a�Վ��^kn�=� �[����y�zz���xރ�X�pj-��㼶.��Y5���2��NǥoS�������Vh�QА����'�\����J��o��m��N��X��:�w_=���G7ev٘L�'����L����D��IQ�V\���� �6�����ʸ]�t�pc�ܘ�����Z�����0�{Cgk�Foc�'Zԕp�x��G�K�����x��5��{� �!h��4��[�}`�g��}��)�@��yϗ|��t��D���D>p�K�*��}vEPQ�j��VCÄc;��Mɫ�Y���A��w���\3�ܭ`�)�� ���0��\�v]�͔;���94 �j�n9z>/L ɮ��m�=����#1\�i�M�O-�0 t30f�a�n��y/P��������q��\�A�{0�6�uY�d�p�D�%q0c.Qq?���d���]Hd��}��h{(q���]�l_O_(���ַ�ꮙ��X�,��ZnB(���i�̐W۴�� �(0���w�;^�7�lڝ�x�۞�rM�G�"ZЁ0�s<��3�����[K�B+9I/o����7�Y��:���ݝۤ�̟yc2�)�B�E"22�Gk]�P�W��ۜ/�����-�k��ɟ��8{|&m�����E�w\��t0� �
|{�Ǿn�2Bgh��B☗�:�d�g���VD��q�}�}}O�f�����61�������nI�'�v�qn��H��Be�;(�����	� K�P�SGu���d:
f�&8�}pz�A����M�r�K�!2d�2��"�q���6�q՝�vu&&�WMgt��E�2�*�+aQ0*Ո��XB�{�K�q�]��[��a�����c�{�/�p��@ ԑ��}��͙;�ڰ�cH���ޝ3���z��>�P/���<j��ث�K��цb*F�^���p�g��K/�&n�F=�%8r\*JU�z3�õ�r3K�k�J�����?P��f�P�98�WU�+�֮��']�nF+P�� ]����Z�U�������'7O��+�`�Sy��j�$֪�x2�?:�F�[ߙ��s�rQ�)H�Q���6�oK���֏�)܇�"�$��dQ�l���X�Fd�[�5D���:�$jt:u�K����h�&�ގ\��a��*q0�cUi<yc�9c�q�/oMٝAEa"�"�wO�ç|��f>�zR�M�i��ms��Y�m�vy�q����4/Xg��l1�wQ�sf�ۘ�{uOg�[���Ҟ�v��o��ۭ��s��nv�-�z%*u��v���ɪ;α��n�:U��Ȝ������C�8g�k�z�t����E�fz:�};Z���m��eO.X���Z��\�۰����W��g��q�.y�{܈����q�Z�Ņ�x�㱶D���p0��:�kc�뷷-WF1a��ɼX�Ŵm��vD;�6��P0U� �	��������;蹯r<�������3O���LpI�`�[�C����l�*��F� Ę*��w�^kM��3��>|�'��?d���V�n���ԜS�U�i�})��w0�6D ~��o����n	��H�}/z���9��h��W�`���) U�:r��Ml�7��������C�����TZ[�[�3y݄�xG�uq�4vSN���*�-ʽؚAj����f�Bx�WB�N�J�t�6�^q�L���%Ġ�(<�s�^���N��͒��#~x�>��(�/u+�ܤ?^k>�y5e��S�V�B��8Q����l�m�W���&М�nSځ+\v$k�5�E���(��L �6���3<�f�3&�ɺZ��\/^֮�6��틡(��	*��ײkJk>�|�Ԡ�d�ږ'V-�FY�-A��oi�ed8w���.�;z�=��� G��}�O+x�s��ا+��������Y���~�g'[�o��\�썔�Μow{_gp���)���F��,��})�lXouY�r:1X���n����%(9Mo���D�<��0+��,@���l�܉�-�tK�v�o]M�87�9����"Wb)$hs�9���x���T�6�e]tW8SG*7:���z��q�÷oO<\����������OR����Il��	�rwr�ō��p�DF�X��oJٲ���u����;�%[�`��Jzq�U�Q�z�D�Zæ]7	i��[��]{���׻[Z�_�&:���ېADIS�W T%`^��=g����yV�Pq��6��9&.[ֹ���F�c١���JH(�T�̶����]�}��x_e�w���0�S�ys1�����ݎ��E�:�'4Q��!��)�o6��c�#g6.�j�l���̽��\�@#��;���^�S$l�Z�#��`9�u��v�:߰�O��L#�ݎU���Ϯ��5��*��e� N��qo�I]5��_�9�JG�Px���R甘b8���Ӟ=���B}�"��	��64a�M�1�_���.y���t��K� �'��:��Bº���bv��eF�D�c^� �Y�߉;*�s:���!m�ݮ���s��b���d��C�z�VC;��eag���wh<69�/;݅��u˲�{��[t���`-���g�^=:p�.lgy�Op���/��Ƕ0Қ3_p���� i�i�/��Y�ǹ��ڽ������D͋L��@VS�A@�ρ�����<ơ����ډ�G���k���˳�#��|a�kG|��� ��4�QUcf]kD���l���G����J��|(��Yq	{�=�Y����5����[��G"�{�� �>:��Y2��]��b���~[�8ܮB9<�{�^7�����n?3�)Y��7c�(�ݽ�g���kp�۰^�NV�o���������#���[�q'6�p��fЭ�܇6���9Z�$��d�W�evp�qɢgK��N�;.kه+������C��(�z�Za�ޞ�v��(6�5�{�$��g<d����q���Kx��y��{ގ@��S�|4z�f2���˽�p��!�U��;y\$���qgvu��� ͦe�y{�{���.�Izs�S�V�m�2j�:����q/f�nsn�c���l��輸	q�ɱP�R̓���w������

�ӎ���M�l��e����bى����:�Ӯ#�N_��6�]�nՐ;���x��/6cH L"fTJ
fR�ou��W*j��Q����ی���]��?)�Yм��d2w���e�R�9oC��o��Y~�4�-@�Ec�3j�1�w;�#�P��9�:��^��î�z���*
@���9���v3+���{E��iW7Ya�󇷔4J��
�����s1�<Ѿo3�ٞ�*��T
������K�����L��h�����VU�����d���T����yϰ�;���X!�ꢢl
�{����qq��/����ƱL���GMb��U�ջ1_	�����^��_�j��st�ԊFx�>�
�C����#�^��;(Vd���6�Nfk6eq����&���Y�^A������+�G�u�^��U�~��h��Z
[*7B,�Z�6�7��A��pg=�_��땄͹��ݸF�h)i( ��~_U��������ᛤ�}��6m#-��yG�r/�{ܳ�k^��h��0El�;iKm�4�ta�8�3j(�ʛ�=�.�㊥��]U0�Ѹd���+�%!��F;��^,n-�+.�(��Y7:O�у�*wS�?=��ks�w0��=]��uZ���6���u���I����2��ю�V�y�bcݯ}��v�Cc��kX[�c�_p��Rd(R%Fc��U�]�K�������L�{@3��O5�u���}��V��iq�h�@��PC�[�Kt���R��,��׾�>w~����O���ھ��3�罧ޠ�`�]���Ū�E42���*B�(&�IR��S�S;�a;�.�I�T*�[FޭO4�T�J����e��2\�z�>�9<Y��\�g��eղ�^����n��Y���tǲ{�(w������gr�?��� �P-�en�9eN9Խq`n���k;���/0yJ��&n��;��&���v�۷`F��c����,ۭ���E�e�87\wB=���uY��{<��{8�y�v���[���ٰ��M�7�������A��[�;�����Оg=l��n!�G�I��b����5<q���݄��b]J����$>5�=)��vB[��4c�qnz���Sj�K�(�:�l]uD��6�d�A�3����o�6�j�wUue)'@Pd(��#!{g���yvE�%����Ԁ��6�ήĶ���P2>U3~��ݙ��-m�X�ii`(�H���~'�Lt���E���U��
�]�n�^.�gl\h��YԶ8MӕV�V�����S��ou�ڦ'c.�wmY��D��	Uuٙ�m��b0x���5��Eb9��-��;�ZkTh>#d�3O=Rx�!��{##�9��<���k�'S�3���c׻�u�׷�b��4 ��YPVm,l�Y��Gvh@��l��v]�lC����u5���u���;�*���}�mf+w�V(��������E ��f�Y�n�,1e�q�9�R;Z�3)�q�FN�aA �2PD�RJ3C�eH���˞Y�q�̘U���Afvp�`G*ja���?l����� ��Kt�aXD�z����o�h����������.��<�N��|s8g�N��)͍oqF���TlHH�4�4R:��r�xg���E����{n��[�{�����[�J;�&�aW	�r�ck�4���}@���´9�xw�w~���`�����Yk�X�.[�mOT��ηR��c7��Z����
!})$;.�n)/Ç�"��5p3&�Ou)��v�o�̵�v�n�v���V����Z�0J��e������o<}�(�S�H���h��{���޸}��ұ���h��:�������'fWV=����D~�C=���U�>��q�v4�ny{n^2n�ѰI���V�l㛨k���~�+�[��K0*9{��B�t~��P`N���ы��WSV��J�II p�+������3z|�ۖ�����{8�oj���,�o1X�y5#��q�޿rv�:��ݡW�c���	�X��$��-�O��y�����9�!�W(�=�@\#+O�/	>�U����Z�w�����O��}��d��q�m�z�����ޘn��_.&_Ot��윱4Y�W;�3!v��nȰ��]�r��)E�%��޹�.4�t���)���[���W����oZ
�V�yӝvl�y�{����,@�!JB��J*s>/43��+2Wi�]_�OFH��a�]Bs����k��7�~��X��a�)��h�z����F�5��E$]� �v�x�_j�Dnٽp��Mukv�XBZR�Wcr"�@����B�{j�]�t����^<�8>so���;4�NeFׯ"�>�g$wI#!"a2�QH�k�*��|�cuZ�Zd�����X�v�����쾺�fpM��DoP*wmoqyZH�Jp��/f�E�w�/n�n����F6;�l�ݷ�lԄ��1��"���Q�UϚ�1h�`:��M�szL���8Oj��x�����d�Wnfv�[�[�H�n4��`�;=�B�����E�����e��<�ӹs,�}��u�`'c*{�5B��m=��b9���@�@w�tˤ鞢zܮ�l���~t_�L�3t��դ���wCJ[_-��]�̊���U�ةb3��qx�m~?,�����w�L���
���j-�Q���R)`�#* �b�D��jrYBק����{gZ�{��郱�=3ѹE��j�++T��Kc�|��)�>W�S5�=lFL��S��n>@�����!kmgq�||�~�Sj�Wmac �\��l3;�3��n~��3�r⫺�f�G��)Q�G�zj�� ʇ ���W��b�|r��)U7�:ȣ	 Q(jI�_��!�O�w�1׽�G�;S�O�5xm�^P}q�2�'���Ow��.^���,���!���勼�˽�P_h]H�ѭO����T9_\�h��50��y�q�M`���1*
� ��� �E^QT���<��/�+�sK���3dn�0#���J��W��Տջ;c�.׏g�zp7M�
���X���.�iy�G�=#=ޞ�G/m��(x�S�҇�p���:y�W����7��^(<��{wQ�JWs���_;�B
H����HQXM�J��� nfuR���n[����p�gQ�w$5B���)~u�6��T�D�b6��sv��ޅ�z�gc��]P<e豶�Og�/��r�x����!��{V����l��uϷ#�K��q�����;�m�۝�P#�5�=�Cۮ�#�{Y����Ή�&F�ӈ�{X�N�]�9wl�R�]ɻb=-�v�%ׇGN"v38�v:Ǣ�޷k v�M�\�S7h�W�)�4�۰����m#a�J��E���y=�ĥ�ʽs�]��Loe�U�^�K����\�囖�>����r��S�+��$$*�bm��ԞJ�U�qO]gV��Z�9Y��b7�2�#u3x���Μ�kW��κ6�Z�Ք���uHuY"���UC���Ҷ*��1V%��ʰ�2�U�u	8B��R�A^[���Z����}���ڴז�Iυ�	��w����m���ݢK����n��}>��%�`("I)EdVf��s��6o�:3M�`�1���Ef��B:��,*8I��U1]�ʖ�C������q�E�J���ku�خ�ӑ�[�ٸvw&^��H����]r$�m]KaA�L�0�QSIs9[]}[�n��9��j��8���:A;;1�	؍h�Ge�/;-ˣʅ�$��0P2����n��L����_�ʷ����f}�oս޸�����^;��|������`B��h��@���T��˦�gg�#1�r�\&�^�c�4/w��:=�|�ܫ�r���ݕ׷=磷�]԰��7w�kyl%��j�K$
]�[$ݮ�Y�+��6�}f�Z"�r�Z�nf����j�U殮�"� R�B_�)��۬^�]��>����O���cެ�p���7�4Bʍ����n쌻�9T���Ys\&Kr��/㛌��է.u�}�̑��H�C(�X���8��e��<��7���v�{4�=P(V*5"���IZ����A�©ή4�w\��;g���kύ����Bq"��XYpy�R����	ֺU��f��{��3&ـ�8�N�.H�ͥy�/MbHQ��t�Z<�xY������"��o�eQ��U76��ެ�ӱ<�'�[�� A���sg�}�zI�a#!��b��������G�-0�v!���F�nq�"lU� }��qmv�w���pl�9s��i&-Dic'FvR��O���|+]��$ȵY�+�v�NoB9����t��qj=�<��H�# ����0��*߶D��ʳ#q.�=u�nR6���r�S�v/��ª�gG�&%AP��s-�y�rm>��ZV�&k�U��u2������w.�s�>��!���Q�g'����erRT�*Qqݫ����c���Om�f������.��������W=5U݇��pV�)g�bp��4�;Vz��na§8u���;�F}��mXPӄhXP+AH�"�ߔ|=}��#�L.��7~5	꽜2�~�I�}YrV���c�v��p�`��ʮ�j����3i��]��r�dwo�oXs���4�\� ��:�ާ��5��!�o���t,��9-!џ��l`���I�7\��̧n�=y���Mo)�s�,�۾�!�|&���
���L�1{�5�
�t�L#-w	�8'����MKR6��{�HyW��?{d��q}uN���g�0��2BR�S�52vO�[��n`�g3��J��v��- �����<�8Mg�wZ#kn��fn�P�Ї5���
%�S���h��n�ICO�7J\9fUD\Ctr��
>�S�5�jso\b��Uޫc$k��g�V��MUHLU���}��*�l���I�C�[��)��ݡ����Qf���������Z�v(m�x�Wu�2�yN����Vi����X*L܃j �)$) �y<;o��'Oh�Upd�� ���u�t�zA�������ͳT;Ҍ�d�e�H�wҲ�F՟�Tn�Vl'��Q��i������T˽��nn�iZ���Ǻ���S�[En������틽��rn�}rLD�GD�Xܴ]���['�Wբ�\�ʨ��$��6Ң(��7p�k�_T�����Ü�FՋv��vA;�]
��H�����s4��dɵ�w� ���裈�o��Tg�V���nu�l�b�5�;�EMi�[P���YG[��״�8��$�scA%;��)�@ymN�h�4j�cG��}��3��&/��Ӻ�#>��'N�·O��>�;ۖ0 -`hi:WwU@Bvm,��&��5���5���~���3���D�/ۏ�Y:� K�_;.�oz^�{�V-ə�� �%*s��>�`
��p����f��Ǳ>҇j��@TUNoWjUN���gH��&�{u�S��WN�\sxeA9-Oie�5�+N�����v�<u��}@3�y�^���\��=w�ë�<��u)|ǿCܟ���yl6#E�K<'��vh:�����e���_c��ĹŖ�֒7�ڋҦ	��V�qp��7�?x�`����� �]�����E���q��$���j�������=58�9���)	T�����m��a;bv�\���A�+��<(��xP��*����x"��O:�?lb���?�)Of�+�U9��j6s��nX�ןd˛���X�B��+7d���0�;�s�_�޾�7�X�S(�l���nt>��2h�а�C_lZ��d^���!H8��)�(%��Z݄C	~��	��9����c=�lg�m�3l��H���V�D �^gn�nG�� _�;�����:�z����Ƴ*�<�rL�ȄHIH���ܜ
���f��ӷ�\�����bG�˻ ���+�/òr��n3v�mϓ/<�[Y�M�tx�k�ǝd�qj#9�3ë���v#��\֌�s��X{���n�:��Eb7	�W=�Ooص�q���8���ٻֵn�k
u���7����ƻe�S�;�o7
V�oNK9ϲAwn��lkqm���J�qqD�����p�:�dN�ntC�[]n�y�P���9줬>r�uWf��(��K����1qW��ی���v�\��6���W�d�m��:���wa�St�X���x��3�;��nM]�^�����i�;G�u�>�u).��䐺#�m���Ʒ$����e�{]�%��8�0�r^0�j�l놩��6�)�;��D�g���`�˶3m^{
ܸtf7�
��m��A�X;r�ɬ/nc��oE����V��u�yݜ���:8����@Q-�L �\jɮ���A��e���4X�vn�[k���v�����s�Lt��7V<R�l��Vہ��\Џ�w��v/&������Y�z��GK��s���l}�=�<�2�+�6)˳��u��l�z^=�X��良�G[Z�]�q�{m�Lv���cb��\A�b�n�n+{y�
��un㔱,�y��h�iRs���gr�c�p6n6�n�mm����{�Ґ��\��oS�[�kZ����]nOOc�먮���:���������v����q��&p��8d��͑����s���/W6q�bd���qd��*&�.z�F�=����gz������k$�y��m�y#Y��m��>�pu�,/m<x��:����.{R���ov�+�l��d�B����u�/[lr�����e������W�t9��b�m�Lg��|pW"[%�{675���$�0��[.4�a�ݵ»�[�q��u�����4%��d��6�j�J� �a����͹�B�,4�����-ip��Ǟ�cQn�{g��ln��Z��uY{\EdGC�<'nM*S��2����y+n��N��"ݸn.�Z��F9�1KʼCɝMΗ]O[1qpnt�I�"�R�[�l&���]��ms�$�tt�sӯ]�����q��1��n˹\�,�pK��Vnv�(E�pOD�sn;8]�;��d�W��9�p�n��gɏ5Z��aǀ��w9=�v��ca��y�xm����A�	�nk���v�=��Y�0fK����nx��y�w]����2��5�A�8g�l�]��_Mk�	;g����u�wZ�H�3�����厎@��#*R�>�	{��E��س�U71E-[˥dqtև�7���F[&mU�3<U��j�%p�N����j�z{EZr��nDh��xѱ]��Q��n���[�}�W����Z���m���EL"�D*nk,�Z���O�h"2_=5�5�t�8!����C.yi���;�]���]��'Y��V���Y.dF�qA�i
�v�<޴0n+9]S� ��	O������X/_h�ʂ����&x����{��^�zz��Qr���U�`a|+o.S��vt��(�A��6��hD��h@�����;z�7K���n;#�u�ۥ��vp��N�≄���0� =�e�ϳ5˰]/�%��Z���*I%��q�QX)\uT�%@��Q$��)Z���_b� ��oAn�t���UQ0n6������b���cZ��{:��k��(�i u��W���qM����8�ˋ%QF�j½�����Q�1��u�t�� c�܌��nO"	�jZR�ͭ�+���>â�z�a�S'Eƥl֣T�j��`�pV�����-*�:t�=��g�;Mu�9���j���g
ꚰk;n���6�
������VΚ�0�=T�BQ �D�V�g��V���#����n_}F�8�����M(5:�R��B�i�Z�qp�ɽ��~�p�Ն"�+�P�ً����β[k[u�6W����Xi���ⶕ��IX �����+W=�f����Fd��KvVAnUsõ�+(¾��g;���H��*�k�(�����e�p��B6�����*o��;7�+{,,.�U�9f��Ν��L��zo�����#o#E ��'={::�1�ܫ����tF�[TI����x@zCs���^�1^���j�}�1�bG���}��ڶ��*��_?�S��]5v�d��K�l�@ts٪����vp>�v���gR�_a�D������*�'6��x�kGg�7)���U�J�y��l午��dL���!�gyO��|\�����(Ӳ�@-;��z�"�\*˩�E�}��U�c��檮�����9�^�bp'�_�.����L񦃝���(=u�74{%�����b�wA��yN�d{N�g���jwh�5usT����<���i�{�V�v���R�7X���ۋ��zP�A��nBm��xU���7Z�VXܗ�~�-Su���┱�(�x����z��֚\5��'���޷l�n�QUk�k_+��F;Up[��,��&�ds�2�Jls�f� Wt�_���S ���%M�V���v�W-��W=p[�|^&lQhd���T}�&ٹ�<��o��~*
�����g��\�;�NL�7uk��o�/w�j��da��x��� �S�7���b�|w��^ޓ���  �����"���]U�lW4��]5����Yݴ��q8���P��Om�ᘶ[fL�p.�[^��l`l�m��{p�s���5a:�Q�e$�T�H8�PKw���{��+I�oV��fn5����3�`"l�k��F����8�so��:�����JIᬼ�X;�v�$f����yf��G��,t�����u�q�І�[��T���<8��� ��@D�������:��6��i���0��e^c�śb��}�=m;��S'�_�F�AVQڑ���3���X���w:����sV��a/�ș�aÛ�=���f�����Wd(H TJ)�,ҷ_5Y�+uR����'�����5S靬�u֕Cr�\d���@D�s��z=3�"�%���M�q��ڀ�Db-�y�^��fy킼���88W���@���٬{Q��߲����_��ў�v�F挻sv�㌶ݓ�mH�p=�����rg��l��e�=�������j��Z^��kx�N^�;<�[�3��y=[M<�۷n�u�F��6�j�;v�7�;�8D�nxܜܦǀ�w+�^.�a�������nP��SO��b�F��:w��\��q>����N���I��ҁ�٬<v�$S�n�\�6���b%��O$�g�ȾI�q�5۔��H�ͬ��kW|?z���]9&���&
��Q*=�wIc���Y��Ѫ����v7�Zb�^"gc���)w=/4eT��ϸ�&"P�8��!$�ו�T�+�.�DU�0���֜���XEV�@8�έx���v�Ny�ͯ�f�ځ��ʙ�fD�H)��f>��ċM���i�Ϊ�� �\��#���t�gx�Xmth2*HFJQ) �����y��8,��D�N0��G+W#Jr�k��8���{�_>�p�(���sQ%�^��
쵔nPe�������R�E���Gh����[����R��X{ܲ-�86�T\� �,�v@2'�pAY,A:��EjH�wE�*6��M�(#�Z-!��s��q6�ʘ�J������ʪ̮�œUr�	��8l!�Sf'FŪ�9���E�V:�j(8cG@J
0%(��\�V�'5,f��[����ĉ�qA�q�"��xY�n�E�Y�`�;��>�8��M�|6õ\�C�V���
M���?mm��»8;��dUFz׷gF��%�?3sO-�H,پ�wI��A�������@i�TC+TL"�&xE�+=��sX�����v�YK��R�v�V�k�\_9��o&��9<f`�����$����!a����m������MvX���ŭ}�6 �\�J"U���P���|�,v����[G���0��w�l�ˏ�<�T�q�B��ح;M=|�Yw0on][��I��v6��%$�ҍք�Ѯ��\漽o3���=t�h�^��.s�O)0I�H�E��iS�o�i���M��)�Y4��P��>��U|����Y����5�u��Q�dB�-��㯇��d}��8�l�{��"Ϻ'ӞGp|�ش+G6涰����2,u��wC� *��4S��^><�ﷷ�5^�9�O��i�*oV/�i��>6�w�^�Ǿ⋑�޼=��El�84Oc��a�v�u�|�3���Ͽ9�D�`7�s��8Mܭ@��U�}�/�[��j��m����۔RT+d-+N��o�L�9����"��w���k���nͺ\��H}�X5��Hkܫ�r�}��~%hÀ�$b(������O����2c��s?;��B���U��v��;Q��p�0D���2H�2�)���Z�묇X�p��ۓ���ǵm>���oY��57���B7P�������1g�ލ���zl��FU:�w���0�>xh*�>%lp�����A u�aCeiM��o+�5B͎�Jn��7r�cȾ���⽋���֜c�2�\��]�IX�[�qb@�)�nG0�w)���{���{��p���eGr�}6N��ݗYִ�Q��ϑL)*J(��2/���a.��v�y�jcj��@i�.�G��Qz~��v6GwqC��ac������{��y �7����oWc��;v�^�ݻ "��qy����aA[�p�e:+K��V��
 J�T�B�QSzm_]q���4+�b�'s��bȕ:��E�9�|:S�.�Sj
m���� r;$���"&��]WTj{[��9�u�^#���mn�{t�ЦG+ex���X�":� VP�ۯ�o�\OZ�w�Ab�t{�Ԯ�4��gS=�s����H>�B�6���:z�4X��^*�!c�b\M��!��1hշ�Ԍa��=��Y���ף#f��C Z�:�.�����(Q�d�x:]��X�m(�u��Q�$�wJ�Y��PZ�@33�B��a�5���.�ݞގp\�t�y��j��[�Ҽl�Rp�
�=r���X�ԨjC�C�
e��G<)T�����m=���k6&����ё<�]�?����(=�\��s��u���O]0��=���P'�I�X�7���{���昢�t�2�wEt����*����^Һqj'���͘��+4������K�8e�K^������%෴R�eYB�to2/�/Y�-ӹ��I�n�1�*}q�i�
��v�X�J���{qu��Lcpp�r�X��y㣖;d�U���͸��!�9q�����'��-��y{;&Yx�(���ɲ��p�Fܷ�J2	��,����+q�=��Z��q׌?���Y���`{vfs΃Au�L���eoVV�1��@WY���%�;������@��Z3��c���#���r�º�8�LD�%
�k�J�=��_�.�VC���
[���q�+�y��^���T�{+gH4���
+�7��}˶O��A�����r�ɠX���jN��L=�s�;g�6���?G}�&�*���������ꎵi-��䨨XaD��I�����7��e��ԋջ�����aB�.)Cڽ$�.�{����{殺��+ű��5M�� n`=1Vv�c;�ۘ氕 �B����RUb��ڥ78kː�u�
g��sѷ�������O)�q�ӵM6m�����p�⻭�dE�OZ�[��rݹ���f�u>ӻ@��������y-j*��Q��H����������;��2��7/K�h5�0�s0�JKc\hޭu��������l� ��5��w�ɼ>����B�څK$�ٔ(4e�x(��=�;#&C�8L��̩%��MKI���4s�5���������rp0kE�ؖQ5l]��(�.��!��V���`�
`�]UC�3�$��@F	P�VP���'Vą�}����;��E�c��j��;T�w�=���]�~���Q�le�|����R�����Q�١�x]��,�R��"�n��bg9-��bq����7����
�q$�P�Ua�ts�R��1 ��Ny*����ˢ�yo#�74��lc��M�\�z����.)Zv��BR��JB��:�ΨN)��u]�pu��NK�r=�\-�̈́mT��+gz�]�N�IR����8���G���#{#��
{�Ļ�!���I)YC��Ϯ��t��9�{2���r�j�뮶cg:��Ա���7i��Fp���[�p���Q)  �$�P�)q찪������{ 3�g̡	Y�f6��G!���(Z'n�h{keۆ=O����}�Np���P�o�GU�ܣ~EV=��|૓+E������J�Á��i��T��Z�:�oMW�i�FX���(o�>5�A@�X�Y6�СA��Qhʲ�N�'��@�9g��}��s�{Gap�Ǜ�gY�a�E^���:g:�ZW.�:�L1
���	
Z�GT)����5���}"��.�X�9��"��r����e��{x,x��v��D��(8���@�`�,C��=�&���E�G_.U�:�����\�`OS5��^�����)sC�ʟ\,�D�;�n�ʄ��]�ܕ��5n�⑲�Ϫ�6��A�L'�a��$<m|���H��`��3r�Unt{�j"�����ojtӋ�TI&�wm;ۂ��d��m��r��\)vwR�ZB��h�Ը}ݝyH���w_���{M�u�IVo�[rs��´N+���i莢��2�]�ug�f����U:tE��r,��m���圬�Zz?F�zW��"�\��:\]e*�����o.#@ٌ݄XS�%�$���9`^l�k�h�Q���C�z���s�n�k'h��݅A���1��jս{.mLx�;=3�ͷ�-�(���c�	�G�}|���m"v����\b���g����9�¾���[�g�{���3�C��ƽ�vɋ��KQg�]�x��e��2�-������Ӽ�ޗ��p�����8^vo��<G/��.*�-@v�&E�.��٩k����F�/�_����{����ܮ��պzy��
W`)�Cp��ŷ�,��}�q}���OՌd{�R�%���}�p�N�Tz�p���ۀ�3�İ�P�%#�o���w+Y4�+P�Υ�?��PSO���e��\������z�j���Ա5i�E`��3ɰ���i�<��hz{MTvWx4�6���H@%B��qmn�[励D��vc�zwc݋�@�ԃ|�*�S��a�V��kj���%���n���[�|�A�{<��Ô�;��C'���6�b�}����,�󻳘�t�`5f� '_�%%M<��5���}Ζn�C�p�F�.��#b��Y�ǵ^�V7���bi�m�B��WG;sv������������/����(f�r'�?���q�J�!̼����3�5 <41- �wI�i�L(�ح�:Y��X�y�u��a��קz��<���]��9-�-��%1.[[�M*��/)؜�c��t�}���Cϟ&Ə�l���z��۵ �-�¼e�A��2�M�yk��ظ�����6�g��g��Y���9D�.(��!:�*P�6t�u�T.�lV�6h��hnP݉��;�]7������z>��Én�,$"�)(��G��a>���c��Vٞ�m�[|�y��as;\.��vWGmQ\e�܍�w�8-@%b�R6`Tۑ�}j�>��g{vpX1-M���\����Ĝ�_��]����E����IYf�X�"*u>W�Y,k��7[���3���X���=�h^iƐdP�$��2����b�>[����7=�g��$S��J����0���:>c��M���}�o�"U��C:�n�����E�,��5B���8��������s��:y�sD�s� ���z�;�p༵�"�7[��%�� �"P�EL�)HC!�v�/"�;;sю��˻WKu�y�^{&:^I[��;:�N��n��si�m��6�>{r=j<nyvo;��Mt(�cE9�4r��6�c�;[��ۨ�z�^�\����Pb�!Ȫl�]�It�s���=AK9�nx��θ�����J��^'v.�9۶�5�r&3��[`���s��ɧ�ع.s�m8�����R����c��Z�g�t�%��{[�������SY�Nk-�tu�Q}�]�b�-6�~�~6R����*�u�B��hM]`>V��1��UwāVi��jùBtLL��% H�(��j��۳���(�c�L��U�Wtm�|���OWt��9�N\ɱs.�n��3��0"	*BD"�)Ők7��͜\��]��n5�F./5�}6[�y��;Z��wb�� �	"T"�W��KF9=�dd��燝��t+u"��B{�/������؄���,�Rh�����m�UJ�)F�C|��f�O��n�P'��֡g,|��T��C�}=�gb�W�m[��=��բdů[�֎��ΰ�^E��z7^���#N�\������c�m	 �j աw�������oN��VA�m��yTt�v�╵��?��F� g�Ϧk)�tb[�
K>crط��A#^�RvJ��� Ҧ���[��+D<U^�g��������!�	N��i������fWN<q�����	��#�pnw������]��U�v�j)��-ۓ��ly\=��p�Q � �qc�ѭj���{&�����s�!EൺU:�᫸U4��v(X�[�1�NB�*$�R�L��U�k8Aʡv�S�X���a�Ƚ:k�[�G��}nu�G�˽�/������9���������"T8R!!pć��c
}u�]�j�<�W���}��������q#�tB�?_n�.�����ׂ:T݇�r���s��/��mY�죭��cQK�sOj��[�V�7�Tqyj�'��>y�Ht�`���/�~q~�=�
c`�Di!�
 (IL�)*ꫣNi��N�wc!Ԍ��5]K��ǄUK�<����vW�PX������e�]����	H�$L��)'B�׼'|"�ҵ���ͻ7"�����r�!��/qï��i����ɖWڶb�cx��$�F��^��0���N�rh��/
�.�7� ��,���u����iV;�u;듷��f���z�Γ"��H�!B���i!Of]d��^ks��������51i�缳v(��b�+4�ىF)9�!a�I)P�3)�ŋj�6�fSZ���c霾�qYcS}F�v��K�b�u[λ���]:gFd����W�DL�P�t�h��\v�Sgz�9�L�/eu�xPn��N��PԵ2R�G �-��Oo�D�\�*Am����(]B����=6j�ZFu�k�����tm �$�s���q�jl阽3u}Wz+v�N�&�u�X&��G��rf��j����H^��ӈ�t�$���`��&d��}�+��^�gfN���i���F=��I�s�^π	��� ׂo���/�(a����zv%��KU�Q�������+�]9 |":�ăf� ����ڰ�����}Lw0d�ܲ.6�aq�UX������b��Z�`�P<���}%$Y�Y~R�4B+7T�2
�
J�i�,��t⑘ze�W�0�����X��v�)͙��YQ|��x��2i<��y��.%TnJ�����Z��Օ5xz�wf��99;N�wV��H�$�B����E,�E=��뮶*�_leP�����C������W���f|���"�V��i55����c��<Y����f+��h�Ȫ��U_��(�Y�@�m�;�-���q#��$�F&J2���W-0����-�ֶn�Z6�FE�{�NsR������]��)�sm��hB�7)u55�kY�v��Y�)��N§�N-��Ժ���Ѳ!����U�y�׮�����3%�!4B�%,��d���-)K�fSO�_B�gɾ���G4��0k�R�ݖSR̀��/��Ŝ��cH�2Li��(ҁU�����jP{�6&(�ݤ�F��8�<�z~�7��0s]?n_nӫ/�QPH�NKI�����"f�{c�����qL�[A=4k�9qե�nޡ�ӷI!�g���n�a�{u�Q����&�n:1v9M�P�A�%ǳ�FU��۞$��]5���A��b�1ۺy�OB>z�����쮧�6��3�����mח���I�9��q���{<��r��xWBY����@��u�ݨ�֖�ͺ7[�%�t[ld+Wez;<8*�kOa����dK��:���7Bm���nwRXîHZ.rz3�V���-�b�M�UR'U��>=��.[��_+;]��H�L\���f�7�n]�/��;�)	2��,�X�h��^�FuF�^N@GS���}(Z�8��ꋾށ��Lo\�ɰL��A0�Hm�X쑶}����u>7^X���-���;��^Y=:�M��,ґG�ʁ�TJ�)e�~��g��q�i�NjX�s�#��[I��ToKܺ4�k�8\��Ko�2�y𝺁!~Kp��I��O��g��r���?Mx�n��|�v�`�Q�fU�U<WJ�c����wq�i�8��r�!6+e�
�y�ۛ�Ѵm�z�ĳ�\�m�g��=�zrq���L�<Zm�˒�f�-h7�Z�����ov�Z��w�8�\*����U�R��],�ͽ���}�<��*,T%.��]:���:��n�.�<ЙB6��7T&��j����ϳοx���=����7��b�V�٫��=��L�Z��I�]yD�m{gQ����ﾹ�ؼ�5␽σ<��fN6�� ��w�պ�q�m �`]�r�/��g���y�T�Ҟ3��{�zy!&:������/|���dW��� 4� �����Ǚ��(/�\c�}�1�������-��2Җ�P��UA�*T\�@�RZ��}�羻7t��Q$![�-Q���4���[�Y��h�q",���v���X�5jE ��r���٬i�\W3��
�	���=�W��\��!$�ð�v��7%,�s���9N�/&/����!�<~�kgq�V��WlN�#y���r�m�+R�������}_t��g�Ͼ����ǂ�$���:uGx���XP��+.��b(��ȉE})J���];���n\3�K]]�'�xy�vw�M�\G�vf���6�ء��+YbhǕ�I��ز4XRD�v�~V_yyWY����k��S�7��c�F>	���2����)��?���u��3�mMZ�Z��R
 ��#�n�{���8�LK�|�sn�|�)cQ�:��f͉s1T��E���99�g9bįRzR�[���$���r�k3>�Bl[i��4͍H�-����y`k�2}׵�^{��2��xq�3�.	�(ng�Z6��:�����Ohz^��3�Mq���jm�a�MYe1�/�����ɮҽ��ڮ͊��v�vY�{�w�a���s�غ��y�O�Hx)S�In@��#l��}ǿ}��7/���gf��z�ݡ�zc��v6���*
A�饿h���i6��e��,��({����3�E;��Z���c���/�Z/+��yW�n�-j�O�/4�FC��nP2��b/3���2ݺ��s�1<�\��E�m�N�Y����梫�2�ӵoF�K��D�Y�OPj́�,��u�*ʶ#&��7f��m�vE��m�&��<g���ݿ6��닾���>���% #
@JQ��v�{F���g��g�"�^K;=���=z����z��3�sݸL[�V���h!]���jɬ񱊞U�Ĝu��sʆܦ���^���=8<�i�L%#@�Dtﶇ�s���qYj�_Y��j�-��1�N��2z�{FV�~㾯p��-rVJe6$/�Q�佸�^��~�|}��e���f�Okz�u��E+�&ĺ����PݠZ��{~�魐5�8c�.9��sbbz�V=�]�����6XkWt�1RD�A$s70�3}�۝:3c_+/-���TK�6����Ե��"3�^�n��A8@8�"�o]dսw���:���w�1��:�b�QVF����3�6>�;�t'�������7�*w ]0�`�F ��[�mf�d&k�v���+���b�Qq+���wW��vk��dՍ�Wso^�mf1����ɠ��a<	�����sǑs،�{Ð�p8����a����3���7W��CNŞ.���Kam��wQȫ��e�k�`�3��{��+�K|K��{����-�]�	*��g��饬�x����{<��(���T��4��a����;�2�$0�#Irw6vP��0`;�w`b�V�\x��]������pO"�>�|�!A�j����n,!v��[���74S�hDȶF1�!�(m�s�W�҈׻�8�;=�q�� Y�vu�4��8{N�)>sV6S�����B ה���8&��h����IG47��t+'AcI[����F@{ږ��{Ŷ&�l|81�a-�
�m�+R��E�
��N�EYQz��xe�|:kOa�5"r�i��'��m��tZ=�(�S��j����}��']ޞJbpgWuut�G��b	�j�fw\��]�*��݃=�������>!��e�@=F��=o,W��2�.�zC=�����|r1�mz׎I�Eg�MQ,�7��iZ�l�sNK��٘��,�Z�q���VP��Nkc� �M=p����t����:Kfh�'�og���ۯ}Հ�4*
4d˕q..�F���cҬ�zwnI��nS��El�w�U��{B��y0��U��z:��4�����%�#�Ф*O����QXo�sB���5�\8բ�N�#�}�	���0{�����~n~��#BUM�I�<�ƶ��1�\m�V�KX�M�rZv7�Nq�pt�9^gt��.t�k��{y%�	ݍ�Z�S��۶���3vw���ɞ�Zy��6Cl�a򛧓	���P�7k8�l�ۛsZ5�K����q�`tm�pe� ��g��-:��7n�SNb��{d�[�N86����U�xޔ��'���mGL��4WY8ۮW�v�y;s��6�u�S���z �	\�ɮ��[�݊��h�n<;��:��{gj3�"��������:Ǭ�lvr�6͞<ۜ������w;kO=��<�>�����`�7���ڇ����ĝ�;Z���n��G8������v��:�vܗ����쪽�Zj'�'�]�wc�y�[9�%��\#�����C�ۆ+��V,��/
ۮ�d������l�-Gck�u�3�A�yZ�7��<��n�������0"�q��d�u�����=��µu�b���NT�]=��Inݻ:�b7-���)�>͏<�r
v��7*7cU���v��[c���Q�
�hV.i�V׵LA<�Vv��z�s-���I��r�ܹ7g]Q���ũ2>��ֻk=F�빎N�gon��m5��qs%��v�\�Cx�p���<�m�Gq��&�Q�q����x�:C6��v���W�7n;u�<��쵌x�t�nx�7����q�u]�c�{q��f�OBN�w<���B��n��kZ<h箷�1�kg�"��0a�'#�T�4�ꕍu��q���όF2)
�/<����mU�=����F�lU�ܕ�s� �3������Z��A�ۮ�Olh�q�m��nd���4�]�t��p=�n!��7d��g��Ong���vw3�n;T�c�x6	�m�h��⎍�uֻn�9�i��9�u��]���܁��R�˳�Z|���u��rv�n�cY<t�(
����sȘ���f����Q6ݷY��A�;�K���i<k�����5�^�,]�d�/�n@.�b*��N�\����4p��N<���ͷ?�k�X0i��q�5f�c�筳xvu��Gfx-�pqşnx�u��qpՀa������zO�������Ӻ�f��-������lj|R�m!�ۏ[v뎷GY����8�m�y3�bq��e$zݳA�"[���Қ:9#���t�6:�pg�G�A����B;S��;v���x�э��J�@ǆ���q]���Sn�i�Tê4ݲ&�[b�U���S�N�"�\L���%�;���ēgb�;��z��4n�����b��uE�k�K��sö�M ���#�u�]�j��]=[�4U[��R���nN�V�nY1�IYw�E�Q��+���ƧO!gm��gln�5���Y�2/v�3x�=;[v�����9͒!��>5u��N�ŭ/�!9���!u��j����K����� ���@��%$%-fpOh6L��W��}s�uv��[���1s5ǣ�z��Ƚ��u��H��;Q�d�&aԖL,�ؼ|�ɧBǹ��Vʚu�7E72�qk�r�XS�f`\��|��^�mEeV����J&8.��=��9Sq�nOIc7��q^ ��k8z�	��Q�Wʶ��wb��Y����l,OTg!&�
61�����]u�OgZ6���W�O+i��-a�Yoiž�2�� ��_�@n�@���+�zol�^�����y��ܐ��, {EO���Y�s˕�>[蠋�jL뻸�S��aRX[�o37�ZT��[�Jm-㕝��@��9d���9g�uQR:M]�l��}��EZ�Kw���W?_H��5�;�fT�##���}�e��HÅf������秷f��{+��c�⥪��q��?=\v,+��f6��\g]�ƞ�s=3��jTb�P��w9�u�M����!�BYn�PW���J7�����?[�Sc�{~v�E{���Mڬ��<t�l���m��els���4vc�WO-�{q�fێ�+@��P��W�r���;�<ٸ��/+U.��$���sf��59y���4G��2�+	f��\��yۛN$�9�⯬� ���7�=Ϟ�;�j�]��y}����u��	(�@�[h�tＮnO�}�jg��Z��7�I���dK^�u~b�U�QA����jR��i�:n�|^��{�:doN�9�3���8�����
��
��둕�"��2#�]�������m��Y�JtYbH���b1i���Y��v��Ґ�Ú7�_���2#'Nod/�����e��h����uz<I�I+���JNɞY�C1Ҝ?} �v�r������U�uL����ʆ�V}P�wo{Ǆ?h�bj#&G�r<\�#=�����Jp�A�6ힶ�`d-=�������pk��f(��\r1V"��Hmu}��f��12�P!��aB]4�m/��!/�)$T��ZV��f���ƾ�hh7B�e�j�U4�+.u������..;p�R���s��h���J�!�$������>�=�B.��d����پ���/)��ņZ��;���Q#BB)��М�q��w���g��k��
�3;�n���|�{�Gp6/"�b)�+B�ð�ޖ�s�$JbP;�Z n1�'"��OD�H��Y���[��Oa�����{Z��P9��k��8�'7��s}O��\\X3H��R������4x��U�:u�њ��dWZC��4Nd�t��Xq%�Xz����2N�%C��\�f�.�`���]�]{o�ɔ��0���"��4o5Y}mOWt��k}� �_I:��_TR����OV�� ��v 	$�	 $��E��U�js�}�om��1�&�V�-M���u�ʄ�s@Y�R�)���;79�+�CSHh$��k�w�Μ3�ɗy�ط(�k�e*#{^E-=V/�Դ�6@���h�#t���Q��;ү9�j��wE֦M���SWV�L�ӓto'��#.���`��@w|k~;�طV�Hb_�)Y�mq�PL�R*� �ǏE_:��Xh��g���̻�܇�C�I�˼Ecg�����=�ݧ��>~�ўɜD�X=G{K0iKVx�^P�����0��>�p�N�dj���"Ho=8� ��n,�T�  خ�nڡ��b�l�n��q�ܑўP���K�y�s9�1�:����"%:b�7n�[[�y�u���M6Чbg;c��U�t�桮�c�`C3yx��q�V1���>|�x�>ݮ9;E͹��&k5�8�<P�8�'k�w��ll�v8�G��ͺU��a�n�kc���7��+�7��{n�<��\�e�vS������j��G\�����6��6w!ck�C0�w��k��§X!�6�0��ֽ��O|=�
��Y`B�����=���7�����a��z��Oʻ<�J� �oΎ_���lϴ5�x�>u㷑�����:�nVPy���dD���Y�._�W܉"B��&R
A*k��o{/�oa�ۮ��-����Er�s�צ���K*��%e12&eR����,0 =�n����_zA�sX���ƷӔG ��5K��]a�YnSp��)#�qeU|1a�=A��q�L{s�y{�su]��^)3���6^�����ˊ"�Y�##Q��bW>����4�kqq��r��Lp�4�)��]��@���{�?�V&T����Ws�W�f8�23b����/*����N:7�Wkpr9@����{;���oq��nV�"T��m�U�6�Զ�[j���o2]8�����	������s6)���_�gwWO�0�>�㛣���*Z��vJ��=3o{+�Ssq�ηI�a���b��H2eD�(�I"��v�/z�0��������ʅ��Wʌa�Ӽj9]�sf;�Dͣ� L%�"�x����j�/��.�)笻��}����L�-�N�:9�oø�
���O0�4���D�
PFRFbTJ]�}o���C܇1V�#�f��
�ܬ�;���d�}�üa`������;2��m�ݶ͖D:Z�E?,[rmD�:�z;<c���2�w]��\t�y.|p���!%1)	��ƞ~~6v�u2�f�OjM%\17�`�'�5w���7!�B2�y�W<�o�0WqhQszj�/������c�7�>qd{k�nS�ގ��;��匦}۟=h� ��GD$��Q��^���.������Ku^>s���2�]��{�-|����Z��F� ce�Fb���#�q,:3b�®�=��-�/�#f)���)��l:�V(ΰN��[Siq�T�ʚ��G���7*%q��8�y1���y\�������ݓ�Ξ���X߾�n�e�a���qO�=�X����Kd�-Q	#n�N9���W!3ڠ��-�dO#y:qM�1��>���
��I�]���[Zj+vzm[��q��+��l�[=:��ǭ���'�3';DZt�{3�@*@������^�qhXzw�(g�X�p��5qQ�T��]�c0	�ﻷ�
�_�,	�������:sH��7����0�̭��N+���ΌN�nCS11��0�t��HB@�J ��T_;��K]�ŻC{��KW�ߪ�_�cF�hy����{����E%u��[A��z����Q-i}�l���ꢬ�WQ�{b�X��@��&lz4���(�,�I���#w�!��(l;u�j5��9pHn�:��Oy�0+v�nuRɜw,����v��Yҷ��������t|>k ��p$�H+!��ި��[��v�A�zk%�����UI���Gl+8λ��X�������J��'%��F��y�m%��d�z�l�t��ۯ\���v�H��.�&�h�Za��YB�׷��ٞ�+�]�׆��W��kh9We^7(����!z�d�f�g�O�rn�tXݨ�Z�I˯-���z=��}��fjR��V5s��.�Π]uf���Tn�\'�m��+m4���t��e�1=��n�e�&�+*��\�>�Yg|�����z2�R�r8�7*z��ހ���\��,>gRe��*��m)�]�jV�i|@St�\U����׷�����Q+rQ�G�Ie�8���ó�6g9šj?':�U[�����o��z=5�������od�'{�ay�ǽ�L���f9��(��
~�:�|Q�hb���$c{܁a:u`�}S[�c���/6Vjz軸x���T��	��'5��E���+�{3PA-GR�η�W���(җ9������V,�v�Mvn7:wO>_l�:�t�ÞzL�ެm���⁻3��z�sk�>�T������؂wf��un�c]�>��� W	���<�:{L�;v��kp^����w#�/�[����&��!�­�!89p�3��nb7��W����۫�ۄ+�=��]9�{�wDlqyy�%q�2p�ض��b�k��7kcblÝ��8P��;.	��G3��"|iy0�,Y��A��;]�mEI�[���ʃ]��bd	�=�����z��6d܆�]��o��g=�*d�^��K�*Z�'v�_$r��S8B��=FU�gN�d�{����&���o�a��NMv����ʪ��2���S}�W�����S�u�*��]�3�=`M�ŏ���u�A����>�r��흺p����J@�lŧ�n�`�#�f,��v2z]|��/��?���Ek=��q��������>��� �*��0�&����zz�Y�k�"F����{ׄN����;F��v�w���T�b�'5�M�	x�kY�h�Z��a	֎�v�nl���N8��L�vnʶy���N�[4�~���8njb�-[�mf:�)�㐱HBC]Z,�p���
�*�Lg�2a����j(���hW�}�2Y�
>�Hi<���Z2/	�5l�`��V�nd�b@��́0CM�w�BYZ�^J��sg��K,#ܲ�94񷼇�&����P�c4���>��>��x��*��}<-�{]�"�̇�ood�ݔ�d$ �BFBE'n�6���XLc��ښ�n;'Dp�;�d��/�a�Q�������y�� ��:Qm�;f& �[{9�9Uj��e��̾�p�:W+�yѽ��/مe��SJm��)M�*޽=�n(�]ڡf�iN+���ɂ|�_T��i�)�#��u��H]��#B�(A��������m��n;>՚�V�F��pp����|��;7U<�d�$�F	(��>���ʢ��('�=]��~;m��7w�:�3��k��v�^�>ys�w�$  A(���ёT�㿿�ʭw�L���'�"p��;�08��F�~�F#dwvj:%��*#t-HW��o:>�}(�^cZit��2"4��@�HؿX���c�6{��zkh�q�CM^#�*S����J�늌�2�!�ůBĦ��r��;�}�{C
ٓ���ͻ�F1��h0�e��ؽJQ�k_�٣$kH��+!A͇�1!��-�eA��ͣ0�F�*-A�ٺ{hX�1���DU�m!x_9Ʊ�<[�z��r��;�n�bɯ�`��"����6t�n֛�-	܂D���lɻ/r�]��7Pc],d�!|�Jg��Ω�4���sMk������U��TE4I⯧��pc���0}T%��Ri���`飱�y�Y�c�s�Hlx�{��s6f�u��F��R8ᝑ8Όל4�ܴ���)�u�lu7�׊BǢ��6:��������q�rP;2���e��'�]���q5V��t����H��2ȭ0@�[V�`��l�1])��­�%UCnb��@H;<}:N۶)�[�Ns��{��Ά3��m��YtA*}�Z'T��l�cc"=ӐX�Җ�����������wPe��g��}oN��5��G���zn�`��M�]�V��|��7���{=�*x�8��JEIH��r��A�`�m�������� �ף�h���`{�7�z��x@g��kt���.p�32v�\�,_v�m��y�T���1q�^$<W��[m��z��[�P��w���W=�<'ےϹ����1��[�ֳv�jQ?{���w{��I/��{�Pc�mX	�%\�ڙ�Uh^����F�]v��Ѷ���Bx6s���ʯ�x%9����j��#N��YΧ^3���ṶM��C��.>>R��"��ѯ�r��`�vq���
�=�Xf���~Rʥ`�K )y��y묭su���@�c;�o�Lhz0{��u�����Tv���F�A�+W�=h h��jO],��b��_O[�h���knŽu�;h�K���P�q���~��������wg�q�3GR�>��بM�$�c-���B���B�g�w���~x�����1��8!Fz���&$�º*PYǞ�6������\�2�����|�۽��$cC㥃���S�g,���0�E_׶�=P�di�b��Ə!�>�;/x;Ϊ���1vX�(�d�.Ii	�hi�Qj����<T����:|�:��+�Fq���(Ձ*�1}U�O��<�\8��(}�)����&�׭z̮E׎5��#��R uBX�j���u��H/��uu��Y��(Ly	6~?����Q��qMɧ�7A��ɀ �-/���Gnd$�-a ��!�^�D����A�x�b�i�Ӹ��=��f��m�y_��>������91`�һy���ՓJ�lt��ue�щ�lF�}S�i�����b�h�M�t��^���s#��r�=]�>��
��z�5�ۡX���Bd}��tڸ�$�C�T��W�����#���c��ŒN�����h���`Z.X
\v`�z0u {Y�6],���̸B�ï��ēo������c�m�_!D[�t�Ϳ����p�|Z�W1����r��a�m+?^}��� ���Ce���+��F蛢(]j�5ǌ��9���oD0��� �����`��֧TŖt���^�lJx���<CHQ�O��5 �0��	La���$0h������� pe-�q��㝋Me'���&ƛYb��~��GB͗��S��޳�g��Nk�<c��F�_|��|�=J8���P��9{�i)bP,L��H�q}1@�n�������3X:(FV��F�4cH��yf����Ta��K�,vsQ"-�y����_���y�K��G$c�ZY�~_1�Q��C�q�dЍ&�J�������/�.͞�h�w��s�-�ȣDQ:�����(���!����;���LR�?i�lŖ��P�O��ęH:�*�������׷��:�}�^��밥i٭���^�zd��\ķ�mi�[��[��̗�zn8�b��e��v�>���x���c��=f�v�p;q�{��;l����`��[q��>��]�tzz �9�s�Qz�[ms��`��=�=�=%���(7����`:�z���;h�.-�wb�f��3���MiV�q�n[1n�9.Y*^KV�n��	�M�a!�O\Uʼ�n;nwZV���p펱�$2�o��7�v^b���x\�8��l�ܔ�z⳷��sAa�E���g�s���4���=/N��6u���6*�B�LHБ�[klk�k�=�C��dY�"λ����hU�$�G�^&<�� =�2<u,8�HB0D�j��Ι4��"�dkb����T�FHS)�qǷ��/*8Gض�ӡ���RDRߺl�Dz�#�?�rcN6��r�5C#������]�lqbLY��]��W��oo枵�~[#���0��SscLe�t��?}���f4rcg+�Ƙ�F�5#�[<EJ�|��q�|5"G��)�Ά�2t��6����0�#��Piʔ�f�4���;��&�>C�Th������C���1d_��'�ي A�Ɨ����cD6o �E��~�eئF�F�H!a�������E v e}Ⱥ��_Z�J�ό��$�:�7�Ņ5�gk�CPpG�	ݞ;wW��1q4 �
�5GLm��Qj���s�M��
�+s�n���9�/5ycŃ��ƥ:�mKk-�� 4o8ٔ�bT�Y�5W��������G�ĄacϦ����4�>��EF��"�G�Y����~�}5<B�W�ѫ�Y�d�����$�������j��$��i�t4�Ĉ�Z�'�'��S�t�5�'껫��Bow�*����8�4�i�!Ќf>g�!r��3��ʃ�}�J~�+0%�a����j��Ђ����mю�L��Lx?p�Y?1c�vb��������c�׸�p½�+�:]>���?ȶ7�'�uQ��u�̼s轙�{�w+�'Ntő���Q܃<X�2�=�#���	,�^[��a�F�D����U��{1Wֶ�����4*0��8�<���A��7�G
�=]��}òl}������\h������C�{����������]d�3�Ɲ�*�[(#�!�G�FL� �ED��V8��#\��{��t4����Q�����C�n~�޽�*�'P�'~���$}��Ar�)�� l���|���GD�ʮ���ȝv�E���Kku�{\r������ݙ�v���b޷k�5ˈ��}��g����3y����m7?f������ƞzpǈ�iQkفм�#\���{�A�F:>�#,�J��'TW^|�af��ɑ�}�8�%Tf 0.��Z��Z�o�/��\x�F܅D��yn��׾���Q|�FC��M���Cf��5�~/8{�&Z���<t��>�e"L�Kd�n\�C58��Ȳ3���Mǈ����_y8y1��z�-5д��˘����K��ٳ]Y3�zG${�¥$����I/E8���c�ۇw��}�m����]J/Qcgg9�cZ���6��G�{�j<<"�t��#��;��O�5�wy�j��ھ����%�Lr�m������(Z:����uT��1��Q���f��,b�4~�}B�4/���&��Iy�٠ƨ�4������^�"6������C�k�e���/��+��H-��ǌ�6G ��r���i�أ�{P',;?�n��ѭQyCTn�x�����x*��t;g�Lƈ�D_e"�5�N����L}&RԐ���ˌ��e��1�x0��3�q�2]WW�ݻ!U$�0Q��p��8���Ʋ���p~>���W1��� ��Cs�1G���&C��s�;q@��n�h�M�㑮����c�<�Ǐ]�='�-0�%� M���*��XB�>���B�G�ns����-f<|p����h-QF��Tvя:���4E��ƈ�J�x:#E��c�Dv�X����1�#sރ	I#S@)k�|�Ǐ_��U�񕷧��Bv�ŗ(���Qc��$}�"�\�w�4���[�����1��/q#���֞�����,l�R�O�kN�	zu�$.�#!z��>6c��O��UbuF�,�}��4>;HQ�r",[���G[���u<+��f��� �w^����{�ܽ3��0'l3��VL�F	ݺ��V��7�)��|��TBd�^����������Ϳv,��sK���+~,mD�-.�"�_P��CLIcic�,�DO�`�{>�ɨϐ�$j�,� q���ٍmE��?\9���T���MfĪ�R�����;��j�G�������9.��-���ݎHqU<9q�uqWF��gW9��b��\����9"Lq��U�#�y:c�
��.'b+�!^}�FXcDVM�[��W݊<�Uy��=����#"I$\h����&,|m_����<�0
]��h���+�J�B�2x�> ��&��0��Yf�� ����Fu,�4tŶs�Q(�FDʕ40��di��ۿ,�?h���2��z��~���i_�ozH�ڤ�߶h{"΂�f�����my���4���@��lX��F5|����U��񻟓l�!�D��|�A�E�"�����i��b�������Gs����D�o�aK�ܡ��/�U��M)�r\���fƐ�8tř>���VF��L!�Y����*�Y�*(d�&Wr�ϤW�{��G`�S�R���q��d�X��<�+[��w�eEFEm=q#7-�C%�6�q��n�����Ogc�f�{��
Ã��Àjy�T͓��=" Tؼ��ފ]�:�.�8� ��S��ڢ�ީ[�i�;J�c^y)��^�b�A9ټ�9���o
�s���B�l�^ư���k�����g��]���gX[�B8�/h��O&^h�^��t����4��nzXמ��Ƕ�
�g�k���t��y���V��P<J�,_�^G�@x�Qۮ��=s�V�9�wVwmS�'v:ꦫ�n���Ì-�y�݀W4�u͍�]u��e�3�u�n�����/����lW$��bJHR���U�ޟ=4ތ��+��YG<�o�\G�o"E�"��{�Č�R����Չ�m
:G����acg�?���s�l��B��Z\�j?dUz��i`-(�,�fr1l.<)�2{�>_`t0�7����?� ��8�1;���8�a�h��{�����>����Luʪ�LaG���96�;�"Z�F�[cN�D;̺�}J��M�g�P���q� ���r���a�WH���Tq����8b��_I��"B%�L�e���Y'����Br��z4�7���q�D�����:�,����}W�x�p���>Q�슑w���2�j�_vUEl�
]��"�w\�t�u��P�Yb��_t�T�^]���݇�c��,�
��ip��gl�r�'�6��6G}�oxo�/n�ģ��]V���ac�h9�c��as���-<I��dK�;����nR*:�%ӱt�m��,#Q�?����<p�1}�,C�۹qkO��>�1t���ō�?;���HiFw�*ƴŐ�2��i|��`؄p����g�m1�<�x���l�xX�����Q:��3��5JV��;&I�6o�|�-�2goF��8 ���è��;އ�����]�<|x1�e=���S���H�K�#����W��C>\F����t+T\ɞ:b�������2���*Q��9�������J��ô���bq6D��}��q�D��Y׽.���ED:@��>�7�/�U��<!��B��/qj�!
j�@ʊT�R�8����uw>��Ͼcf��1�/{]6��Za`�ﾛ��H�(��H/��j��F���By���~��#�F�G�;���3-	P`Z5m&�^4���֚�g�uk~��(��4�?_��-�ҙo��Vzli�#H�k��_5�n4�#�h�}^�֒GįWj��^�f'�2��)UX'�Ksvsu�1��}�l�1St;������j�{���62��yǗ�z#Q~7���P�ے,�hq��m����Y�"��=W�
�5�?\�G|~�w��N8�zu����ˉ�U�	�ƦU���"Ǿ��l||ki�'~��I:�"4��S���x�
�L]g�o�`�d�"�{�*�0�Y�6��&Ɛ���kՐ# �|zx�_j!��5*�ퟬm�:�C"=|bƉ�����	� ��W�֐C쩾wݗ�t��{C���l�= � ѻ����������d+,�5��۶�]5U��n����VEX2��rj_L=��q�-9B4G��0�#O���q�,1tO�&r;ccu� ��Ym�����[��8�y���P����O�K���-L�#_��z*t�~"�5DP"�
=s�x"�+%��驌C邨yς)I��b
X�{��[�{J.<[ϻ2��K����X�½V�g*��E�G��0�ޑ����,r�#�A�XC��ƫx�Q<S6bq����9�5bS�GF�x�ֱy�n�����cgcr�r�z��te�l�˄�X"�-t� �8�מZ>>"��ng�q��{�g�3u�X���>����*���<A��6cD{<a���,)���(D�޸�S� $I�4�Sg"ȓ�Q�����CO`�>�G�h�r�a��;�q��,�/�O$P��yaĬ?1�2$`��U�]�hV�����|5��t��N5~�Ӗ߫�)[)j����OJi��m6�񯼮8�0}�(�ʃ�~q6�g4@��h{�]���I����%����(a�Z=��svDA�d�LG�q�jm�pY u%>���恕Xo�v����f�����}5�>\E�"]�*��#k��6�D��=P���Yu�S��w*�={����&�q{L�G`�9Q�q�.ګ�;R�U���W�n��A���:��%<����g
��\Ƒoe}9-�j��4�V�����nrà}����������ks	ۓ|'75Ы^#�G}��"��:���YAǶ~Nc�"ӯi�(�?qe�S֫&��m�V\D�%0ܰs��c���@��ɶ�wn���+j��b�.a �I)�1��b2���Ϫ4P"�'�h�7�}�
���mqa?Wƅ
�!y�<t�1�}^9f�/�5�i��K�P��tM8V�ӏ��Y��ʣ��Á[�
�ߐ�1�hY����C5E��E���·ǈ�H�=j<���Ƙ5g��A���g�(���E;9L���Qf��ϔ���QV��f�?���<�!�i�(��Q�x�<WG�	��������t/�*�HQ�:}25Ɵm�^��>��U^����X&[44�r��t���H���3h^��}Vj<81C�1 �a�K���{|k���W[0h�b��ug�l|����%���<aC�U�6~��n�����y��4<^v�5������i~A�L#�\3�>]�bz���Q�z���B�#�
ύ�*��C�N����ka!�&�i��F ��d�����G0����a���Oj>Y����W�b<c/��ޡzv^\z%��JK��4�!��{�n�\$����Czڛ� ����}�WsY�$H�
� ybz�^>����~�S���v��#����b�\��#F$s������bjr�]	��HFi���fټ��7]bדA��ꚥ�@Y�*����ۅ.�/#p�9��~�UsUh J�Ȉ{��< �'��Q�p%xZߜ��A�W�І�N��7+�P0��;��7�G���λ�N[��d]b�s]����Uma�ʟ�qO�9�f�w���7��}��xx&�4�Q��;�����Y��V�g��txn�3j^\��	�s�@�������u�z���}���=�{��p�#�)�=���f�6�M.z{����^�J�e'p��\�ؤ�)��e�y9Lo:�<�J��ĺ�f]��|�-N�ǻ{#^n��T�Ouư�;^^ތv�.����(�nF��l���
�j�p��ylq�o`L��=�êK椧������[���B �����k�*cv�B�0��B�=�l��2ㄚ���4���TRf�6������ȟ������x�(���-eq��P�#q��x�M�H��
o�t��*H�z�b�N�Uw��o����wݸ2t��'<7�qr�����|9�]q�a�Iܾ���|�cz�^����;5*�o���CR�v���ѴJ���f'�5����~ʵ7�G�{�v��&ޜ��q-[.f��d�M�S�����&5�?(�	u+7@NŲa������H�e]�SWq���mu<�Ӳ=���p��9��}�'�z�6�<Ȟ��vN<>H;��u�q㗞�{<�v[�����(�� �W[�R�I�|�Y�n�s�S�x��D�7m�Y�y�)�Ltm��ܻ/,�ogb/& ��)�����rX��X������v�7j������t���Q�ge��ݣu�'m�09�ns�M!����<�k��
4���dS�Ya�Jt#p��u��n1��s�u��w��K�t��x�E>5c�&7��ش�n�n;�0J�ˉ�u�����|�۞�'K9|nVn����umΎ�9�Ȧ�u���b��r��r僸�M����>����d^� ֐�ø[E�g�E�e�iESYv��7�WAB�zI���csͣڏnxnض��&��m�n{rF޲f7gnՈ��Ov��Z�^�a}�������m&�.)8z�m��؞�9��X�s�{>w@u��vx����8���֕��xN�tWs��v�<�k�6��m�\p�����[!�1v�ج�[jf69x�8�;�h��=<�MՌ㥞�W'ct5�6��6<>����Z�"�
#���q��93�b�7OVq�vy�a��Og�Z�ջo8t�����Y8�X�n�%m�99�[&�]r���wS�t�ۗ�CP�ٮCr퍙�S	�]G�-m�.5 ���qՔ[\��G�ONu���\�q)�j�nyE6s�TO<`�l�-緪�gw<��a�mS������c@ٞx3Bm���������^���|v������L�ħ/nq���9�7l�9���Nwn=�������v<q�΀{%tp�m��J�����cu��sݠym���b�[�����9,�n6j�erq=�;v�<)�Rur�u��]��^t����1]��\cs�c�;��u�LsOv����n����}��ܬ�����km@�2���	x��䷹s���M�`�����%�͵�zca�e��럝�3�c�z�C=v�m�{[�WqѐC����{h��:�l('h��Y���vd�^/4V�8x�|O\=Z}�R���s۳���ೝ��A��sQ����Z�+nݥ:chݬ�k�'L���\��ଡ଼��M�f��1��xڌ��m��E{=��� �P�6u����=v{1.9܃��m��ay�O;m�q��؉�;��������iS�Y�u���Q��۰��o'����&*{����ƭ���[{k�ز�;��o�b$�
�1�}�*8}CÇ�P����6>J�����i�~"��·<gq>E��ڸ����'���2��#ǩi�40Ǿ�ha��ښ9�cw�D���=��_ۘtP�!b�������-h<G���=w�³�	1dP1V{��kOK��m�+ 6 �����t�"��˴�qc�
>H[��֕[1��[�R��F�ןx�cu
2E�³£G�5҂>����Q��$ �Qm�sq��Q��E���&<���i�	��fO��To!dm�E��s��yE�#Hν��۬۰�����G�iE�\�*}�KT#��
��:�;&�$H�>�CL��酽#K���H�H:=������.0�zA�}�B��i
�K�}4�V�R;@t�$�tߏ�����73�6�OK��{�4�)��ٹ����%c�\�4nY���lp��[xٍ�,�-vx�ҧ�D�8}}�5���6�=�Aw��d�#jS��w���#U�K�F�ş��(��jn�򍖲�q�yZ�^zk��T�]�_���}F��(�f�l���b�뎓�y�+�}��l����ws��M�=G�m� �'����חU�"��әH���#5�h��~�b�b������s�T2#1p#��}�s��"/�wE|��,A��:�3n�j�T'Eh=�MW�Ȇ��w�#���o(�=�UF���U�C�K��W�j��6oh��<k�8ő7u����jc�;�x�ۖZ�����J�@���� C�s�ђ��q���G�!��T����3������>g��#�մp���ãvpQ� MX�u�M@э}Z�ۏx�_'����V1�I�q�,1�+N�����68���\#a��`QG��1gٳQ�3m��'j�EJ���	|P�V�p�.�?{"�X��q��2�����G����P��D������ˣ��N���q�<��E���C���n��:�傉��`ԀJN���=���^����?�4!f(%1L�������1�zv�T4d�Q<WH��["�2(��4�P��<l���>3:���R�Kk�wR?��b�Qy�p�ei�b��O���5�F����Q�u�G�6y�|�e��*F�Dx{�YJΑ�SQ�N���D��{"_����5T�ctm�Cko���G����L��@�<��@�1�(8��j=u���1�1za�O��c�\8	��<N�6�l����j~,b͙�9k/@~X��sà��L�E��4Gω|c���{:y���Ǐna���# !ԡ*���7��m񯉶��֢�R�Q2�S��a�F3�bm�ud��x���|�q�aj�3���3�5	h9^"�n��жT]܌!Hf��|�}/���#�v*)�5����v��ʜ_M�j"��Eed�,�!m�!�,������,����@��LBbE\4���v��4p��;�<E��(���ha���>��A馚Q���=��9���Ê���:=@�[nͷ�Ä�n۔�>�X督]��a@��u���tqמ������ᢲ��;MBB�QGR�ϾT0"��x�1�jx�NH���o�6����n�=5G�nl��'/������iJ�d9��ΎQ�q`�#�[��Y��~���<,g�(Q�?>�a�'�?n!��(ß��C��b���������͑��-�ЪJ�Z%6��q�Q��Y/�n�=�#%���-/w���B��Q_ �>O�m8D�g*b�����
���Q�.:qx���]h������=.��mn�k�=�ut���Q��}�#�M���0�O�[�:c%�*��ϾUE��3��|D������>ԭ��]aev�-�[)�� d*IQ�4��I\5����ȳS4��1�p0��������N�u`�^��}�20��_ �l��4��fKE�-6�i<��(�2��*cq���͏-�yY�X���||���A��F����<G5�P��i��Q�e�Eq��0��\�Y\��:�F����=[����ʷ=�e�rZ��=���v������:9�9��ص��5�E9:ֹ��j�#�t0�Jq��/�W�+��F$�CٞϦ�=>�ŭ�V��fH��<������P�$N���c<�W̅��;X��:��^9�5|����I�-��f�G�F�:+w���,���1W���j��QÄ|��UFlX,�	(�"k�"���k�K�(���	��Ʋ݋�-6��g�MA�8�J�|��t �Ő��c�m��H�#[̇'Dj��40T�	z���u6�ч����z��<B�')$`+�8�1�$Q�M�X�.����4őCIB���ޜ�Tw��$�!g���>���B#�PNJ��W؈�y�#�uG��?��q�s��Yl{R����V4�Y8F�xd"
�����G�#O�P���s^�/c�.4}B0|�f��4/ĭ"�e!�����C��!_)�/{� F���A-Q�g*Ðj���Y�q���6���A�w�6{��"[�}GN����>�Y��2����`�����)�է�
�[ #LQ	�vlc��;Z;+�q���b;5vs��\��m���9�u=�yNH�8*�ٵ�s��\�\�m�Z^9���v0����'��si���f��Ymg/���\v���n]rI��:c�V�S�u�ca�.��N5]7e��.�2�j=�{v�{!��ϫ{O�Q�Mn����r%���.�U����v1�m�M-iwj�rd�u�Mq�d]��#��;�
闵����I��.�!���/;�6�\�v]��K���4�2A �ߍo
d��8٬]�o�Q�!�A;��C; dI�A�o����~<G:�G�Li�LW���f�F7�[G�.<o�񦦼��?�Z��u�~f����cvb���a�Ŋ�G�y��#m]&x�1���
�����%`�E݉#μ��N���t,V���.�Ƿ��;�ɧ���ƈԆN�"�>��¢�!G���r���r~��Hj��[#�#�qp���3�G �!�Y�|��jQnK�tK�Tƶ��*��+yν��?��ڮ8�sf1l�1ɇ�Zb��=Myx�>��$���	}���/��Ur��4�*͛�l��a,�%���GyY�|����١�|N!��j�^�FI�!��Zj��qD�q�4Ew��T(X~H�0C����T�Ε�)y1��C��Ń�,ǵRoC�'1��KLlv��t��bݜ��c=����W��Ç�����Z�X��a��ω�i�b�k�����o��1����.0|�\��tw^�8�>@q>|1��(�0�o�Zt�F�����}�8�P5E V;E�q��2������/]Y:�y��dI��.�&�̠�)��Q�����{l(�JAΒ܃��Ÿ��7�vz�����<k��o]��<98#c��6}��4>H�<x�7�#W���䃪,�g��91���W׼a��!>��<��Z~�|�)`[���W��]|���V��K1;��0�וv��Ieز>Ey�vb�dV�44�y��Y���CLH{$�:VBϼ~D��MI�A�̤�F�G���sb8�kא�1���0�B�1g�}�MG�=����[��t͘�(i���>���������<����c�i��'��b�N�Q2�P�(�~hY����'�0��m�v��򯻇mU�b��p�Ju�M:E����ɏ�\+eq�`�C�=�||X��hMu���8�i"�a�NȘ�vS�6�F�n�!��y��7���0V��IRR�q��������)�|��2QQ�d}�Y�H��@F����>��$Ut;C��|,D�����xp��0�Z&c�~b"I#��KM\ri�1�MU���]c��4őCV���Q�M&G�7��W�pP"Ć߼\<�"��Ʃ��KQ�#��6d��01������'�"J"v�����^�Qi�}���&�����0����*=�(�+�=�g�>�E6����3�0(�t*���ZA�(�E5d��[X�}F,@TD&����^�;�ve��qP¸tc����AR\%z�5Y#�n��1diZXP���U��0��f��L�.S+P0W�L��q�q��]~j��ߧ?Fa�0�"]��A�_�1t��W�(T�|E�p�"\o��8�-��S/�v��Q�3��.a��
e̢��i��1<�ϫ�t4�Gڢʪ5 +NN_�y�Q�Q$�"�a��ő?&(ŏ�f7�����?h.lb����͵�|b����J�D�N���o8R;[7����v�|�lk��F��\籽�)ie�F�`�,	��4כ�Zj}�_�0Y�ײ��}r�1/>�PcV�qo$C8G���<#�>.����p�E���Mv��+�!�#>�䜩aL��)��T$�x�jI�����L"87��k��t��#���>�BND���Y�3� (�D�{EF���@����~|x��[\wh%���(.0xT�X��
�8�������1������f2+���>�F-�丳x�t�bG�4��}�+E/���F��.6{�;PGG
�(0.�ǵ���ò,��CO�g�<~:G���$�>��q��!�!����Pq�-�c䄺=���kD��IߕkҐ�rβ���M�8C�[�<�FZ��m-1R��eM������UB7uښY�yXNc��>�%��
�0���,%�5���lv0�(�Dՠk��E���_9Té	���X��N�I��p�H Z3|�|��E�L3��Z����h|zУ�<1G�ϹX�hf�����m05�����pV�Bt�9l�@���a^֣���W5;t�nţ��u>���H��-�%�p�c�F�|E]_|�N��������P7����c����[�'|c�Q�r������Y����'�x�Ǟ���5E�?�;H��tU�x��`�#��d�i����Ie]eY��s�,�[�*lş�"��֊�x�/�2���ʶR1Xa�H�y�k��֧����!2��A�{�G�:�"N�o�C��YB�,}��>��E b���|kd�6ЩthN�����:��^�s�a��9�WͿ�	FY�+i4��^��:�l#yl�4Y�S�|�\|N&a��	_�.�Q�0�#�XC<~�5�q��O��1���d��ϧ�y2,}F�X���lG����/[+ER�}yx�Y}�����{a�l��1���X+ԯ�$�v��7#)B�x����X��b��W���#>��#�jc�ة(��+B�sْ�	ǘw�|AE����w\�Q�2���)��!�`j�b����u��OU�5��کMP�h"�+��d��T�<�C���l�Ӷ�룁�m���;�Ӷ�)Ѣ�ӵ��'ezMF�>�o<�{i^�v���#A�ǻ69�X3�z�����n{����@��V)�U"���p[�y�qu��83��C�9:z�Û2�-�c��Ni������Çcdy����,����ɣ\��:�b�=�q���!vuv���H'Qtak�{M�qn^@&�:
\m�ݢ4/�n���hl���B�����n��>�;v�m��hr���kg��f����,#�6hI����p��iG6�_��f��4����/g�@�kV�`����_ah�#f�$me���=hi=5*�8���;h��{yx�Qv�����{�Mz艫�$L5E���F�&�x�^�O��vM>���BA�C|~�o�!��QX�i����qƶ�U٨�ݕ�GG
JV� �{%9�!r�� `;���>={��d�dG�����>�f=Yl��o�#�x�^{�E���$bG��N�ݯ}+�C�BX�Akk/�V�G��od���!��އ#�����MI�許�H�����3�x�,ً�4�p �8��Z�K�8���ĉ�7~���:�R�+mi孽&��o������fa�t{��O1�%�K�#Nyi񌐇���Q�Q�F��DϾ�Cǎ��q�`���D����r��dvK��vZ�W<�5�\OOd.�ݶr��d��z���� �WX��a2����ig�g���+Y��N�#)	��a�^�ϕG��D�^"��ƻMY�1��V��d�����/�Mj���1�Z��*���Rg
�$�,�����cJ6���,P>~�qC�o_�oރW�zb����d��� ���5Θ��+*7�ݾG}�b���G�~=�زP�K���p`d�\v���9�����6k�>�{2g�<C�����S��B�~w�v�0}�F����������Y�ms�e��JH�GIg"�:G0����[f��:h�em%o��؋�8L:��#�0���#�{X��gK#J,�Nl�_�p��4��.�R�x���/J�ŉ�L-��b�9xlɻb��ƱٓF�2>��^��"LN ��
�ߝj�D���P+=��(�#H�7�
z��M�4O�](�[2Ʒ�#^��`�QB���]c�Ĉ�{���i�T8�G��<p�(��!�A_u������Y�WK�4�u�r�Fj��3m��8WH��O|��������(��f��*RHK��	�ނ��q���`c=��Ʈ{z��a�h���iQ
�
RG(��]6L�ǼŶ�g�.Е���ܠ�@�z/�qh��Ȣ����Ƚ���l���"Q�~���cK=��yS�q�F��,"���Ҋ�h�XS X㜝���>����v�޳c��1RNp���d8ߌ�xet?�pbCE"�y���i�*$q�<E{��#H��eC]G��&���&�E �	�G���L���0��\�x��C�����Y?P���}�{�w��y�Uw,6�ZS���E8C����s �>�X.�z+ >ݠ�5]�ɣ�l\��F<��קּ����?A�!}{�<67�*�rF7�;�G��y3���FM�N#�RX#�4 ��t������ۼl�\ϧ��\}@<f����7��/�L��<N��{o���h���|�n+��4Y�|sg>v���K�C����3�z����n���`�׊�Y�.Y��/`����^3;� ���t%��Vv%Gl3 �#���)�Og	�g����ܻ�7y����	����K�4�p�^GD��z�Y.�״\U:���;zi�6���Nq�M[��q�JW`���vVsG"���Y�p�����O������Pv��#g���<�P�U{|}�ͮ���T�=�gpZQ��x����!0E3�� -n��$��;՗� �Y���ڍײ^�r��h4�mƩ��`IA΂�|y��G�w��\5[�{��I�Z���5W<����Kq���!��r�����ǣ�fD���d����A٣)�=7��:�ǻ���~�nP=�m�<f��7�M��,�v����wkmM1f�M��١��W%8��xpS��od
O�O-�xj��P�����^8xA@��O&���	��(:��ψ���m�KC7��x����ա7M�y�q��Μ���`�KnH���9:�A�L֪���t���OZD��`V�I�n� dԥ�dS=�|�b�_���G���#
�p[� �"-��뿧���^
FR�G֡���j5[#��7�W��ϐ��*�0��im�G��U���[;:\d�Rq��b��Y��|�/P�E��xh,C�[�E�_�H5�Wٸ�����i�*}�5�8�|�)������b�>�/>r��z>Ͻ����2E1�L|D�|w\��h��f���90h�$;�~�C1q\�ȚC�{��JV�Di�,��itǣz�����J�!Aڝ`�o���`S�MۃS�4�w'���ͷ<q���GH��"RI�17d��z�qBD1��H"��D�*����
���9�l����<��G_}�a��eε��YDi�X`��-���AKL�lql�4�\�x��(Y���4���;(<��6���:b�>�D���BN���Q��>��M;\B<�1�r���o=�{��y�|����B�K
8�pٍ"�fU}��Ɛ��TY���xW@��a\�;cIu��m���<��q1\��t����8����e�0��⮋���U��GG .��vi���~��eԷ4P����_h�l��5'�c�,�D��F�Kg�L�e{��s�,!!v��ka��V�6�U1���`�}��[,py�e1���N`UHt5�	��.�y'��q��î�K\/E�v+^��fgyWĘ�6^����������r�!����yQ�nE%��
F�`$p�z��1'wd ���$g�g��"H���Y�׮�
�����}_�qLsU��q��u�営��˄"�VϾq���\�!�a��p�㔻*/M��)��3�=����k- ^^���5^4���l~<E�$�)6b]��CLYck��ފ1]L��j����L7�p�:�^�\ypV�E����P�`�+�N�3gĞ�!@��i���\X�^j	>X8�����v�Y2�3�Y�C�Np��q�8����ݳ��pCǁ���*+�p�z}7�����I#�̀!��)��#�ag�D�s�{��0ɣD�"W������)ƌTE�^�)}��b��Y����$GW�b�u�V��T�S���Z��+(褬�Q�R�G,1�圸��&��<!`������2�*W��騭C�Gg�@5ޗ�<-i����LH����b�b]��C���2�gF�Ir�@��ne�cH˶��5�a��8Pg��P'��%FŲ������x���S�.+Z"�كAs�y��4xgu�"�X�[�d���
��W�#6��!ם򜏈ᭁ����p��F�u��^�װ=̕(�������._	� ����9��g�� y`�����"=�F[I���u�G�َP9ۃP@&�B���:�s��vMɽ��1��g�����|ݺ��
̗8Bz�*Q��t��Z
�5[gn]�<X+)�I��q<p��k�;n7]��۞���uvk�fˉ����q�n`|���AN�\�5^�+��xB����3��������Lvc�#j�]km�LY�g]rvtt�ig�pL�3�Z���<�Xy�.ɑ�$y�pt�#�WJv�Y��QnKB�r��R��y�_]��Wߕi�a9��q<���E�:�!y��E8��<9
��Xp�ˤQ��"���o>k�k/�O���HZVV�Cm�|��Մqp��/7'�+�}�a�����In���gH��=n���7��<D�d7��P�Ē}��x3}o��j.�ֽ�e�b��(ظ�s�͘�Cօܩ��p��i�6��*�x��kH�c��� ��{g���m����Ɖ�����s#������Ǌ�����l�P�����Q�0�[�r�⺚��E�w{&�ǈ�!fH�7����(�d��'��`��B�;Ra
!D2Hx��ӹ�`���]kO��]�����T1Ec������6C=Ha+>������f,���"�I��r���.�¾����#��C�t��Y�����q��G����RȖ>����vϰ�N�ee��pus�x۵V�ݹ�Bv�YϠ���ܧ]�=��ӭ�|u��6�5֭'Tr�����P���Y�u	�]�B�o����M�w��q0xő�u���ڹ!������(:b�<o!x|/�^!-c��JK���o"�ӏ�ͭ���q�P߄�ꞷ�Xc	م�g'��pr�e{���g�9`wuU�CGj�*2�F{��f9`�&����䭔um�m�:�-�}�n\)�A���}������L"{��d�rV�!�k����Q�m��Ӱ��;���׷��e�.w�Q\��Z��]��4fL`����h�~���~=1a������:����ch��d��dx�{ם4/��ad{�
>�z)1u�4����~w�!(( �H�Z~~�lk���$��ݚ��҇쿹X�~=���Õ����h��F��B̑/���E����k��4p�w�4F��{�J����7��(b9G �5����֞Uٝ�E�����0�D�a���q��C�4cC`��	c�����nhv���֩�O}��8aC��)w�}L��n�9��o�d�j��uT�)[�^�Lq얹m�a�WG�#	���϶ZQ��'��qZB`�{w����][yt����+N��D��G�>���=��M�\�e��y���D5�F���X��,���v뉮���Zx�ZS�O�E�Gh(�T;>fc���'�5�)�bm������G�Y@��"ʧ�9�Ԩh1-��3���(�Q����c"_ۆ���.iv�;�<��}��u�FQ �@�w46caE��Th��C>kʾ���C�Hޝ�XϾ^�����^6陠[�D�ٸɁGH�'i�̟o��~�:f��g�p�-͜�5��W}��r	�3��x�� �׀Uƅ�y��y>"���!���8����v�ƞD�N��~�T����4�D�J"J2�(8���͈���y�X��/3�0�Y~ҍ�o��ЭCNgT[�x��lx���\��C�\�A'�)�����:�銋A�؜"_���i-RP�K�k����w�UƴO�-���`�(4"�G����My���A���>����~7�GvI#��p��q�θ�+��&;�2wu��}F+nΚ��&�N�n�;��p�S���<��v4�lvz��� �XC���-���b�A���i��3�(�����Z����r���u�а+�4�!��� w����uf8XHK1/��F�A�W�u�m�-5}�k+~48�}�J�v4�GH{+�FR�"����b��P��ۆ�#���t;;'���������{=��@����r۱�J�*�(Y�g�+�9Ж(��"�O���C5i��4nP&$H$tXt�x�ʼ.4X��ن��T�>;cL_l�!��!�F}�,�)���2�Kb�,���1����֑&o~��Nz~#���qԆp��Q��E���D>~i�i�.cDLc�3N��.ɚ�B�.���G{"�^u�ݫ2�:]ll%|���u��rV�;��w�[���90�P�-�ge����7�����\��&8���Uy�Q�8e"�ec`-|�Ⱥ��f������ֆ�˼�ǈ�W�g�V�}Ƈ�g�*a�����ϧ�i`��D�ك�ZC./��"��/5�2Q������A��&��;�AÚ]� ��M��Ktv����f�r�DQ�R�6�'P���ԑ'�d�"�Y�~�b�a�@�tc��ޗ��(F�@��1�W�.��`���=�;����6</�ܜT**����'��h*�#t��+�P6t�c\��7��}�㬌"��.R;��]>4X!��E��=Y<cZY�TqrD�Q]_[��9đ�Q2�N���Z�}ji�}���6�J�%�-��'Wj�u"������V;HY���h��Vuߕ}}�/�L�?�aV{�x�O�GH�&ŬhM}�
�8���^s뷁g�%m,�8V�em��da�l�*�O������;�W���b���(�0�:�ʾ;�KH`�"�)�VhA�W}{ݑ� ����Yki���e��.�����M�!b�����@��4�,��㲅L���V*4b�3�)P��p��1�2jU�2�s�WG��;��
u���D�2���c�zf�ٸbN"�'wtΐ��%�S��t*�j�(����1�b�cS}�̸�鏟i�okc�7�����1077s��|	t^P[n7lV�����\;���N޷��gFObϨ++u�̨WRlm:n����&��r/f�y�gA�ݺ��n.���Lh׬��7=��y��z��\�*�8έ»//f�nS��)�1{u�<pvw���>��TŰ*�{v��ݞm���-�;�J�U��!���ۄ������2����k��m�M��=�z�=Ak8	��Ú��j5ұ<�Y��a�[rMg�3��f;7o��Ӵ��Ϸ[��o-�72�����#�e�Q��>��q�0�
<}oEY�RE$��;�V��5�_�aR�|s9x�z�0C#6~'s��>�W���g��!,���� O������f(P&Y�d8���hE�*�� �w�����1��X��O�t7X2N��Y���7�q0,$+gs����o��>Q�G
P���,�#�*#K"�=���xG8`�H�\��oƃ�C��ځ�=#~A�a{~1V��s�Cp}?t��Cԉ�1C��8թ&�ܕ��a�٭��|[�Z
�h�-)m��O�t��W�z��\�~�A��y8���Dň��`�d�2\1���(iM#�]h��(����|�aL��&Vmr��E=��ǈV�:|<��}���갅��eq�����v.R}�q�ل/�Y�TE_�m �Uû��]���Κ����C�}j�2�E���b6c�n��EiAf���7$�����Tbc���26��H���!;i�q0=��m�ک	n�ص���̶�	�[B���c`1��Z� ����q�1� �x�PŦ,|�f�^,��+f�~��:�@�`H�,!�u��]�SP�]yws�~R?I�����&�X��܅��.�8Q�;���8耩o�}����|�ʳ�Uы
D;}ҮU��.r@3U���r�Zy�o	w�1fn`d;&	:�	��`�ed��a��Mu.���������W�}�B�u):D�N���Ma��Y�#�x�~�����0r1��{!�Y�"���N�A�A�,�{zk��i��	︳���"p��(�`���x�Ela�`�G���Ɛ�`�����.�Ӧ�!{�nk������s=������[DV6%�&fhi�#5;�	����]����^������8ay"��W��ί���Y�����u�3�N�m��0^�*9�g�^�CP8}1�}G�f_�_��+�YY�ڏ��+�u����X�Cr�DI�4�<E�����7�Z�+�dp>"̑^�b�h|5
,��������wT���L1􊲂.��o���I��ۈ�<��y��Z�[/l��mj��.����fN�I.}�;M�h��"���H8��o�MG������PCU��{0�a�$ؙ���(x@C`�d��W�>�p�+^$��9���!�x��=QIme#n�)Xߧ �����ˋC�P��SW"�C/����Q��#���K�#鷢��T5�B6E�}�q�#��/4���k��m&w�o���#��--`j��Cؑ����r�E�.�t7#���(oX3h^��*��;7�]y�܃'�ͣe���4g�b
�e�.j$v�8�:��Iu\!:��ݧ�Sa�0M��=Ys�w��1�:�u��#櫐�>�[1�c�+ڇ�ę�3�g�[�m�W�+�К�^s��c]�#u ���Z�?y�P�B��4�Wfg=���`Zp�9�+V�_?
�b�Zp_i���:fn@�3^θ���'ft��Q��y���I�$��e1dw-���w�X4��Tc|}#M� �e����w]4l��Tc2̣�g�T/8\�x��P��ދ��ǈ��;�.����e���2� ���9^4��<p��r<���Ȕ�`����^8���3mv������ /�k�=6�}"b�����"��3�x�t8��$
�
�B�@k��q�7�Ѯ#&cب�ޏ�u�"����=�U�@���3�K��Vl�8�F��Vڿe�5Ǖ���eW�}��#��օ�]ׇ��(�C�|���¼dyE���`�>�ߦ���Ŝ.�E%��B�}©��H���(�e��|�hw�s8�'a	en� m��<���l9���8�%�s�T�����'G!Dy>�{L�<��D�NGu�������R_�Mit��?M�T-�2��7 �[ V��4��x�"҄;�|��'R:7s�7Di��Y�Y_}z(h1�d��}���T�
h�{}_eH�$1=N���W�G]�{�7ԝ��\鄺�;��5���~�����ߑ	q=�`>��Օ9��r ��oEW[w���=G^�'�\>��D��e.�<3�fBAl���m��8#A�g��+~�N�r� �[�b��C5��g������`�(L��dUA�1!�#1B4�x��7���h�e�KLH{!	��jБ�#9+[��ی�ycy殺2K�W9n�\fN���Wn1ʔ���gR
��4��Ϗ�JM�����dq@ю"� �{!� XP0 c��to�\\o2%%H\���#Җ�r�����Gu"$O>�a�Q3z�ΡKA�L����2�ü���}u��44���h�A�����LH�gD1�b_S+��qa�d.BN	���.�<A�˗������3��*��:,�R$���%��b�����<��$?�oڲ8�Cr@XںQ�;I�k�?�����'SB�6gD����g����%������Z�5J�;}��:F�<����s��m=����K�,�E(�;�}p�w�]jD��H��p��Y��N�(��!���13)�ޡ]�;�����#��#D�q���>�R��v��@����C��		���ӖI�p�]W:,߬i��L١w�F�=����Z�=U��Q�u��A����5@�
[EȨ����t;�j�ϗk1=�w«s߀�>@��]��������_��ziS��11����"s��&�:}=��O��{{J%l�Â�f9�f�����{x�w���L+V����'��6���3tC��r�"�N;��k[�Ӧ��`��]������e9��)CUF�x���t���x�o�N�����ҷ�=�{AoA�w$�X�태���<E'*��/�w�p��I*;_&��~�̦��sި�Ϧ��-��:�j����:2+�<��'P��8�^ww�a�Ur;4B�r{08R0���>���<:<>v��r���ʸ7bXb�+(�j琦c��Ȳ�oX����"R�gwl�ģ.I����T�w��{�XH�����B��_G��|Q��c��L��ދ�\T����&�z\K�8B�̎��{�K/<i��e~}�1��o������3i�v]��Oh���ȹ,�7�(���1�&qS����Ț�g�<h�b��?W6Or7���2CY���Y��>ƕ#�P�QZ·��YG�K��.]����i���� ��peՃ�p��I�X���U��f��
5{{0�%*Yl	A�f/vw����4��F�-�ye}�� �.��e���]��r�'����A'����ݲ��{΅C��7	�������+��F�.,�X��U+��a�jL1��*����v2�2P[W��)E�!�E� ܻX���_�/_xx�|�6_� 6�Y�qw���v�{{�;:Z?�X1��bH���Q�-�mnn\\v3[�ݺ�x�;�s�w���Lnh�=\����v��s��y�(b��������k;]���mmE�H��q��;vD\�3ۅz:7<am;��]�zNN٠�7n��q�6��̃���9�T9�B�=L9�d����3�u��ϫ';�<.���9-V�EWmu���*v6���.�v�CcV��`2n��[�u�����۴\�������NG�#�k�7���Ō����r�VL� ݚ�ڛ��ˋ�ݼ � ��1Iu����5M��mC�z�̼ۛvzE:�a&K=氐��#/�b#��'c9w�θ��'���<�/Lc=��s�uO>���rZIǋ�)��gZy�v݂��M<λq�뗐�v�Q���>Ŗ��m[��x�k���6qv���GX�[O��6w7Hlu/ ��C׍R�ig�d��t�ckЛyunz����e㷭�</a�;�8��vָN.ջS�j��2�A�e�xy���7�`u�ܽ<\�w��;����0i0�<<L��'b<��]����+�ٮ�s۾֩X��d��Z6�	:�q��z�G<�x�1�j�F^#�ԇb��;A����E�h�=��S�r��\0+O��C���Tz��Cͤ�牍kM��4��Q�x5�ر��M�}[�:�}g�]����7Y6KJ�Y��zS�lr��ף��\i*�v:x8�;L������;]��:����x��v��㳓�F5g�ö���')�.��n3���Yc�m����fxN,i��=A�P��#p��t��C6C�<jݱv��G�=�vx�n�m��Ǜؕ6 Kʦ�!�ㇲ���W.��ڶ�����v��t�Vݗ���a���Qm���[E�\��|4���<��դ��6v�by�ƷN7�x�����Iɻ��8vU����u��8�����:���.�\���ܐ]:���/OYȆ���)ر�)��]�k�ώ�-pEh.��x���s��5v6g68@�6��v.vz�A�j�96���un.�8�KK]p�M�r���Gn݌:����� ���E��N�ok[zi���7��l;u�w��\[����Icb�Ɛvnz��ˋ/W��\Y��pS�e�s��Zl�z��Sx�Lv���v�� M��Ǎ�i��nx�ݣ��\K݋C5^}puF���͍��f��Z���b�\�����.'c��ػ\5)y�m����խ�61v�9�ݱۗ=�'P�DYŪᦕ.%�!
��F�~>�ŨK$�"Ƞe}�E5Y�e���S���1�8D�˹@�z���@���6U���j��@�_}6,�12$�&�7w翨:bPL�
�G�ֳ�b�ҋs�ϪpY��|`w���X����b�3��j�0���x,=]��.�5C%�O�`����v,,��k��ԉ��qd����ŶP"j�)mX��A�"|�������'2m(	 P��=��^��9<Z�����G����hτv;a|�� �����_yr����2�ln�DL��3,2Զ��2Ց��XU�ޜ��n������4N���A�C	;M�̎�ϵP�y5AYu�/>��39���v�����H�m�w��,�W���-�/8����E	 �z�C� XbO�X����,�U��qњ%�1+��$��ٱ�*c�qU��*w��=�i���<ا�=7����^*S[��r��I�:S\������nv]\�r��]#��E�m�뭨
� 1YE���j͵��M���woX�[ ��C�)�L���Vh�3�-ԏe�����	��G�Y��!a1�]p��g�`�E�!I �}���j�4RJRkk-e��7����\V��-ѢwbH�V���0Y�r�Il@'�gA�d�Wk���OxE�۹��OS�`�c�ɐv^=� ��s@옽�=�Tg^z>�h�u���<.��Ў�܇&��bG��
����
f�#B6Gx��j��;9�:�gW��=����|x�g�+/i�D(��i�V9�@�^��6G
���n;���I��Y�C��f`j�+� Z��{�v����U��� �!VD���Tt�3R$��}Eaⴏ��,K�����c8�j����Y�ܯY�,^�C�x^�-�`\��{l?��TP��#L���}n�7�^Ǣ�+���:i����i�FuG��4I�`���(�e��r�lU����dq�D#՛�ょ۲�[u�1�(��g���?
���b�,(]VCy�+�̝!�T��L���V4�s�6G���>�W��;�����v������h��%�q�p���㋐`mCn��۵���Lv'i{[X��Of⒈)B(l>�1C�	�^�Z4`Ċق,/��}鯮Ψ70�:!L�޺�C"�u{�>���r��܄�V��F���u����Z���-p�Z�YKh�Α���1ʌ�"���Tq�^��b����Q� �M��
�Qdf�E����V��$	���f(ϫ�t8�_s�^������jF���/(�+(JM����Dc%��!8����4���2�B6\:��|�Y�C;;�����
4K ���`�A���jo�t#�2s�&���k��(��8u�s9[z]e|�Ƙ'�q{n��Hv����䎑0�������TY����c����`���h��W?/e���lh�V���b���QճE�sCs��x��+�$iٞb�A����h�FR��*9i\��5���!ƾ��׹�U1S�P�9\x�W'�}l��Z��$	�u���{hCg
4_��4/�!�9�I&�u�jB��nM�[����1����P���B�9�e��,��|w�Ucvd!�L���E����	��:�,�TԴ�pk�X�#���m�nf�ic�؈kPve�:M�M�FZ��5h�}��i�4ͤ&���㎜1���j��}��0�j�)29m[!�#���s��F�׵m��/���ŗ�+��;v���A�H�56Ӌk_{�h�9���y��>t�,33�퍬�;�3ӆ߻<Oo�3d|����_�Uq&|�#�~�P��9����'�~y p��p���/~��Q�)>9��@c�>�lvt�a�A2�,�-�7�2(�^����U^��ƞ"̑�ȳ� ��N�7��!��R>����ay�
7{D����"B�t�_�*��Q"��T�\����\��A��h�`Nc��2c}4۵H����Ј����݌���OLYz�����zY6��������p���zb�_V���|D��&G���� t=j@�6i�j����Nz�����2έ���ʳ��K�03D��9�:����*����麶a]�Ɋg�����Z� ��0��=������cV�&����F��8t���g�k���Q1�a��S��|]]ث'�D�C��MI���Ƈ�K���̓ �����D�l�(��g�kI��_�g���kn��1��=l����6i�Xƻ,S�7�����ɣm
Ec�ZT8��@6��拧��Ċ!_}udm8�M/V}��2��=�$�A��Ӗ*�T�m�4����j��#�bcY�^�7;ޡ �������*�7��E�e��"�2�H��'���?�����|e��#��$j����n�O(�i���t��gΆA�@�L%���E�3�3������le$jrKD���g��%SEd�N�6�rz��}�Q�U�I;ۡ���&(D�����d���(�(�F�v
F	��{E��j%e}¬͍�E���Z���;�zG����&�Q��|�m�Y�[C+�hU��G��0kNF���f���賩��.A�O� ���U��RI�T\�*�C{��Ɲ"̌C�+�^#~���YW�Ǐo��*]zYko�_Q
��K2�rظ�ne$G��h~��U�8-F	&�?]���1�.��8r�duǐ�ᡟ^[��PF�/�ț\��;��w(F��i`���ˋ+'��JF���eܺ�q+�bߢ���9~M�����x��3��}��X=2e5���ˑ�V�>C1oKA��N�HG$EPnѶǷn0F�G
HvNțz��h��r#)���n���ۥyb̓cq�瓞l��sθ�ۑw��7^�hˀ���!��b�N��&�sc�a7��1��gֶ�t�;��ɷ#v��b�x�/�]m�k��]��g���b����km���f�b���&�;�݂�i-�=v�uh���j��8�f�/!�0keC��5m�4S)ծ��Z�Lk�n{���&�c�a���gf+��.�n2�uM�/u��t��1���TG��@�>����q�f7���pb&����$Kˉo�4:��3�߾Lo�2'�#�$M�y[��|��$�C�G�60|5���	���%�X4�
�w)�\}�k���(�*Ԙ���9Wٷ�bVs�ϝa�Q`�<Y�j�c�e蠖L7r0j�֘H�u��XG�����'0�9��"��|����,+	m�{[kXc\v�H8Qq���Ō>;�|�#�[�FY$^k�2�}^a�*�=�Y���t�|����-&��+}�s�"���\]h&�i٧>��N$� �A�q�VD�a�^�}����4�x+	��Y�CZ�z׳+�#�<Ƒ'�a��'��4*1i��������߯�bw��ִ���~q��0�~���cW�_-��W!\m�RJ����ܞ:Q?�!�}|�H<�َ"�|~"���F��?[�B��8jMO>��D����c�H��f[+����ռ*B!_�G.di��f�L� �����),AN�ۧ<F�+Ә^�ǵ��m�+�qB��f�+z��b�̣n����}�ߜ���8��:a�d/��5`��&���B,J�=������(L ��3��EYϫ�(�]�p�ڤo!v����Yw�]u�:֞2��7��B�`&����i٠N��'���|�I$r�dx?{�LM�ف���
�ݍ��8�c��''�A� ž:���g��ִ1�	V��!�ƽ�x4�l<6X�w�|G�$*J����l�nW�fB�Ϧ��[<P&Rs#�,N�W݆��� s��sbHex]^O�2��e����g�!
�Df X��Z�c�v
+T�����C��(Yg�Y����f�tx��5�w(xx�=������o���Z���9֚�\�=��ʛu�.���T��	rT�,i���Q�.�t�y�Dh�{7�8����� ���
��b�:G|��h�۶(^ ��6�#��dfc���/�}^�E?�lǅ<�#N��_}��Ԭ��N�X�=��yr?5�=Lad��_��_&E���q��=1'��U�㊻�0�5D����$j��Hq���kN �Lu/�/�yw��̯wZ���*i���ښtT����K��N;u�������
;d�7!��UO+TuP�*�
��^ۙk�kMLw����<C�.��&��
�B�qe��q#X�ϸ�|hS�vJ�Hc<G�X"l�g_���F#�"��$f���۶ێ�v*���;4������{��
��c�R�f�Y��������W7�4'��N(�'+�ۆ�U�D�pX:��G���V�Q�$Q��N�N����N��_$˖��d6�Kd��'M�L����;�~W���c�il!����Q�(�{ʼW�p�[��7�l3J��7R-�i���n\};�����qg����Rx���{Ց��r��?��#|}a��%�v�i��X�����&��}���V�1����^���SvIE\����qp���+}�:�J��y �^�:r��̟�_h��"m#��TC����è��"�+��#rj̕᠉K3Q'>>���QmH��Yj�Ϥ�������(�{��i�8Ր���ߞ<tya��H��8b�L3�c~��AfLQpx��!�}4,"����عdO��5�q��>��d�I�g�m�շ��N���
�@�j�h��x+Iv���v��'���t�<\zl��̔���e�T���^�O.4���S��s|���dW!CT�&�x��j,�#�
��,Re��kOb���"}q(�D�\D�ϳ��Bx��df*C������Z"�Piq����׼5�����ӂ�����r��b�d�-��q"ٸn��!������v�$�|G�P�_h���X�� �ϧ�,����y?��-�+���n��4�������c�N�'��!��U��T���c�छH�Y��![�F�ۜ��}��)�bB��$�#��kb�Zy�]u����祙�L �,����,�!���̘�@����Ь�8��������9a.1�}~���|�&�kL�7O|o~7g�,�h�C��&����,
��F��VD>SO��(�>�\�7sH�,�iS��w���5,��/.�:��Q�����,V؋���z���C�@�2�{������t$,,uZ+@�:�����Lߊ�q����1��?X"����uC\w�d�`�Ѵԍ��4"��>�P�a��Q�((�^�y�6b��P4J� b���vA@��ݖ�d7-�m�St���GY@���M��1Z��DtQ�&���..�C�̓��E�����,K�Ǫt���ϫ5Б�dI��5F09�ϝ���kdQ�|fOX�0�I��$F��ܤuD�D�*��X��S�X!��)L���q�fr��N$Xī熅�Y�2@ҵe��P���w��E��O�P>#�q����QX(��m�{����DLh��5���s�h��,q��ni>����E���E��֖�l�zk�m<x�6ar�e���^Ѭ25Ef�%���نCFe��vN�#��C�2�_}�j��采$i�+�Um�~�� aJ�D#���ߧ��F{ex���aGw�<s�1��J�����CG��A���B�p5���ɰJ� d���.wգC�]��䪴T�9�5���j�ݭ|��4RIEBB�K����h]�Me��0���64�]д��6p�>I���oA���M���0�?�Ŕ�?{>�`�.�,�H>H�H$�����:F���,L�
�>�X3e��e�Yۗ��QX�������X��Aݚz�Hڣ��o�|[�Ôm�cU�Z�ߨ�h����.�*��.dQ=��v�wu�Nh�B��;;aݞ3�it��r���{hϴ�;��e�j���5��.�n�G�6��6y�gE%n��E������v�`��wn9}��Ր콶�v�9Y<�`@�[f83�ռ����6�	ՕYN,qV��qq���o���y|�m��Ұu͞�ù��e�'<<�y��v+���y�8���h�k�F�]�	�ijI�\j�랏p[�A�}��";)b�$�c���I�X8�!ۍ{g�{eD�/km�qɜ^[�ʑZV��f��l��:8���Q��8��3yu�݂uQ�eA��I��B}���,yA��,�Mn_����߯�B�"G��fw�E֢7q�a1�^O�UIkU�2��ƞ#fl�4h�+��}hg�T���ĉ6<���<(}�(���6�ϋߍ¹!d�Y��}�.@+�Ft����9��΄6ffc���@�^_$93co�U�>)�}f�N�h�1�� ��T8��eYſ|.3�ga��4Dc^H�$�A)p�}���G3��8�Ʀ�<���P��F��-�������j���$i�2���`,"�v}!��#>���4�l��Ȼ�"�﮴��H�-"Bk�^.n>��4��ǌ��z-�11g�G:�q�*�d�L�<k��H�A]	;�l��Ri �^`�c}�8�/T�Ŏ��L1��e��D�u��C�Bu���5�\����H�y I���vs����o����Ի��e�u)����d�6����fs=1�;n]�1Oa���1)��D�#0�ZFEo���`bV�FH�c�VKS�ZFoD�*��C>�V+&��$�c�.���%q�G�N���
�{e�&���'���|�����f��c�Գ�2>�אX���I�i�7��e�*��Lm�P�t(��ɨبC01��uE���J1�ʴ;p��nFRuGz���}fOb�/|N�0)"()��^���{�,B���A�q�� +_c��}1jW1�B�>H���u|>"W(
�̏��"��	�|d쑤�Ye+�G��ȳ�ȸ�֚�]����c�X���D�?O�V���ɻ7�&�E!��$d�9b��r>���T��%�G$g,4#2Y���P��#�$=I�8�h�s)�i��x-�������ⷖs�>���\�=�O��7��t7� �!�fH��]��� Α�I⍕�=�n+W�M��$(���t��ip�C�P�Z˗�m���0�"A���|���VW&(Ic����S
�<X\�8�G�>�a9�Y@�6Ԯ�3vbҪ����}���&��CR$��c�_Ɔ�A����rY�f;���#PFx��C�c[i�[Χ�_NUx2a��0��6�����s<�Da(��nJ-��]�Ӌ���8�ji`�䪈�yu?=���&g*��_5h�BRub��yVvQ'PD�F�(�y�M}q�Ds�d�̀er �������X4���4�pzP뿸V�w:�ԭ>��?��#lHo��8�pMII%��.�6��o-�j5*zqُ��x�v8��1���A�r4�!�^ۻ$H\Yt��/K�^�֓�6ظ�1��;�G���&�$��xz{}Ou�˾1����+����PmW0̩IKX0��)銑ef��NXӈ�<����8�Moٝ���!6�.�CD��j({ЫtR��T�٨j���h��˃b������b<�3��Y�	��i�^:�����J��j�Ǖ���دO\���8�:.���]�t�|76��w!�����P�ݛ���%̤�q惢1wP��f��gpZ	`E�9��|I����s�� ����$�W���t�{W����.�F������\��?��z���޳��a����"��ee�S���Wo�d�f0��C:h�$�i��h�l\FD�q�;PU�����:��.�0�֠{�z�̂iW�p�}ɩrx�&����!�!��e�{�����Q�B�l��t%�[���Ȳ�*�.=��j\qo��%s��`9�ͧ4�c}�]�H�~ʷ��piѣR� �|�O³�j�Ƕ�Wx��Nz������:J(�Ь�Rw
��	�x���X��Mg����=��󻣧rn)���J2�W��]
=�����K������{�eB75�0~ޗ�F�ط����u�ڷ������O�f���sT�+�*5�T��&�V�ܻ�~�_!?^{����^uJRz^�R�
�������Ր�]��H��}�?�S|��S�����;+'��vw<K��C�{[���=粆�|��FG�4Im��ow�%��]�wwx��5}u��P��}�J�������*{�m:��;���J�N�ݚxP	�="�*T�+�&�N�Aix�e���w|����o5���[��f�"��"�bu���o��9�~4h2�Z��U��29��M��.��I����X|QfiY��~���@��&0Ui�DcErD�ٚ�/�Lљ�<��"v��=�+V�8���ӱp����vM�Ihm83�#��@���=���RG��[pJ�W��.nT���j㌓n7R�{>��8 vZ�%�����v��$ƥ��QDN�K�Տb�4����>5ă���čA_!���m<�d/��PC��!a_}ΰ8�sd�⦅�spmm���>>����V)V�GV�vN.4^�n�9؆ ����HG8�rr�^ǋ����2��i���@`Ih��ֳ�k�~0��Bc�϶la�qG��V& �+>�5Q��m(��tUc@w�6*;}�mƐ����}i�jB�A�?V|n��q���hWmIQ>�s��%��tfQM��;h��Bm# ϳ�w��
�r�x�s�<"�8����y|��\i�,���#�}]��r�H5`���\��u��M��_q�|�{�*��C������LK�KBX��%�'�9�ȓ_\d��� '���$q[%M���D��D�w��htřO{Sݓ��R��+>5��W��`��3���=�L��P��M�g��$̲���G[(gM���}:�׷�q��N�#����>J��&8)ata}��M8���"�fA���j�"p`���O��#�N��&%�U�\���s�z�g,j^��I,-!`��l��6{:Bz�k&����w���J�`w;����>�/��V��D�Fɕ2�U/}��MҕZ�T���C�c
���Dϰ^�n8����AL�IŶ3�/z��vF��{o��9Ebt��>)� ��>u`�K��.��"f:��H���7�#���8��_گ/c}��nn,�۲Ik�Cdm�}l���]%y!���s������xP ���x�V@���~����D�ǞR�m!V}�6/RAd���l�7q�?f��� l�������0_�*	ՙ��:�=��L��C�+~5$qΑƀycU(����'��75���S�����hL����۠���}?v��'2�S�{�tՂ�!&���򅎁l���ؼ�ԙ�@qL�
rd�3��������S;y�mk���Y2 5����|2 ��+� �ߢ�ON�OZ���,��Y#V E���$a��'=��4<p^�2Qq0+�'F�C	ѦE�:�X��I6�I҉6��m��;�{o�*��JE�f��V�gʧJM9���:���綉!���u�_}��f�z~�2�
 ��D)��P�d,�0.�w��+�Nt'�$�Գ�wwkŀ����'(���nS��7K�KW��l�Y���ʫ�͑;W}��ꋿ=���%.۠����l�Ә�r���st�!N�-���Q�ץ;�����>�kV�on�B�� 0�$����M�Ŝ3�Bq1O��G�5��ҭ�f	NpJ� /��'���5�}}��-Ж�=c#Z�f��g�9����t�%�D��^NG[`�iy�4(�0�;t�q�]nxx�P�l��5ү=��c[n<�˱�E�۩��f�7=�v�X�ՙ�f�;a�Wof�:8�^{v��V{c��l�р�gZ���[��zm�ڭý��썧����T�S��a]��o9�KE�k���l,�Z?���>�>{c�x1X��������|��k�\["�fu�k�s9����&���nL,	n{<8�v�z9��h�kv�ﴢ������Ŝq�zhӋ�Ÿ�y�b�5ᨨ���NxԼ8
��`�b�QgNM{-J�5.����+-�[`��ǵ��VZGP��^
̪����s����X�D���5�S�(����d�!�#7��_\w|N h&%=�w;
%�����%��-(�L���˪n�{V���<E�r�����*���L/Nr�� Y��3u��/LaƆ���o]YU���H�J����</^P��R�Ɯ��P��x�v����GG�=7́F�H��ְ���|/�*Ek��.	�"�BBR_<��wNt��{��9��UZ�_z������
�6��	$$+377[�u�'��E��7�p{�S���
��Ȑ'���cH��E�&�@�0�罳^��
)�j�eF��3��-9g�*�b�-nԖ�g�nr���fݎ�8P�uv��7gqs�M۞��u֒ �ZJWX��s���ƥ?`˰L�11�dc��R����H�"�ċ��:�{8/��	��1��v<� 1F����eÐ����&5���j�k�Ͻs�r�0�m��r?����FYM��扇	�sʽ{��%�������h�׽�{e�����W�Cҋ�S�O*�}V7D�t�1�A ���V1  [A�{E�9�j��"�0ȅ��N]�F��������׶���i�bI�`nB�DS�+���d��J&$�����N�e���9X��U|>V�$�f;�BA�1#J�Q�]��,i�K�55���3KE"����.v֒�W&7kL`:04�f
V�f*S5<�cr�d[d
�c�G<n,<@��#�kA]�2�רڟy��oq�=~!��Uئ4�Ҹ�����)#�c��q�=�&�B}5����֌w��mn�-.#@(D�bufPsY��a�c����LL��1��i�{=��mYU�� ��:)㱱q�nM��*1��)ϋ�[۞����ӝ��IĨm�J�%�kޛ��Naw�;�Ɯl�͑t��_��(��&@S��5Q.*t������M%#�wa0�a�6jbmD�#�:�J"䆛�;wa�L�)����^�R���whX5q���9]����fZ��t�.@�%@6@8�"�ԑ�HMi�u T�&%�%O�!K)7.[�3(��F���p*ȓ����ދ�cd
�_�,����z�lO)z=v]�EҖ^�"��NYd_cĶ6;/�zL��_:����rs��
����]���Xd�O&dk��:�evɾfr�?�^ڼ��f#��YS~�1����mԼ��-�4���e+W�L9m�p# э�v�Ht�8�OJ�����X$!D!혋p��x��E[�>�͈�2����06h�'哙"GV5}��v>�܈@bٓ&4�QB�����ԀG-
K�x�j�(��@N��N�`H�DΑdY��)����װ
�ꨡ�/�]P��~ј0Ũ�,�� �HX�ƅF!�"�f���Κ�z���b��n��U�5H��=knŸJ=Zo�rܹ��]�.�]��:�ƱɁ�H$Z�[b��[�k�/]�`d�ͮu�TT�!LS��7@� ��T�H��
���)~��� �P7n�f�n�P.cf*aDR}S�"T��@�]���J�yi�wǸ��-oMS�<z�[���ƹ�!�:�QCDŕ��!"��\"�Z�*"���"�(�e	��r�+=��03f.���VA2��I(�C)u���������s�:�q� ф	�Fҋ0� �e�&䁸"ͼ�G{Gyo�Ј �Z��Ϣ`Q��� I����3�k�*��G��K��9��X� K�r�7�p7-XfRE�^ȿ`�����cq
���UW��ndL1sD	DVy�`�c��19��sP���އ.?�8�d�zg���	�ZS�ZJ��4gV���q��2'd��J�ˈ�JuGd{�
���-q��/��wz��o`� � �&E��S=^�F�	T+��]x�N�GK"L(��~�B2��d	aa���W(����ѹ���Db���q�n!	f%ϰ1f�ȑ ��H��9�Y��&0(�d(��JĊK�n˻qaz�n�f��ϋ;�#U�\^��'��=�ĢZ�%���N��4ژͥ�m�1�%�d`(f�L�sΣ�&t�gH��`(�N١6bu�N!E>���C��猚	��"b�U^�TV���[���*O:]߽�uR�\�ذ,�D\��VB�?`���9�Y72=xٸ��Yh����X���!�`]y�H� X@�p& �@8D]�������=۴t���;�]�%����jȯ
QFV�(�Y�\�dĐ�Q ��=��sc�u(���}�����C�E*��PH�>��"�D�����
B ��T������L(�ً�aE��c����h����Kk��V5��>x�I)Mx��a��^(z���YpH���y�ÖL%��t��"`�!G�9f��Y��6f�$�Ef.hh��ҴY1�h#\ 0�'pxO����X!��Y�.Yx��1�{4TY�1
(���]��M����t_��P��(��h��Y�V"WK�ix�	&�_���4�a@3HaKQ��Ch5M������[����{N���0�(;�̊�5Z��iW5�V���7A%=#A�h��h��ȗ�=�ʺ�W�U����GH\�E� ��p��%��@��#�=A`�fr�[d�j���eoh�ƛ�k�����z �v�nt�[]�w-�G�ӄ�ar;<��ϐι<�Z�]�!E	�c�z9���;q\�\m{P7��f),�/Y�v��3���i�f��q����3���`����S�����vy^ݱxRt� ��j��m)��5v�+��r��hLÁ�EĻm�jLf��[Xyw���(�3ع�����.�5˽9�]õ4�rs^�M��E)o��1$��H1d �*�CK�4��e{�B�t�dC�cH"����E���R	 �!��2�B��F��e�4�$� i@2�M�\.�����p,��Py��Z�#&0�ʀ a :[�Q��jQNتp̀K@3 ��~up�)E��@"6��y�d"
7 c� ��7�hHFC%����,�:��"\{�^���n�	��@�y�:c HY s���2$�*_�P�x�qdF�I1f"	0=���D3"�D�t�ϼ���G����� Vr�n��!Y�J�hdQ�@QH�ZF"S�-�'�4��P�Y&��E'[��D\A��s��e�H
��	�y�5t� #�&)�� ��~�Їp�za�!�� !e˧TO��U�")�Y��1�"�@ͨ�Ha!D���s.H�LJa9lTi KX�H�0�6B�?��QF�$E��2�)�c���O�Dh���H� q��2�ӠH�`T�� �W�� j�D�K� H��)�evmz�%�SKe(�'`N�~������A��\=x���"� nݷ[�Y��ݵ�aL�	�ʲ����a�a��s���D��b;�0�,��
H�#�@5�B�x�Q`$�0/�N��<��(d��z�\��@�$E������ƃ�<a��<DV�E�&0�PMa�BZe�$��M���@$�6B0h���Ð+��ug�2��Y3�P{�{�W�ח�����[��٨�Va�h��*�媦 B�m��ь����l9ۙ��5�[��-��q����D8`�f��Y��X�Qu�D�"�;ӖP�܌7@ (����McH�����
[2o��2A0H�@Z``U9%�d`8�&R޵q��lJ��m& ǟ��@�0	""AI@��"@0);��b�j$ڿ{l������,�@�@ �^�`PH�a��1@
	����-�2��E`�n�i�l��mFR�o��f(�/]����07���ʿMb	LE�&0*`"x�^�j�Aa�(®}�[`���Lݐ#w���F��LE�L2�xyX��i�,�lTa�@� d�� �g�@��3�P$B0�CԶkln]]�\C��M9]���
��! �[�P,A1�y�h	��0$F(=�j��������Q��D�e�o[cZA�f�d�X��x����F�G���<]��#����/!�۫qOJtn��TJ0V�+��X�K�j6��:(���E��>�Qb�A(@�P�� a��L`{�|(q�@dI�i��B�Mg� �3�#x�eV�s0���Y0|��1t���4����0$�S	����0��aQ@��4�D�Dh���:4�r�܃y�ؾ��p� h$��`%ٕj�c��c&a\�F�{�QRH�f@J�H����{ ��b:b[��<��o}� 3��8�H�����jD�9$�-��ZX�X�Lx��J&�3���H��b�� a�Lj�LY�ƘG��p���U�)�S|��|�{H����/�'ŧ�1������N�+���8��Iz��b]���81���[���O�d�I�U�������@�$������H�b(���@Q;^�j q�8�&��8״<�8GF))m�2�0�b	�@Q g�L�Ί�ѽ�=5�&)Ks�@00	�#�$�10��֪�H��b.TE=�,A�0��QDʳڨ�n�	7U��QD ��P�Y�d$��	3��{�R�D
�跄��8�Ɯ�I�(�D@���#�� Hd20��dCʭ*v��r�w�)����  IDi�RG{��@���F�e!���Q��ikM,q�\<c/	V�ڈs��+�-��h�����R�X��m�4��n+v�!�:��0r��h�D"uL���J�Z�o�M�@г ����B��8(�D����D'~5�1��2"��4��
 }G�*��.�^��qF"#LGJ0@� ��� �(2@�0&ڙ�dB�{�ᕁ�e�)����� d'�0�Ceb,����3��T��y!����Dq	"0� IC�O�j"��`i (&"_�PDa�#LE {޽�BP�L��&��wN�{��+��bZi`["�Zd�ѹ�3,�,P�@F�Fd��x��"�@�Y�i���Ӊ@�C E�z�� ���ؼ�&�]����
 .�c�DY��"&��DH00���ڵQD�"��c�$��xQ̋޼��cPM��.��ǎj6"�m�;Y�:�����`�b����f" � 
 	!��٢�F(�TDY�Dq�"#�� Y��1F�ȁDCf�_���mR�;bok}���$(d�'��KI9�A�u�$�(qu�:K��ĵf�R5�h�nv�ho�g���}{K�]�J����q�]�@q�@� ",� �~�ǴX� �������a�� H0/��t"8�p�,�FN� F5#^&l���@I�*����@`G Y [�MW1� �D����4����@f"4�(�B i��w[��5�v|&��(�,�f뮭M�뙠L��\�q�#p�b��l�a�س��u�F�D�#�Pk	-�,	cH�1����"0�f  F� 
"���K<j q��1�� `F�<�@��yx��L�Α���1 W�먁� 
" �2"�J�<K�Z��[R�@�� 	"a�� 8� i��Q���32f���� E�.1M�������s�k��S�K|�׭���Y���&�'�97��D@& �
�x�/����$�b � @�*�R�-7)�jY���1 QF""H�� $ ���" �"� 1�D��t � E#d��kj � I�D?_�P��� @dg5HG�6��]��*��'F�U��^}S�8�`��P�K�I!�k*��;�+ˡ���P��ĵŶ$�
��S�����*�(o�:�[��ߍ���9�7�� ��,�՚$�����P1 q��� @F0 ��X��2L��%�庁b Q�,���1 wg�T@�&	 3Z�P�/��͹�������J��}��\���  ���� U� U_���U} U_0
�� �������_�$��(� ���U� ���V�
�����U_P
��U|�*��U������PVI��c�� b2` ���������\�(��-�m�d�@іڶ�֊Ͷ5P֤�V��!� %k
�Y����ݬ�m�MehȤ�gB��6�*�E�*����k�aT�J_    z (   
        @      �  ( �@  � ��    (  P 'Uﻪ��7��lx��lͫMu��.��8��x���[��s�E⎍=:��wo]^�������N�v�J+��E*�\� .������`�M�f�٧��4RT��  /0    ��@     u� p      {0 =�  m�E哳^;��=:�ۇ��osT�Ï ������p�{mc�b�[��֔���m뻻�֖���
�����)�   �  
  z��t�1��ڗmfm��	��ye�����W��i��{�x �{,�\^�����+V�x�v���v�����v�Q��Z���׮��r��^J�k�m�e�sm֙<�]h�����W1��9�/[f�b�Ӷ�G�� <��vժ��W^�;�=����7;6�3ݯ/WaF���ռ��M���$�m6緧��0��̴��@��J���         ���n�u�g�)zOq�-'����Z�^vWE��p��<�y��cs۽i�y9҈�ˮm�Y. �/z���7��MRW&v�S6a5��Ui�;��6��{���v���ў�Ҥ�:��k\�={�S��sl�����m� ]��j�w�ݕK�<ڧh�۞�Kҭ��Ӧ���A�@(   P   ��6��{�Q[[k���Y��������i�mk� =��Dk�9:��;��5��y���"p3��� wWM��w]3e�����b���%��v�����{��1� �Uv̶ܵ��y�^�ն��ki�{�7<*t� ����^��<m[m��z���c�o^��#Mj�����     (P �{Z�oy���u.ղ��m���-�M[\� 3�k2{�<^�Z��Y�r�-�cN�6� �]W�y����R��'()B��F�9�v�5����kc� �y�ޝ�f�-{��:)O!��޳�����#�]�1������Eǈ��Uk��^h:����i���5�n�������7�(J(
�)�"eJT   E?!�)U  MT�z���y@ i�تT�IF��� ��A5JJ�F L%="��z��a ��o��m�y�Է\�F��Y�	�Y�.{�<ѻ��	����9��=�J(4��e�(���QD.袃�(��PbQUEU�Ǿ�������ї��ui�I��_{�7��۾�54j�&��ycx!�Y��wB�3UK�&���'ۭ�p9����V[V���$��0\��Z\�7i8Q����r��������+�ER�i���]]�c�qN�u����J�\71E�W);���,ݩ�Z��s��Q��y�z�%�-�z�����S�9����Ǩ�s��K���ޘ_S�kϵ�g5[�`m�golW
�nP�|8����4��J��W)ôrU��jR���A���`��n�˪���fZ|�*am��I��/�`k���r�|~�3�q��ج���k൹IJ�T�h�e�V�4�oٹo/7%o�Q��V �y��P�P }G�:�` �[{h>cF:����S��P�q͐��2��ְ��S���U5�U�bŉۘr�"��v���n[�J�ͪv�6�=�ƒ~��̄!Q�W,�ݨȴZx.��8i�y��'wZې��침j�Z��o+b��h���xC�X-�W�pQϴ(c:���
 &%U5����S#iB*�#�F/�n�J4e�*�8ݟ���q]D�AYr�bf�o�Tu1��V��6�
�Hkqލnl2�0�v0�v���!u�-]�N���f���;"Z!��SZ*��������lMͻ�׹nC9�I���CO[�u"�P�ҁ��-o^��^M�
�Yی���j�n9G2��{��vǯi9l���1uvt)�LSJ�xO�ddR�^���D��)K̳nݯ4b*�5�;t�f�������g�Avc̈�"���16
�(.�Sـ5��o����4��*�Q�c=�m���;�y�{Z���kw��vKF,X��aMے����9t7�]@\�Hhʦ����G��]�3��LK��\N!V���fH��q^�� ��
����&��*��p�b�]��05�-�&bf�ֲ��&)���n��t�ݹ�N�8�B�>���;%G�;�/"��!ʽ�B��)SE��;�_;�oRd���l�e��+U
�����b�<�칄e)P]���t 	��N�;9�\d�b�`����I�2��R�4[A�o�	�Y�Lx�K��h.l���X>��Q�b��ҍh�k[�
�,���3U]��W.�!S.�<W�*�īHJ:+h wS���j��\o��:vy�4�ǘ��Ռ��f���`���)�\l9��ug]�h:�l��sL��2�I��e�q�K2���šV���N��+ �4h26�2���1Y���Y�Z �0���E��]��<Y2�8��˅P���NN�ntqݫ�n��u�B$r�޼f\fйB	��,�3��˘.����fԓrV��qZ1��-���D��56�R�
)豰J��b@��fk��t����Bj&�C[��!`!�,��U��X���
��E�y���V�];"SgE)�rf�ܵ�k�c�	i�y���ȁ;�W�dmc�ʄi5�ź�35�r�ttn�apa�l�m*�SCǕ�t�����gĠҼT�߶MGV��ŷ5�˫v�
'b
m�s#ɦ�j��YPV��,[��ا���/cA�r�56�Kμ؈��;o�ڼ��ap5%՛��4�����,wP;��~�`#���w4�aK;��6��r�Q�)�����m囍V͗E�Q��_^G/'���1�QS��JȲ̘)cK��ԻE�Ǫ����W�Rf��,L����u�̡��l�oND�P4#٢:����,oRt�l�eX9�x��4���o{�;�*��s�ɹ�n��ڎŜ�܏tCiВ�;����#Rn+�bQ��Fv�h'C�S��,�;zB�&�h�U*S���M�W��Ehe��޲Љٟ*6%�Tm��v���E�x��(�"RQj�Ea[�o�b��y�_SYQ������P����B���)��cҲz'l�Oޡ��U	p�W��L.��2ɫтL���*M_d�t������؍Q�L÷&��,T߲?�n�а%�xA�)V05���%޺�!�TH'1�k\��������׮��4tW�������g�!���5���M�8�F�^�Cɏl��bū̶�`���Y
.iEL��Ed�CP�KiF��|6�w��Lc\8�kk�*���ek�]�t���͛�1)6k�7��qP'+#)��6�l�"ͺ��髰�йGv�kf�C�)����[�:\����R���Si�BR]�K$�&�M��#vFKWJR�gJ[�/m���7G��O�,\K�*���>��h`؀X$A3,���vU���$*�cV�5Z�t�p�
�0P�YX��ԆD%�Z�Ȱ�B���N�rfB����9W��wL.�Ƌ)0��Z-+7d��F�������Rɣ\�k
�:�8���l8û���:��Y{���ת ����O�5����3���L��[��ŕ�0d���Z/R�8���-E�l�汊���TBi��D!u�+v[�J� M�[�i)� �R[S�;4ʗ��&�e�I�u��Id�P�L��K��d��6vMF�ڕs^aNỐ�V���IH����Z�S�U�+^�8�ԕ��UVI�6!�p��n-�v�f)�tJ��{�0�Sw�<����Yw�e���C�Z��S���ֺ���I*�	fe�K�5-���m���y����׎�ڡ�Yh������,JQQ�I��f���#^����9p�_5$�r�6+��V��#P�g��L*����ɴ��nn�L��Z�{�6^0�
V1c��6z�3aR����2m4�KtiaӇ-�X�r��$��/EZ�1@E+"��l/�d��W5ꖘ���͹���&���o�j��ANP�y�	F�5��a�F�RhV�Yn�]��2~
���Ƀo[Y1k�i�2۽����kk2�6��_^[�L���Hz�	|ʽ��H��Hc�f02�U왚d`�(8�6�;�lD��L�76ZZ��9t6���keiv��HjT%TC�Nˈ�Zt^��B:µ�hc8\�K�Rh2�mSHn%�Y��Z/ъ�Σ�ˤ	lK�P嬥Sɜ�Be�@Tq<�7t��'փ4ST��*8뾣ki����[���ŃJE%]����<�����Y����cn�˴��X�c��0�Nj��I��g#�pvsv�S�43����o2VB��A�(�1�@���fec�Hq�zu!S�Α�2��Eѧ�2�ɤ�� ճ��I	ye���C�aR��jB�ӕf�UeY
�ڮ�_R�KJD_S�F
9]Rd�j�ߞ<�rY`�d]]�JB�8F��9eU�Z�Q����J\��k�WY��25��Rku�YX�5�ض.��&�m*�Ӫ�3��܋]K%کN6b#3@uvh��ƭ��-��V��u�~���O��>!k>~kkNM�A�������mGi�!S�[*ؑ�tձMA1��v��Z{����P3v�]cvS�c��P;bꯕ.U��>�e��t�ߩvH��س8Vm<��l�S_�{�r���Zs0�y�)�L[�"ۊj�h��H�*�Җ�M�}[�E +>r�ԇ�{-����_���U��)Ej�Y��e�\��-�RCBf�E5j�H�`�[�2�ABW�M�zY	!nj�F]ȍefX�U2
ˮK&���y r��|�n�;UU[��d?V��+�ҕ_��(��#�[�LQ��K����]�92�oێ�ڮY1T�]*�E��#6�UB��J�6�ޒa��d/_����$�|���*��Pk]�+#ɚ�<��~�o|���Tg�<[��n�U���)�<7bS О�	�i��8�ˌz6Q��W�(�A��>�_��q�OuJ��L+�a�oAcje��GdB��o�Q=E;e裚ӻa/-���<�|��W��b'��I0[��Ռ'=���e�=e(^Xf�KOʆ|,f �yk�nupUw]��c�۾��%�\�Ҟ�{>�34f�w��ݵ*�������ڕkS���/C]O�\��W`u[�B��<��Q�[�`�l
�\���b��ڛ�w[3-[BmJ�q��� i�.�P�Z*�6�@��iZ��u��o�,�mM�`���C>�-+FE����v�vŭ���Lܕqݜ;s�W�����StE3Q&�0�3^�1KN
ċ���ݵsr��-��K�5��w�2�*�Cwkn��i�&�!�\Y��|m�@̚��қ,c���yfZ��9so7C�v�dg���5qnQ�XA6j	S>/sw]���� ���34��3���=ͥ�@�Ӹ�ba��qA�K2����Q��F-hYU�.�&vs_T���_:��]K��:�Y`<�X�E_ڝ�Y7��vY����L�aU�
���[��q���nQ�#�s&lB���<�����
����6P�	ˊ�`��$�o��CF�x��y��J��S9X��b�*�i��"�$nQ��N�a-ɏM�L�A�~_QY�x!iK�DvB�@iE�hr��?Q�l<-��7x�<B�2��/�ђ�C^,I��@>tq8�f��f}��% ��C՞AL0b�q�M	١c�]����9v�r�-�We$� p{ef�m��p�jitU]���7 ]e;&� �f�Pc�7t�0)h�Y�C`ڙp��<TԲ6U`��R�wmQà�ߖ���rE��"�����N���R7A��>#E1K^��3��`Wm�gPP H��sh���e��R\eA����K�]�ڷq9Z��K"�M�aWd�Q������" �̺�]��(s���d]I&ŉ%��`\ʚp�c,�8H�q轶^T8:���Q�c1�3mD�&�ɔ��sZ�-p`�n��"�H�{���Q�t�fS4H�f�w~{��~�'�ҹ�fR!��<����Ә�U���Y�-�ɕ#S���F�?s*�﮳�G��ی�L�;��kQT�:�M��eݰ�~+(+����b
���Q��	�÷��3��M����36+�:i2ʭ[s��"���U��LU�����{{t���&�t�ᙻ��w�b��8�Ԏ�FSV�S��8������>��2��X�w��j�e͘��n��}�UV*�d\4�xf���D+G"����@�﶐��>B�FW*x�v�ꓥ�FϜz$�h�W�*�|�{���I�)�7=s��(�rϪ	��qUY��[�<~4�A?I'b���^����&��HVM�@u$�k{K����+OfW�r�ڨ+���Ͼ�i�h�ٮuA��J�Hu �Z�絪6�cGr��A��n̪��/����<DR�3֘���'��/n�+�u��J�\j����pGYSb�z�C�Q7���XbR1(���f���v�n������%��0�%ԑf=�L47fmU��s�Fȕ�m8*�S��Pʅ�F���+�h�g{Km��Jݳ��^{��c��L�^�K���D�*L��xr�#�h&�j�� �7�Е"ˑf��į��w�]�Hq<R� ����G1u���"����Q2}��W�e�Q��T�c�`�ۇVc,$0KHQm]Vj��t����wW$�Ȩ:�)GfX��~��qK��R��۔�xmH�2�=����Zv���1�u�bk��Z��勶-�zY��ֱY���m^��f�V�C19��aaO���)uk��LyQ�B�� ����Z�XWG4K�{ql��֭��4ۻU1�����*���-�d[�,�J���C4ʔ3q86��id!^����Ye?I �+u
�zK����[�  k��ƮT6��l*�*��h;ʭ�6�٧�v��gח6�k��7��2mix#
$�Ze�4�8�"�kz5��)���i���*��/�!��4^g�Ũ���E��37}���*?hFS֠��S���m��m5�cn��r�ꞷ��h�-	�j�KuZ�8;��[[$� �l .����˓�K 2�Y��P��g��Օ���2Z)m�odng��`����E�����غ~�
��B��5�cday[�׶��u��w���~��Z#�v4)�ED�3�l`�I[�K���]����;�����-Ͼ�p$��d��=�l_k#>�I]u�����R�߆�U�<&��4\�����p��A{"�@6��e��m�������+!���U����5j*u��M���n��nF�B�̮Ok��o��;{r���}�h��S][� 4;nq�R+,|!�>cJ^�	�U1U0k����e����f�'�% CWĕp8��h��M���L+3UJ�z���ra��͋!Ƽ ��Dk�b�:�hq�\�#� �j�Q�5l*HH27�ͤ�x#ݬ����˼v�� j���Y�8(IW2�nJdG�e;;B��3���V����B�ٴsL_��?}��
���מ	bP���*�lNә�����8���9C���ᰵ��(#�(⤙4-��-�gt��B!ɍ�v���r�M�1m����5[�t6�����zF�,O	�ׂ1۟Bn�$o�B�s28���B�2���哒�����n
���[��)�����jB�J��
8u�T��7�:�
g3n�������v6e��e��Nӽ�%:5�
Czk-ұr�)F��,2�����Z�)P�@ۭRG��2L63��3if����u���u`^��{� ǹ��	[��Q;���o3�	Ř��Q$�o���b\�����[��"�	�+�䖪ڽN�*���������*��Z�T��UC���
��4�j���]�
���[c�A�Z����*�&��c m,�J�@uUmJ��we����T6᪪�����
����m��j�������j����4E,AV5E��;iju�zw[Qڝ��^�Ul�UUUUuR�T�M�b,]T��k���|��$��R@sU[*�Dڐ���UڕjB���V�8QT�-[R��UUʵW�����V������UU���U��j�j�[j�V����j��Z��Xr�U*��k����Z���wuɱ�<�&몐�^��
��yۖ��k�.�(�(��&�ەj���A����&��[v��R R�U�,''u����:�k�O[��1p]p�X'�E��k��=���Y�^�\u�Dn���`uϷ[��`4������w<�Y��n��X1m�I�u=���뇱��q�{v�v�c���8익m��o)t�ܘ+�Ʌ��Ĳ��X�j퓨#��&�'�Swk�u��3�g�C�'�.e����]\�h�M���:��q�s�V9wmì����8V����m���;���r\��o\md�۫;vtɌ���r�t���v5�k����kˋq�>O5]�I�c��r�)�f[1OQ�g��=t�c���N�71��oE�.sy���&$-���&5w�#%���5���+׮�0$����v�΋Y'�=F����_�����]dM��r���wb��볹v<��c��K�;<v<o@�ԛdc���4m�t��;7�����8�s�!��s�n�9�[;�u�ݶ�}s>1ӻn=�Ox�ؗ�5���7h�Psn�ev�]����w�-Uy=���;s��a�ظ&���;u�-PnU�3N�����ȝ����r����x<�b�۴T�f]ѱ�nt��nph���h�������s��Z���?<<�V�F����d$�m��Nzٰ�-�j7�"�Ӏ޼>�z�g��sw*F�s�܄Ұ�nb��b,����by�Ty6�N.ѰTso�ƻ��z7u͌qg1HTw	����{L��5�y-���%��)��\�������휏ps�}v
�b�7k�2��t�%/6�0�CJ�iMA#ę�˷���ְ9�z_=����;�]�����ۇ�Ɋ�`;v!'qj�i�u�vSO]�n�Aڮ{v-vMu�\�2�F0Kq.Xݒ���kX�D쩵�KpLvI�⳻D�7&q=�j�v�Y����+��h���zn�m<s�㦗�nwT�[m����[��U��c��w7��YW����ZJ�"4����A`�N��^�lOC��ac=�v�\����.��<[��'c���{d�]��"�m����K��z�ad�;�r�y�|�[[�V�v�3���9v��ws����'�������EܹN3�N�����[�yu�e�N��Ț�;g�0�n[�mq��t�vp�{x�����.v���9n��y]��p�\V:��nն6�Ga���WlP��E�:�#��O�r?s~��N�v1I��n/[���N$�s��3ڋ��v��)��3���k�����l�e��[,�U�M[�����qq۫��z�r���`�뎑��Ls��VkM�q�f��T�s�f�����[�VзL�p���w��=�%���.��[gu1nFx�;c�+]���^�Wi#g�5��Gln�4�4�9��i��56��5��[mv��K�W��`��@]^�B9�q�sŞ��)`֎.�ܻ�;��;k��v�v+�e�Y��\�+W������y�ҷ��]�ű<���؊^�qZ�=X�"���Fx��m��m��v�Fz�+.��P����<s:��x�ҌWI۴�Q��Ė狳�xdl��Eȋ��ٍ��b�Iz=��vR�ƺ�bC��7����Jr�;����/'m���u�b��n�QMEݓ�a;6�T������vA�=�@�N�᳀e�W�r�W�[geu�{�+>6��.�q�Y�8�n�m��2�~����jlf�7k�5rY����n^1g�������m�����ӪNb��β�:�X�N���U۵Ӷ�J{5���kv|���S�ݛ<s�3��c].�s�Q��p�pg��a�{T��Q˸݈^��u��v�C�󷙗��`�(o��r��B�pt�3��ӎ݌n'u���,��`�=�{7Q�ZP;=�ofn��]��W�fn������K�!ܛ�F�q������"�gn�.�=n\�9�����n�v6��\N�5v�a��Y�����^ڰ5�;�#��m��wi`yis�p���b��h�<�l����66�ݞ�m�Q:��qj�&� �q/ȶ*^Ymļ�܃f!2���6��s�Og����n�Z�ň��/u��m�����sm���V�m��vn��(n;l�+�7[8װ���w%ΖG��;q1��d5tL�&�R4�Z�۠ձ�����^�ۮNڶ�\��s�'j��{�z���J��=ŶM�{{���kqhb�k]��wiv���b9���B[�3�@���v��]�ƴ;��QQ��AݚLu�l���ѝ���q�)�vquljy.ڻ�N�\\;�:g�wAZ�q�v�<�X�Ng<<��dn:}����	�����ll��k�n!{�vl��TA�7/�;�_�8�y������n��i�ګ��Dwg']Yj��12dI��aEw�p۔�a���a� �^����#��=Ziƭ"��;������y��s���)�1/�ꖬn[��k�\��H6s��΋ǷGI[&V�Y�)�N��/tdK�:r�D��3pstW����]�g���>�\�w���Ng��v�UZ���]N��ܱ�a���K8��x;n�"�G�Qy�ug�uv�;�;�6�nA�k���x�\k]<���Uhޟ`�����;g��܇N�{gm��\V�J�;	�QΆ�!�:xٗ���nطmob���q�g��7G:qu��ukK������OM��$J@W�T��z��oU���u�q������8؇<�&�1-ٌ�0��3�q��[P�J�<u��s�<r���2�YV�w>��h�f3���m�������v�۰�k����ʖ����n���a٣�ͅ3���z��\=J�c-�gqըj�Lg�MYE7���b�&�p���7dn�ak-��[�2���9J�leٷn��I�fcXA^ͻO1�>�
u�zq�c�t�m�8K��m'���n܏aU���K�0z�M�uΓ��V��!�7-��`�y�����Z��"���9�vX�GP��Q���ڼ�֮cc�u�^�{ F��Ba�jk�8M��kN3����r�nK�����1�{�������#]��X�v;<��������;m�
۞^��g�{t�Ļvw������\�A���mN9�Y��[tj֮HA�5��7<�<rv�N!S��]j�Js�C�r�.g���c5����MY���,�y��tR<�<ۑ��5	7�Uyz�ra]-b�X�v5�l����[Iɼ����T�. ��X;k�����۞�k��"m���r�El�-Ǆ�U�͵� ��d�k��]m�{7�:箯f#Xs��������N��3��T|��zsۍ9^۝%���numEY�\���V y��x��l�d�2�/@�R�AY��-��HzF�E�MFӶ3drtՑ�m�W����{:�.=s`���i����7�Ä�h�Ɩ-e��*: ޮ��v��1s/����0@s9�Z0K��!sͣ)��a�Yݔ�q0��r�6JD�MO�Ht���F�����n��Tx=��qt"t�`��x�`����8.l<��{l8�Vpd;k�����s맶�\��X���<����n�u��C�l��vCvkZ�e�%�g]:��m���Gn3��J�ݝ#��n�"�.h���+�l��8�ݸɭ�z�:v�Dnl��:��[��;� ��6�0�(��4=Gq�Gvn�u�9�n�z�/���u���85!�v@Nˋ�uv�u�����{l����(v��C��v=���Ô������v샘B\��3�tx�o;qC5�hv�8�e�v�[��-�Ÿݞ��Z��n]�z�;<]��a�gjc�\���竻��"\�i�KԹ�șP�9<9%�v����ܕ�Y�h�=�v����iO�Cl�v�j�z.B!��5�y�k��.����/:�-��'+m��mۙQ�ٕ����z�l0<�/6�>D��fc��Is"�\�nˌ�#�Zƛq:�#��g��e5����n��a��ۇ��ݥ��hvzľ>�����=�y�W=���V��ƺ�ɘ��2㦔#mG�sڊ��[�c�Oo�=���:���I��G/lv�v܌z��lOm��8fltVgS<{Q@�:����s�6���Di�n��I��4q��~�<Gc]�!�y����6t;����m�3[Iq��>�����]��^�8ܱg�z�n����SF���F���/p��6��w#�l�m�g��l�F�v
&O�dC��a�yk���f��m�ҋ��kn��nev�S]��s�����Cc�O܅�NЁ�'�]��r�c����u���E�*n,j�ݧ=j��n�`:oG,��%^a���c`� �3Pr�l��/
���R.װ��lu��M�.lj���a�F8�	D����㩎�]�a`v1��u�غ��\g�w�XG�7
뚵�v%��u
�+��6�X�5�r�e~��~t;]�0��ms�=���n�p�p�	�3�'�Ng�pN��܊ma�-n�)փ�sԷpB�4���آ������nq��s���+vpl���[aq.��@�u/��nQ�x�s����;[q�f����\��:��W����t�:;z� .q:㖼��t3]�%{�;<���UG'�i��jb��4�l��ŵҭ�r�b�m����h��<���@-0���}���w����l�$]�Q�PbUTF�c���L��wwr�-ɍa��*��q/h�4��D�T峣zd�ب��7T� �O3s�����VV�UU�H���s���ôav^ڃv�u���1�q`y�q�&�v��ۧn`�V�p\v���3ͭ\�������Ս��$�5y���nEïw��u۠B��յ��x&�'N�'��c��"ۦ�盱�{N�sn�Y�=��WgL#D/D�[s�<��4ѭƭ˗�u등����G��ۤ�ڃz�-<vN1�í�;�x
�9C�5����]�[�Ʈm�i�5����t�unnn0����WQ��)�8�����qQ'p]�-�<�f`7nS:%z�(�U�i��.]�k�n\��$�����ַN��lvm����mR�82�`���[P]oiǮ�a�3�� �JX�\G9�#�� ��2����n{>�Z��:!�t\�ݰ���8�qpN#sz�=vy�qْ^#&an����d�L'Z��on5+�n�Lg�;O��1��rk����]��r�v�էs�rm��d�'�o[�S�
K�^:���x�8��\���[��sV���9Eb5d�c�����{G������s�>}`*�:�]��p@5W�F��;�w\���\f�p���zE 6Ɓ�u�$C�%m�m���ya0P�ڷmq��nͬúr�j	ձ3�*,��K�H��f7T��9�ݎa"�lF�]DT�0kEu����Q�5�c���\��κ���l<��i�{+onQ����5ͭ�kk��:�mr���NĄ�u�Ě�[�{p�[�x�ۍY۝���S� ���Fso4s�s�a9��Q�tR܋���<@�Gm�ӷ[8���ծzz��r�'�ܯH�ݰ��������r�K���vI�Y�.ca�ۃ]k�n�Ne\c+#[X{pk=\������P��]I-�x:���[���nݵ��c������skW^]�s;u�wnò�hm�Fy�ۍ�mݧ��v�v;]�@�-�w[��HDM���(�����ֵsDK����K�&w�T���6����k@Л������ܡ��[6<��y�� ���37��6#�kl�]����ՎPo-�g
��۸�n8�!�aܳ��b��ck�7\�n���=\�a�%P�$�-:�������q����O���s�\[�1\7�8l�.�e��Y�\��t��2k�[���n"�&����T���5�w��mە\;�|d�qÃ�g���d�a�0l��v^x��+�������j��~��v6�6E��Ͽ��+,�/iH"޳w��5��ۡ�X�''���,��Ğ=�Q�I(��~Y]�P�A#���v[[�M��k�e�B�ds/.�Ȕh�3H� �M ��:XÕ�B��k�x�q�Lf���v0Ax�0�G�y��@ h�4 ��pV�Eu�9��I��`�_�  >� �4�{Cz���aI�qh�Oچ�
��t�[ﾼ4<���g��ӛ�r�$t�Qi5䉰Ey��:뷪n:�J�k>�4n�+=|�-"�!���@�DI����TW;�Ӱ��"���o����D��VcR�Iﾺ�g%�m9�r�i[�=�6,�?,�ر��r9���8>�=��G�g.Ӓ���'�s/.D2� XF�Qi�U�#) )2���3�u�t�y�ͻ[�{���mw-#�?B�%/vi��Hi@-��#J����Vb��p��T��2�`d���ݭ��勐�3,p�Y�d���v�d<�{��^��6586� 1(���u��+��<�s�9*U����hy3����jr��h���A$H�L_z��� �65yd7�L��	�@K4m�8׹�?x�8
(�`�J�k�P����%�Ec@�D�dQKݴeU�u�|�]���5���:%�I�W�Z�7a�EA:�}�����ˡd4hI��:�V/��P�v�b�hc�d��,��n�;�ª�I*Œ���V�j�p�2�Ԏ�W5~�V�	�/Z�};�����s�ז;����.(ߥ}���oY&a�NB>�E�l����٬Pψ�LH)J44t�9�J	a�l~��ٺ=��D�i�^�*��`��$�@��ܠ��4�#���G,�'ф�F6��q�ɣh?1�uZ�~������(|��/��n2���Ͼ�ڼ���.�Vִx���Z���VV��8{�{�Y���7��޳K\�tž�����j^&��/,��2�zH�K?}��U�������԰����ap	��$T��@��c�Z�V!
��	�3���Bu�"�a�!�D�ސѢ!d�����ٙM�{�',[�w1s�ʓ�O8��n�q�u��w=�w0U�z�V��ugNM�j>��{����������5ɿL�&����A�^AXwPdYM�5HO���N�\���V�p��@�"��+���Վ��d2�oXڛ��~�w��œ	�\�E,� W��ä��e�dg�jI�E���	4m �£���d�L���g�i�S�P�A� � ���vS������㒴U��gab A�����0���nK�h6�N6�$��\��R����VN$� �jnz��d�mh�NG��/�'�0Dg����ר�l"k!��I�L��V/���.����o��n߁�ʸ�/��!�|�N���o���r�k�H�HqO�]��m0 #��G���u��}�.�28��Fջ�4�7�^��5� /��{v������9[C'�
�\�`π����P^/7ܪX�r l��p�ꝚLy� Z��*�ZPYo�t�B�e�h�#��%8���EO�����Z^M�=���ݎ���6��8@QiI|� �y�1��}���:�Rf�Q'A7�Ox#�NtE2����3$;6���v������ug�i���L�:ު6:�=F�1��0��9$@\�I��6~�y�5�T���m\lW~wY�}}�HȦ��rB#��U��]��5粮j���/Q�{�}3rm�AG�Υ��3,5B7��rz�!*'0�L��+3=)B��ux��B�\��9ߦ�y��E��"*�,���f�45@���Y z=�E!�U�}��Z�S�XC�[�mW���J�c�J�E�� H �7;��7�L��+��ӏ�0{���J��)��:TP�QEV��YWX(���Cdm-�I�;X���<E��i2� u	a�S�Tm�#H��8���ӛFf�<|,j��_f�)Db����bF�@��1B�|��J�5�Bl�s ��Dڮ?{B���Mdit�{6�d.�U��B�cu��;�iፕ[����R',���Z(v�p�tg��^o��v*9v�����Wov���[��]�uzI�k>!2p��L̅��sj��ϯHce���g/[k�-��/���<�94!��� DN�z%��+��K�B	�>*��:��f��D���8����ә5$���vT��V��=j�Þ������KŞ��6�܀����K���z�]�k�g��"�:^y�?+��X��D��@���v�� �����O���Y]}[G�Đi����_$@q���1��UdK>/#1�.��K�=0�N��=}���C������\x���:�e�e����l�:]�,�������l�ʵ�KX��^���^Cof�ev��|�KA�Wey�K�m��%���a�C!�Os��+�k���i(@�i��01� ]���i$AhtU�YE"j�\��<���wn���cϚ̧Iky�ν<���w��)B���_z
AZ�R���P��e��PV�����U�ѥLQ	������{G�Ǟ�F.&����n���X�Sz����dn�/2����w/6�n�s﯍ix���D��GJ�-P�i�$.�Ag�A�#H�4�
=i�uW�Q�'1�[Zl����/�ػ�h*�`����}����T��9a�/�<��#9b���3��e�^�.k����{`�QKM
$�!�3�j��	�6/D\'6ۛݳ/W�<<և��{������n��Ym �c#��Mt'v���7G#v<��p6�՟:�����C�N4WMzwZV����Ӏz��ƣ�/\mڹy��"C)�3�Ѻ�����n7K�c����v�@�ẚz���wO�Nܻ>��v��)���a:��&Yk��r�F�o)%��۶:��0���K��7�)��לq�\�u������s��3�8���u)��/&.3Z2���wx7y���z�p�4������e��*�Bq"L�~ a��/��8*M"�D;6�Po� �c��A�L?(q��/=��m�4%���[)K������//%���$W�'��Q#�ˬ!@�b��M=���4��;+��$;IE�9W/�VB8YG	 K'g�V�����%� ��׿RE
���l'DSN�n7�	, cB��=ϱP!��@��}�C�,�o���?9]J�����S?a��ů+:S����ޤF��<���l�0����!' ѤI���k�S��Zޯ��AD�9
�A>�*ɼ"�|1�����B�$}�`q!�<|6-��h&W�U�g�FDez:#+�yQ?�rF�NO����A��i|*N�*��X�	!D����;��\(�Ux���P��#( �/���`"�P� zH@#'*��CcE6@�F�U�cz�s[����w�'w%��+�dˍ�ܾ㫥�\��JA�';��ۜ�G�7Cp=N��'K1H r7RJx:]/�"��8����T:�*�-�����̖��D!�}bV�����х\(��mon�4�=�l^�`��0˗�r8ar)�aG "J�ZU��"���fz�`"��t�����.6i3�����Im�����~�G�]ɓ=!q�&�D��V Lֿ+��E, �����+�di�Q�o]}+���$>����2,���弔�X�� �����5דҠp���#qU��5s9=�&���_�pW�y'$WȒ��}�Q+�A��6��ڴ�]���~h��sR����4�(�ɻ%�� �ʟ���9[�:4Sߎ���0�\u,鱗��f�@X'���H�/��w ��~sI�W��w_EH�^�}ۇ�!���H�mO��I+_ax�T���.@��8�a�"�D�Q��L#������[����[A�.�]�SD���K<h��
;�ǈ&�*��(�g]�++��k1E��@p.h7�?\�|,�6�bNĘvM�`�$k'�<�<��u��Þ:�⍸}��^vJ��.��Z�c����%�V�'����8&u$
�r!mC[�Uv$�@����f�gY����/���C�G���ӇOȤ�G�U"}�[�6~�HJH.ɴ	!�A��؆NK�1�{fa���4���٣����M<�G+���+��He��~���T?a�����X�qO�O��K�n[x�n��7"���C�}_R�Us~�F���j� t+���H5 ��=�,:���
w�v�P4�"܂���cx�7�/����(o}��[�)_)P�2�r�t�[b��^t�)h^ �+Aj��9>Nd��#�{�Ӻ��1̷0�92�-0�c9H�����8*s���(��U:��Oor�sw�4��8Q&�&*{�(�6�h,H��襁��>,�@@D �`��-I�#iv�x]s��	p�3�}�5Ÿ
qZ��g���3Y�5��}(�Cڇ�zR?S;֥�Sŀ>�?l�Dik�:F�����Q��O"�B�Jq�Qz�:�}��nۇikhX3�]3z�uv��uxFe�I%��^e�_"vZ'�?G��}G
�$��P!{;UX60�F>Jć��
���+�n�0�``���܂��I���X�<7�.�����N�x2�V�ɍu���~��t3��� y�Ċ C��8���4	�Zq
,���T*  ��$4Ȅ���n�'�\��_Ϛ���|gY�s.�R&��EB���P�KӪ�����!1S�B������ӪQ.��W��OD3�$�r���WG�I��d�m��/�˼r�������W��#����H�\�K�B�$`$� ��=����+�h�,���;L@,�"��f�ȉH�~~Ք�n��aۮٓ��N��,���ý;٥�n:E��m��9͂N��f�T��8.�ƅ��ɠ6�e��Z$q�x%�<_Ob�	^�C�H�pc�WµYGʐY�K���G���C3���4_�2P�>a�%�Q���!�A��ǈ��"vf+�>�+ D˿L�ʘAl��� (��G��l��d;u4�}�!�<ݬl��v���	����!v����#�����c��M mmWr��PB�<�$�,�Wv	�7�-��՗�V1�D���(�4Fb����B�V��?��~�3//&I3/2�y{8��i[}��>�ZOt�&�eq�a���=7#�,�H��!{� �Y�~_C�uʦ�|�6'z= p�ͤ}�禓ZbD9�����8�a A�5��s'}��i��Q�P5�ր�e�}�aY�^:t��U:�40 ��#�����mG�ے�}�?_s2�w�6�s2�)&J������O�zY�7r5�ڽ���閭rήغj$�n��F:�?#qO���ܠn��O>ݛނ�4�}��GT��o��s�w�.��8��~P��DJ�c�8q^J4Q$(h����Q� ����X�M1rD�7���4�E{ˮ��{_k�©�c.�����g��'\��v�-����IoĄ�䣴�7�px���/����6=!��T*����&���-��M�f�p�Ԁ;-��,
CЛ�Cvz�x��{v��C��l��k�v��v��r�ta<�nD��F�]�q�g�ڎ�pQ�"��h���ׯW���mַ=y�n�Ջ���:䵏q�����؋������kÇ>۷Y��=�g�$�<������y�nɻ��@G��ۧ�m��<`7�ԇ�`f\�g�h�n۰�z9��;\��d��z�vI^�ղ����6��!��l��7Y%4���V��_�@DLK�~�}��v[l�>���Gǝ�2TԴ[C��
�j����dpB�ڠ*q������V�@��ӧ�=��ancA��0a҅��9T�(	hCӮ� ��w���&�}���+��#�]!Ap���ຯ�?^���>��>�)���{�kS~F�D
�r�F\+f33�52A������W��?1HON�_w��8�	٥gf����ᷬAx�%���o�{Ay�2�&&��~&e�yn]�L̕��>��j�M.��T�v�G�*�T=��YV�_I`�mv��-U�YD"A�#P�L��x�Z�B��HJ��I涎kB�&˟G�1s.fg� <ޞ�4���gՋm|Ι�-/^�
�b/��U㠅H��_d��Et�?#�����^]ʻV����ڲ����.��z�ڠ�������X=�//]l�x�z�τo�5�mK����
��O�.�Y2Zۘ7-�2�ϕOB�K����U�D^��>?a��ئ!G		#
:�* ���YuY��;�+�Ax�5��$ο^�H�h��8�Em�����m(Qŀi�@�"J1;��ux#�N�=���tZf���g�S)j�l;	��鋞wc
�՗���u�ƙ噴�r�9]�_P��'�LL��S�]���}q��~՜��Z������s�~�j�u�����>C�dT	7]��'��i]��p�k3`�j` �?Ϊt�$�y�iׯ�ǎ�~������h�H�X��Q����z�Sl��i
����q*����j���@�t�q6���^���'�4�ϼ��x��p�fe�M��\m���{��ϮNC�d���*��C'^�#ꃆ�I�;����iQ$-A�Nuf���=N���i����rG�Wӄ��ʷ�̻�4�R�鋩Yvk٫�oj��)�K�dZ�Wf����/O�1�H�ta� As�X�[��a���G���Yl1$bV~y���rsY?|��%��/KH�^a�g�Ë��� Y�&�$�Z��'@���v�&��\���	9�(Dp�0l�^�=���,Y��$	��˭U�84T?��_xv��v@p��X�5�r��H���%�cv�<�>�m��r�2�Ï�m:��h�e�߸��E����{���s_���88~D&�'n��]��9�"H1"קX��(u�$E(��x��  3����d��92fe̗�F�#n%�m��E�|g�p� �^H��,���H�|�'f�}����~!�wPz�\6RV���+e��l}����)ͦ�Rk��Q�kJ����hk�,�Y��%մ�]b���7ٕ��#��{�����CqZ�h�ua�Y���v��]R�[��%�]$�#�ݠ��t���r��(�s���G�pP��s����E/\���{�6�կ�or^�G���@��'ӫ(n.�;)I�6œQh�cH�� ����F�B߅�[b���˼���}�:�jCÍv���"�_W2aplBR���^�c=˫�Ze,$�:��vW������$.;�µ���,H�JH�6�1���Zi1�o�k46o/�1��c���`�s�+Oa�Aк�׊�Ke*����s'�kwp5S�9+r3���M�Us�;�M��Se"�4OJEu�l�=���������L����!f(�
"�w)��⩒�9����Z�ټح�����@��aͨ�5w�`��V�g��e����ks
�P�Ǿ�Qs�%��Ҿ% >-�vo���e��x�t߱i��48�U�\�0t�f+bQ;SkD��y��8t�=fy��HZ虴��S���T8b�[��Qs�7�'&�!��*��M�'����V���u���n����̼���QKᨛ�nL��{���,����x��C2�t�����.�o�Ѝ'�#f&G@�N�K�}�R��f�py=a��7��ޑ*���Jz2�},�`��K3�7���B�i��1��Z-�5Q��s�4P�����h�DJ�(ԅ
P�y6�((i ��Bџ���Tm��Q(�
P��ƋJ�:�(Z6�-�%?~�����dr�$�sE
Q�(�DJ3.�����a��~�&ge��B�rCh�䶍�����kmTJ��Q(Z-�!�Q(�
P�m�%
Q��~Ѣ�(���J����@X��~r�M��(D�lA�H�3��r�G����P�F�7p4��J���\K���m(Z����~s@}����漖�)B%
P�OJ-+�J7!F�(Z5��<̼��^`���AǉB�"P�~h�h��(�iQ(Z6�����s3�4P�GZ�Zw�1J.J1(\�E�
P�h����~�{�x�h�{sTm(Z�	�!B�-��! ���"�ե
Q�����M��X[G�(Z���F󙁃��M(P�a[�P�G7�ކ��P�y�	B�)��iB��z�B�m�i��(R�P=������+I2�a��i�c �ͧ��;ﱟ��KǶ퇖,�"su���κuG\�����e�(R�A$��҅(ԅ
P�~h�B�"V!���k��j�Q(��-�q��h�B�A��\!B�-Kj�9�q(}�_��B�(q��&%
P��4�Umh�B�d��y
�ߵ�MQ��w���}��gC捉B���4[G�
Q��A�-����8��(��i�=��-4D��vJ�)B�戕�"P�F�$h~u�w�nf^Yy�c��tm(R��U֣Fڱ-���%?%D�h�DJ��_�E
Q�(�DG���o�s�k�J���B�<�m[U��\+�B��[���j��h����5Q$h�D@{�-+Z�5�P�F�ڴ�J=�?h�B��#GZ���J5!B�-��#iB��A(P-#G߿w���]��J$�
P�5�����C^;X����J�j'�h���z�����f\$�-o1�)B�_4ZU��J�h�f�zk�TJ5!B�4~���ꍵ֪%�w��ġh�DJ�����h�Dq4[V�n�~��(R���(R��Ƃ5��~�'���*�Ѧ��(H'�-J�Ͻ٠�ƣU�렼�
P�cD@�D���4F�m�҅����~�4$J��D�k�y�1(\B�-*�,"Q$(R��־�.��dnf��2^Y�6�u��"P�w��h�(R��?o;������|V?4��"P���]�;�@m"D�|�iz�K�%�([��4\�(�"P�
A��w�&��P�@�����Z#F�B�>�-1	B�-Kj�ġ������rQ�(R�hٻ��h�DJ�?k�y���ބ/�s�{���o��L��ށ��]2N?x{i���/6h�󠧮����c��������0oM@�E���)y���F�+��
�M e�����j��
P�
P�cDB%D��-r[F���J<l����fF�d�m�̽)Gd�4D��
;%��Th�	�҅J�B�J���ݚ�iB�vB�(Z6��
D�����#F�#hB�7��o�g��.~>����2���@P����	�&���}�{�4�P�*�J��j���m1����x�OZ
Ƃ�����Ua�j�^Ha��ɒ�/������.��juvݷ3u�Lf�'n�wD݃\�Z�e��#r���r�X�2�r��W��G�(R��m�AH�(;�im�4cDh���z~���P�G�"sPjڨ�)B���-�iB%��r)�&���M��%F �(R��6��
A�
�kI�%-�%��~�)�.��ｙ�����4cDJ>��5۔F�ՠ��-*�d�Q(R�-��>��kޕV�I
�N�Th�B�(y*?�۠Ǝ�D�J5����j�	2�f�:�(P���iB�j�G�"P�]��JM�(P�4O~��5F��Q(Z�������k���~�����(R� zB�(Z4�4���<��w��(P����IB�jB��j�F�"P�
o��G���^��P����D�h�G��J�B�)B�ƈ�)G�}�ހԂ�rJ<ե�T���Y:t�i�A���)AJ5!B�-oG��dm��r����ɪ6�)B�-h���(䁴��-h�B�g���E
~@�iH�-Tk�
�f�Z1(P6�(��8�*�7�}�j��G���X�F��:�9�ٯg�?f��G�(R���(R�]��h$J���ܣ�-+�F�U�([B�-�j����b(Z3{���m{ܺ�J�|�D�[E�
Q�.�Ѷ��-m���?�ݿ���9���f��D�h�DJ2B�%�(Z3�4i�_�u�����(R�(R�����f��Tj%���h�#V�iB�w��B���h��д-Ti�����q*%@�O5��P�
P�G�"QrJ����s�f�����%mhƈ��D�v�h>�ro��ow�h�B�y���q�H�-4D�B5^��2�"P�OJ-*j�
bB%F���9Q�~��/"ff^d�u�P�F�ܫj�E�ii�u��-"P��Q(Z-�4ƿD��]���4J���ֈ�b(R�(Z1�5��jB�i��p�l�h����j���4�m(X�)-�-���J4e�B�h�Bյ[��7��*Ѝh�Gd(Ԕ_�#mTj4y�%
¢P�Fo���Q����Gd(^�!d�hġJ�"P��Amh�B�-{�F֨�R��6t�����޽���T%c�u�we�x��;՝%�QV�Y[~�M��;i-j�j�BCDE�ؼ�����~��}��'9���YjCn�K�Iڶ��޷�}79�6�ݖ-��J�wg���e�����K;�n��`���m�i��d��b\oK�sr�[]�\�� ���Œܞ�Z�p���/M\v#�:��3��lBog�������ь/v͔�R���&;��'nyiFL�u�|��9���U�,�n'.zL�����1��>�pj���O�xQ�[����x���0ܣ΋�x�������0��XB^9cx32��P�
��PKJ?���P�B�/�<�P�Zj�B������f��P��)B�ƋBҢVnwVP����6��(��ߵZ(R���]M%
Q�(��׿j걣�(R�H�˅E�?rj��֪>�t���o=:_��
�Hך=�$J�!B�#E�F�h�Tj~���/�-+�2Q�DJ��]X�m��F�4D����\�G�����d˻3�2�VfY�6�)B5ƪ4_�Ӕi-�4ZP��j�oЫJ�h��֚����4P��"�E��}9����}!B�.�,8�my��B%���+5�}z�iB���B�(Z6��---�(R��M��%�s�(R���(R�h�DJ�4D�C�^p"s!B�-w}�4x�,h �j�Dh���߽ws߹[h��B�d���t֓�E�[DJ4x�Y��f	32�P�G�"P����J���~oMm��J�TB!�-����MQ��J=%Z�.��戓r���)\����B�ڴ�J���h�J<��҅(D�k%��o����f����14ZQr�
�h����5F҅�`-5)��-ha
��yh#6�-�%�߻�e
P�u�%q�a�R�B�-h�B�"Q�iQ����/�9�v��s#r�l:�(R�HP�~h�h�(D?k{�=�7±(Z<��({�����B���)B6�F�5h�B�jB�%G�s��������J��D�J�2�ZTJ�&zV%Z�?k_�e
lC�[GZ"P��Hk�F5�Tb�iB�9���~�?{����hJ�h���@�J��)B��;��J��Z6�Ah�G��������$�fd��h�J��D��J�h�`c�FHQ�A�Bў���j���Tx �A���[F#Zh�
�߳$(R������u��_�Q���gw�f��"P��N��4�"Q�-|5Q�m(R�L�X�-���5F҅��A�
P�[Ff���Q��h'9��ZM�[mj�����ހ�s0R��h�ZKJ�F�U�j5Q�d�ҵ�w�h6�I
�h���<R�N���o�F��)T�!A|�ڷZ�(��Ӻ��m��'q֜��n�ɭ�z.+�t��%����?%
P�B��K��4D�J�C������Kj؂�ƪ����͔)[�h�V�j��\��%GZ#V҄J*!�
�Ϸ���J��'�Ui����my�\C҄J�Z#Q1-�(R�ۿ޻�B����>}�o��>x�҅(D�J��D�CSvW�(m*$i����n�5<��X�#]j�P�[hZP��`ZF� ����m��F����o���pr8̍�KÅ
P�|���;�k
.B�(Z-�%
P�B��"m�k�?:�j5Q(�\ߵۿ�������s������nu�T����Dw�$��ᔖ�ɡ����J�ĀX��-������#��iv�'V_|�B���J�s�0@ĉBѶ��m(����6P��9r��D�j��%^�Un!��J�r%F���MQ��d�r�ġJ�4D�J.B��{#F�#��%k߿a�4�+b��(Z����2��r�!B�-C͵�@ġ��CIQ���r~�3/1������8�-B�䪶�Gc+Im�-"P�)JP�cDm��g�����Ԛ(S���4��j	B�.���jB�HV!3�;�(Z/߻�Q��h�(Z1�!�־�������m+�ݔ-�ƶ�N5���C���6P��<��o�-(R�IF}(��h��%b	p����h���]Q���Um�ەh-F4����U9���� �	m������w,��W���p@���ˤ+ي:�,x���졕*c�����P�5�� K��Dy�{��Isz3�^��Z�⒣fW~�cxe�x�L�3F�v���V��a�2$�]�e�B�b���7�ux�d�A"r`����ہ���P�E�A�f�?A؁z�u.��ve���T�-���2R.`�Ed�"ݟMn��E��d�l��N}���'E���n����v�&c^|�Z��э�o�N;!�\�I��ҺgR#[E���^#+f^t,ovoJ��kݔȦ�0��}�5�!�\�Wb=g%��W&,�q���α�7�m�����ҽ[h����h�E4�!�"�s{��|#DjI}1|���AZ;�A|	]uʕ���s���x�N�~�F�ɇ!�A��^IZ�*�q�c.=�W����!	#>?H��ϲ}�e͢R�����9�/��]A�.^v7{�V\J�c9�rvu�4d�k�l����}4��t��jm-��5�J��"7���n��,��*5�'Z�8}b��(���9��nj�>l�6���Yu.]���*���>3*`��zG��ҁй<���*H����`�{��>PC�@7=�8�7�h�~�g�箊��Lfm\h�ϸ�+"0�"JY�v��Di@�.A�
)_J"�k�H�ڣ������$@Qzk��8�WI�S,ϮcL���z�X���i��<�����@������1��ۻ�|��߽&�ְ�{9L������W��c��n�1vx�:�@�v�nH�g���7E?������~��0Q�&X 6��"D�_AvJA(Z�Ȣ7���p�Ӎ����Xq"b@t���H�n� '����-�a�(�MG�t$H�����4�>���n�]a�c=Ƙ�d#*��@B���*pq0��U�GWh�Fj�F���Hł4�,�I��qn׸�q�����h�O�i�Ԅ��F0�~�6	#H���Ճ=�?����Qy�W߰Se�ӱ�>D-Hմ��;U��D^+"s�a�R�R@4������	�;����4d+^�rk�r)�P�}�}����)�@�._*�8�f�Z���S���[���Ptkc��җܥ\��]W9 ��{2,�갻���xݣO61��ǰ�ʲ���\�=�o������2M콴0��
�w*
��@�S�<o
 ��9�i���I7� bX��9��M�kofm�QX����]��|W�ꡄI>\E�5;�
W&fM����t�W^^"5|,��f���&׬��!,=�qѭ�*{jz���S=�V�u�v��K��� �n˸�y�Y2�-fL�a�9y2��E��}�������+�V���[�L����s�5eg֬�Ȑ�_Q�X�A��� �>�H@ ��i�s�^	/̛64��|�Ͼ��жZ~[���:�F
���ZOʰ��I��d�!��;��
�� #�"L�����A�4�/[�t�0eͤ��]�2܉�w�p�����0(����X8����g�ɮ}3�1�Z/�m�粒ڹ�.	훊Ń�)$	ĉ�4�N"���20�#�>k�2�䃅�TqX��,*��kDh�(t�D���K�3@����:
F+�cW�~~��C-c@���ȇ�`W�p��$r�L�d��#{�%FK�,o1�o91�+���	'��ݽB؜��M���My>����q�f"䌓�.)y	�o�Ͳ���ո�~ϛدM�G��L��,��r�v���6��]��Gx_w*���t����X��S�w��[>�]���3.����]��26��K��2S���|~���m�RW���f�Q��3���ڸ��v1�U�㧛�t��Sxu���C�z��q��O�f�l���K�Yw-4v̼cg�\��^���%��Jg&�n��n�v8�N��d�u��}T]��A��wn���퇳�*7Pܚw/Z���!�5y�t���bN���˻Lgv��{OF�5��<n^�s���f������FNuu�n�W���n���J`"��壷S�ٳ�*:N,�zۤ�m�:6
��C�sg��Ys]��3/.엊d̳���v���M����8�d[bvT�{>���ՠ�I��|����0W�J⨟�x� �n��l�:)E"��?E/va.]�e�Xq��y~�:P@�}���t�rc���G�yI&�<;�7�QڱF�]�Eҥ����v�����0�OѪR�]A��h� 6M^:�t�n�!���\ːr^["���aʴ	{��p��A4�H(�Z�~���t�Z~ٲd�׮�M�@ Yj��@g�)��Ȩ k��]�(��Q����✍$P2񙍚x�j����n�ͽj����!��-�B���Y^͕�8��Be`��Xӫ�G��8cg��3�R��a����'��b���e���E����Sr��_���}� �Vys1:B�}@Lz�C�\H�A�s�+�"�e"E3�܅�?aR�v��Ćv�{_��E��G��a�\�mUW0�^;���d��� ����Ǣ�ZG��%ɗ�w�3+Od[k�X�5���Z�v��,t��b�h* ii~�t7�ī��(g��ꑝ5i���u:�jyT��.;�!7K�>�$\��32�&�u��RH[I�y�>`_9=�F�'����6�(t�d�����G+���>���Z]��U����o+F����Қ�=���U��}�>�2�J*�|_��A��]��b(,A|f�ݔ���AԉR�7��^#/��FV#,8Q�����%��ř�x�q��6���G13���΀���E ��] �l�*�spi�<̽�-^�j�H�o+��ù8�V�(���Nz�GS{��|/��NC���Q)���E7U@m8Nǵw2��w�� �C!ڳ^<G7�(M�4Ô�����d�����ig��;��{4����w�U4����t/��^�,�`���	Ƞ+��#$b�:���+▣��;��(1�Ɠ�`�表�8�%Az��Y�K@i���v��;3��q�}�'�͒'�qW�B�#�$�t�&bt�Q,��错��������[bB�A@��H�w��̇� ����8�=F�ӧ�N�>A�Tn/	yqf-�/0��}�n�v�m�m-f��\&}�����b�X$�fr�x��K��(Ș%c�_f8��Kұ���[�+��hB2W��ܹ�n1��M��.��^7��伻�Q����$�S�<�o���vs���V����>#�׵�Yl���~t�G���/����c�����M�n���`d���_�N�}�����I�}#��//*fb�x�d�Ťq���F�G*��Ֆ�E+\?bC����օ
�p,�C�kZyHǊ{u��Y���vQ��e��i�XP�n���Z���{�q��L_< ��M1hq�F�=�S}�%�k��!]�����!�8�@���5DrD�u"CY��Y��U��i�y$nѴ��]�H�d��Q��#�Z�����^��Y�>��C�8�W�%_j�S �(
�@���`�+��4�ڻB��uի�U�j%��.��=�"q!Zz�܄j���R�MR��]�|"�aH@�n7��di��G��Z@��@PtH%w�C����*wT.Ϙf*���:uχ��]F�0����B����?0���mC'}O�;��Ț%�Ŵv�8�okW�^@i�;��X��U�u����3�ɘ��9�z��e��}�.��{�^����Y�b�!@�6s�ŒI}ө�/�[Y�@Z�;H��O*��U��x-H�+=��l��ABr�׼]���P$c�P�@���(l�39�W�p��˳F��uD��_Ka�u�W�DQ�+�o��w����rm���fJ�ٹ�X>�}���g{r��^w���܍�HKu��33,:�q]FI��2���ݓ����%�J�o�MtP��>���=:��>k'I�W�]��t�u|px�&����"'5�s�d�&��wŭ��GMF@wG��N�rt��@�����R�n�7�j�����-�*n��qL�]v�Nn�^�{kGzŉvzg���Ic{V��i�D�;Ѣϝ��}�k�P�oI��mD@Ѳ�5���U�u�m�]�a�� $�k��L}���r�E�Ii��9���f\$B�����F��B�X<�b���=���brg|��9�W�k�	���7�QT��>u���d�X�l��e`A� ��B�٫o܏�Դf��	._�Y�t�̥�f,���V��Ю�pl�b:f+\T��hj���U�{�����E\IϯN2E1_k�&���cD�D���7�=Nj��w7 �2�%�`�L��0
�@��G�����k��ؾ��s$%���Bd���>��Di2NE�Dﳍ�[���}U�Y�C�v!y<_��_#�2/#�s��~.&}�<e!X���i`�k�:��f�{�X��@�}f�E�sj]ż˼̽���WO[]��+�	�:P?y�M�@�gn�ZO/�0O�:��AO�ǂչU��n��*�[}ʸ��x�$����F�RD�P!)� 3�6� �A.��9@+��z���Lkǫ6�eA$�1Fʟ$:��EEe�p�A~]�\��f��� ����b���e�Ay�eK�	ո�/���y�PH�����$桄Y:���:D�h�3,��gA~=[2�ΞU��X�jO-��2Gz:["��5��z(aX�-B�E>�������r��<6g+�y[�V��Y����X��D�m�$����/nk�ɧ��ڽ�}���e�Jh�%z��q��Z��'��-(�/�9��u�g�3)�U��A��٫mm�2����^	b̺x����F`��]�+�2��31[�,�����O�L����;�p�WE1�_��7�P7}����[	�{,R�jI�Rx������!�૲]5w��NN�/�h�N:��b���}����'oחX��B��A�ce7�j�=�صW���(v5���6;Y��s�|�i֌[��	{{}F�K����T��Lj�l���|kwss����V�*ųlK,\��.:��<����M�Q����/`^QdR�؟�W��C�=�Ȥ6��'��xlc�0��"Vv��#Ǭ�y�PS�FhWJ�}�q-1��(���p�Gz;��'��oi����N�Q�ny����7	�w� �t�w��n��v�ܾ�.Nu���J�"�%"�0�k��W� `*	C3��s
 l?T9W��hq�i��(MW#�U(�k��_g��z��^�;�\�g=W�[�h`r�2ܹ-��M��kj#�#.*�vX�L!���z�qӧ45�f�&E��y�ȔU0!O<��Q�H�vNc�nG���i<&�N��/a���@�Oc`�p�5h�U#���,ʍD�^��ᩭ3��{���9WD�kl�U�=X��@.�k��*�STٍQZ�X�1�m�&Y�Pİ�UP*�U�0�Kh̽]m�Uåy�\�6�;sG�\�M�܎��)�n]Uu<n�e�Gq�^ҭ�f��vǬ���ے6	��s�nۮn�;�h��lO��u7V�:�;gqd��s�݈��/qEn���`���ú1�m
�ȯJ��;n��i���i�M�`�z�6��ݦw^9a�7N�Di\\Pv�e��e��Q�Zַ8���>"v�s��]s��U�[�k��n7iY\M�S];5r�wl��\tN�[�#�Wf���\�[s��&ݶ���r��6���� �v9�[�{��8f �tm݈ۯ�����S"۫)��\n�� �6�R�'K�6�.y�ѹl�q�7oȤl�ݙ��c�z�]����h(�;b<�烝(=�s���+�ڶM�6K
긴W�l\2�f���nL�r��L�L$n��j;/n\��xz7�0������I�.:}���*D�g�]��l���G���ىxѺ��#�e�l5���{ho9�P�;�\;��ۄvyj^��\�4�l��}�}�9	u��7;�۝y&j�9q��mG3�䗐̀=u��v�m8n݄�6&nO.�lE�p��c��v4*�s�y�mC�Y-�p���x��;[Jz��ݵ��U=���l�&�9m�[j;H'�^M�/�fs�ts��+pm<q���꼷[sn-�.n��M�Z����d�7ox��ڝ�ոMҝ��>[sm�4�ΰ�l�����W6�����.��9����s��k�<�ɽW{m]Xn#�j�M�zy���]��cQ�ln����]�3N^��n��LL#w1Q�_;��}W=���	�$���v�QӮ.)mj��c��J��a�{C��=�q�z��`�9�Ņ�nH�8ʎLu��K��Z�q�-��v���[��O;���5qV�:�]'Q��[�ۃ�\g���]AWdf�c`C���L]�gV�n:�J=nJM����-��)��-�YΑԔk����ݫnH�Y���㓄���V�t���q��n:|nɞg.��ݳu������� l�ڹLP�mt.�=vLy^km�]�ݍ7Qv;g���⨮�q�&��u�9ԯ�M������J���n<r��Z�q#;b����[t�Y��Cv�.a�v�e�Fvq��e��9�:�s�d�Ƨ�
�'n�@;��Ĭ�����@��x�j�v7��̶۱��]����݆8,mځ퍛aG�L1.\r��&a2˹��=��m�m|�:�@)~ܖ��#u�$J@�Iv���oq�ı�{w�G7-_gn�v <���˩�,��	t��GUޫ_Bv��#�F�*^�қ�}�^Kr��0���n��JX0H���r��UY�:��H${��b�Nv���g�l�EG���/��H�bX[�B�)���'��os��'�������wpms2Fd�%�[�;�����oy
�!g�L�#��| �`��ī�� �$\M~�
���
�����nWW�oc�;}"�"F�������d�H�H1� DbC5�EiV��M�m0��B�:Q�L��L�I�vN�v{�$0$טF�82֤>,$
ｃO.�V�����V~%�F���������HPH�)�[��`�_g(��g��llx���PN��7[� �-�_StFB�~$��:�c���*�Hf�������8jmn9-�Ƣ3����k32�f+wl�-�e�fF�G�֙3�m��u��c����ƛ�:'�2R�\܂�F�n7�X���#�����٘�/��LAV�&�X�$��yy�F�d��,����/�cY�/V��-���Kϵ�~����_���Q�8o�6��fZZ���ǫ�V��ȻT)��T]�]��YY[@�\4���9e�7�
��I�ng�T�ќf�qhڽ�nS��q��o�ά�y����# �����*�t)@<���!'޷��� E��$u��Cϸuq���L?%����=���UR�KҠ~~��~N���I}@F�� �>|�xU8e#���Z��5u���j��ǭj}t��|� q�,��ĔH jA����v����@�����-�*}8�Ybݼ�q���y�P/�(c�>ֶ��)v�Z� ��ő1�6n���O�� "�#T�"��쭤>���*�Θ���'��R"or�^�0�w3m��n���r2A����n�=���q��X��A �l�*��7�
�Xw��1 �1,�+[6M�B�/���Us	3҉�)��w��/���C�yc����27r�0�Ѐ��.@�m�ێ;f�7m7�9����8'��+LѶ�k���.I�lra"�2��ۿe�O,�����v�vH"j/��d�p�5� ����v(2~z�̡y"	^�Hnپ�=���^����(�]�v�L̠�H�2~ -��}+���S�n�C31��E{�h�J{����-�i�UVl�_y I�I���Ѩ3�"I�^bI��ԎA�x��P>���ylU��I�CƏ��?�*�-)��p7!A�T���}�K�ʬ�r�|BEU2h
�N�|i�*��P���K�:������t)
�`��<v��>��ʏy[�x�X�>��*A[1=Y�����������E	���}
�)
0�0��3Ҙ�ä��XE�'�#���G�n8!Hܑݔ�`;������5�������gx������x���t%!`�ң��'�;:i�2�����$�	���h�����0Ң5�u񫛿K���]^L���DQ��,��x�߳Mm����r Ó�U�(�J��Q��Rdq���Vw����?�� �I e�+�v����������ۻ�׹D���+v��`F���u�K�۞5��t1���^���f�ⴕ+��I����Ix�������"=l�H_nJ�������(� af���^���x��`Y53hQ��9��};������|��7��^�H����(Ma�I���(�j'�I�j68C?#�w*7^ߐ���K��h�K�bI!]x��N�i��Q�:
b�A��z�i�����j@t}��S��۵�
�E�(BA}�5r��d4'Ȩ�^�`�(���R�x�I�I
��5�K (鍮W�c���E!�g���Y4����wn�¶��c�ou}(}D\� r��u/����Ve���:�N#���O}^�L�͟c]�P�@&�����W�/��{f�"���]w"�>�~u�Q0��/~(
(!6�̫�9�_ck5֨h�N\�^�:�^�����s"���V�:KT�˧u	�*G�y�����ă����XE�QN�wn�x��[���y3.�.��X����J,�ն��N?w�hڌ3�Fr��F�oA�3ج�1#��-}��ޅЈ��k�c�O�M����AY�B��DR_����f��]��e��K�%�m���'G�u�{v�܈���!u5�y���ެ�mE8[�2I3�v^��ۻTTo�w�{W޿�|��P�w���F�ǒ���VkފT=Fz��n�Y�FZ@a���{�V�1�5f��}�{�!��
Q�������_���'PBf�m��]��{7��ːZ��LH� ��AvI�
?n���~�ؾ�o�T^"�(�dI�f��G�m�o��b��|4{Z���w�c��7r�奭�>��Хl]۳l|�u�I"�c�*���B�e
7s�V��w�Z� ly��p�Эe�P���4����Z�w�n�u3~�.���&`��&33�E㻋}�c�x��wݫ$#����rIY��x���~�Y�^�q�z��%�������/�G����[�r1B��u�O�bć0�(�HJ����m�NH-8��q�N 'n{�Y�\�:A!m</˻׃z��4(y�?"II������y H����q]�:�+�k�d\�@�N$ ��a�h�w�F��s��@�̧Ǎon���O��շ�Iġr�ڥw��x\j�I���*���qH�L��{z�x���3&a!s,����6,�κ���[�[�����v�����]���y�j�K��l�K>waĆ��3�\b}�n��ϣ���^Iݲ���wĈͭ{���j�pˍr������$<h�pg��z��u���:���mi:/]�W�̱pn�R�a���sϠ��e=��`y�X�q�]{N�ȝ�s���P�1�N�q��I��Quvxc���P��n�[;qa|���n�m�U�S�X9��f�k��Yԭ�G���$YW/,���Yn�wԀ�ȼ�m���ڏX�ϽyO9w���V�Tc��n�����u�}�{���5�ܧZd�H�Y:ݭ���ٳ�$C�2���ka���#���Q�݂@8Q�e˔U�	�^�t�X���a`���WڛG�`#����d,b5�7ｷ[}�ה�e�4����*���p?�tQ�η��<'���X�ք�7M%Q�/�6v*8po;6}V��}��G�U�j��υ0N׷ޡ�y���Ve�s�˻;�v�ZT��s���}�a��t������Ӊf���ٚ�o2f`܈�%(F����x��� D���P��H��V[��$��`��ĝ�Df.�t�����i�l�� �BbVm��#2��b\@G��k�I$���rGB���"��ڨ�5/V��!N@��v���aS����Qin�ɃX�s����*[I|Q��+�8вwnӤ�������7:0�ۜ��\[�g�#�盗��=b9�����Zu���۞dmm�:��<lO2�ql���0��+�e#H�2^����Nl5���h��ϼ� >�uW~F�C�A[�R���9��g)+�����Wi�Ah���t�AD"�P0��$1�&��Ã3�ÜZ^�,�콸;O��>�No@qo��h��sMJ�� l���&ϩxڨ��5om&F���Ӯ����,�Uer�MmV�#��ʱ��ٹ2���F�y�������5r��#���(�`�������$��M�?[4��	�!�	BE.�Ě��.˷�/0�q�ݖ��,im���޷��6�z"X�ȉ�Z̢0�H �of���>�v����f����M��#*�=�s��6���H�L�������I//-�p��qYŚ�:�(�qw��û��D|=/����>��T١�����6�X�Xf� ����0*�qR� �H	Z�[����T��^��NBi���[����d�#r8��H�ы�.���'�� l(aY�4=x�}���a��w�U�hn�I32��id���f���n�e=���;S�*p�(Fyv���ֹ�����7=0\��ք]��Vczުp\�t�M;��N�~�� ��po��{��3��=`���E��C���^�?wى�F����� ��aձ�k3Q�����_z+�/��ǩ��IV��XW30����[���j��D~�:�3y$�Ԉ$��{������f� 7k(����K���7�e�'�f,,�k���M��_��U���C3ˎ;�H4P�L�HX�n�@R�8�u���ĉI[��z)�G�IJ����'�S^���{]r��	��7��7�ٵ4z�51��ME ��VuٛOS��3���@:�t	����W��g��/F�Z���J�ݍ��c�gY3��㧈���	&Ѝ����˭9���\��ޱZ\e'����2�]��-e㆞H�ҳ��f^镢 ۮz�!Q���4+f��:O����o�&�%�G$
r�]l���EW���7l�ʯZ�l��H���AƯ�v?^[q�Kp�� ���q�H!jh��Y_���X�3R�������]4K���GDDJ�a��׆
:Q$e/�i
?>�_5�몀#G�&��X"�G��'<�kj�fb9Ɍ8ڌ��6yݦ�v[sĂ�d}����ccy3�E���lt�P:Ye���I=+ܮ�Դ!��HZ��~�n�Hm��2�ْ.�܏��1V^�o�I�h�
�m��9�ci|b���ϔ�L�^U��e��$ᡧ��)� 4(�6ppV�Ak�y������4>@|��}��m����A�ڸ(��P$4�ĄD����7W�R$/yhG)�E7� �7���:�����c2�3-7N��T�!(�^��b��7�#)�}>ρ�&�'
#ñ>�0i~��a}��_;��/5
)n��G!���x��F�왩�������$`�G����A|�#}li�����2sA���I#�I����X�6�� �M`R k��"�����������=��ևCN�Y�!ƙxUY�ٖC�$�"[�g{���ןr�!x��(-x�{�4���<!���f����c��;,��ϔ�g��^�fc1�2�.��KV(��P��~�6/W��I2M��K����s�ט�{%�������;{=�ul��"�x�5=ʴh��B�V��7���Q��˴s���y&��C��]�x���ht�����=�]>�7t�ۉw\ؼ�fd�9w��7��3����2�#�*�&�'
��ě�p�2��ή�%x��yմݏ��WZ�t��=�1rk�b|�*�������pJ�b@9$�
����2ِ�Yy��U9Od~�o���2��I������ 3�U�x�M1�}��x{4�:�QR�y<#@�D�һܧ��	^�;��K1��9�.^Y�m#���*(��v!`�t�@� ��L�Sn��ܪ�U������O���P����cY!�Q�S[?�P �?Wg^;�TB#=��	z��.5��#y�[x�y1����XK�C*)W/�X$j�QG�}�팟�^��Fb��5t��4��F]\�9�˸BC�[�X$
o�tR�l�u���߭�/	��Yr�oh���:ڈ��}�9��.�K�B9'ܺ�7^��P�{���2D���F�o5���H�6�)��;]A��?�
��cp0�[�״�2AE�/�ͺCR�w��L����+�>kl��C#aC'�qN�V@��km�ք��lȳu[�lZ �` "�E�I�I���wV�.����Y^9iw��ڳ��-W�s�z&��^�����G'ZЕ�˵�m�\�olg#�۝Lq�ݑ�9�f��F{e7����lu;6��ѣsȋ�=��y��xx�AФ�9<1Ɋ.x]�c��:B;p�l������p]<�X�x�p��q�\\��?�Z.�%I5�q�Iv�ƺ�3���;�B&8��ȷ���G1�m��rm�q�.�gS�<��F1�ٚc>�;�W7t�޳d��I,��9� ̼S��e����43fC7?1B衞LDR'��h�Us�`�ؙ�"t�H�L���V깷�۾`�/u�ƕ_J��ۜN�#�;#～M=�͐��e#.��^^�!�'$(�����P���rϟz�ai糼�m�w*�<yH��$���"�h��	h][�����$�&�Wm�u���!#;m	a3��#�\�X��@�4�����6oҢ��48�k�}/ҊrA-�_e�\o!ӄ"�_;f�|�V�*YH�!}j��( Y��3�~�\������ɣs�[qD��{�4�UH�x!������Z&�Y��~�b��!?H�'|��h�Ң��<md�����W`�.��l^���<,~���f]�ܼ��u�vE���f��	�7g�����Nj����߬�b��K&su�8H?4���Bx�L"�zMbn�}��fI��*�˚t���|������_�[�wKd�� b:][ۻˮ�n,^	�(�U��7\�w<i�^Ʀ\c\7Y�g-�K�����d�k�֓�3-5 ��>KP���MmSq�]^�,i6��$��p.�Yv�\1� ��J!RM;+�X �I\)��ީ1�\��x]}�x$%���6�鍧�Z
�E#�|˥PS�0�C��������poi����^cx�����P��Y_b���轢�N�߽Y[�-�+��5�J�JTD���m���AG�@�W�肺�>l��a���Ǯ��T,�$�z���D�9z��#J'ըwj�ݍ	�[�ew,����q�-���~_�~{��lnE�����X���3�j�2�N���j�]���e��{L2=��~�U
��:�(nXl!��!�u�����󈟨��%s�{W�Y]��fU�c3⯠J p��]�w-u:](;��[LRi")�V�}﷕�6<lZ��9p/�8ݢ���@��*�+�#9�k� ���m���%ٌ͞�G��p��y��4����!ٗ�5�}�4�LP�i� +s�bK@��ZU8�l�D������=f��81C����_o���y�}f�
���Չˊ:I��<r�>��%�2Kr�._:�^4�'��"��lg���:�GD��7d�c���)M@�
1��Ģ��;򻡇9��� '\q�|���@�#D$�k��XM*�Wƚ�\bu�y��o�Nd�b�A��(D�M�#nGv��*�0�
���l�� ��0���&x��}�&,h��k�V��Z_�F�k�v�dA����-����h\AA����H "��Z�f���E�Iw330�<fKj��4�ke�}��v(Ϯ�P����?j���my#i�����Zlw+8�WK�#R,�vS�gl}�1�ooqʜ��W�-��<�+
�t���Jf��iϝ(J[���`��`�5�_^fM�F�3�c�@��m�RL�x�*[X�w�|V�*�-��|\A +^�!���O��]�����A8i����@[mkR�.y�n��#����i`���b˭���L9{�r]1ӵ�1m<x��Y�T���n��[�%\^gO��A_��u-�7RL�]��{F�jP=��E�v9�G�^���T�[�髢2V��dV+t�]S,v�׻o����T�����>��y�`���0e��܁w�ά����v��^ݴ�⭻�?KRll���{���+,�A��Sn�P\(c�M��dJF���TA�ʻ}ì��wNgz�y��;�ĩC%��u��1<��Z3����HJ�Il��+�2�}ף))�H�W�}R�'<�m������^̼o$���H��Œ4��*�/;	�s��R�b��푉6���+��̺�Ȳ��įK���
�K� �G��v�ޱwec9�,k��r���D�|�=ۧ�:<�Ԃ��<����5�=J�=�j�����5c݃��Ә{�|I���h�_J�ʻu�[+�n�kV4;i�]���;��u����*w�k�`4�t��s��C�
ZC7!w2��4v��̛���Km��؉R
�Y�S%�1�a��o������-��J�k
+C7r�|;�rS�ea��|����z��ek5����ig���lY��:�<Zu�/������PL���$�{&�/K��� �O)�Bշo���Բ���_m�6AĢ�u1�s�x�y��!
2�ήo��I��Q���t� �"����{����&y�[^Mצni�*+�>P��KT��4�+��w?�{������%~�R!��	���X�0�l�?Q&]�ȠH8GU1F�o�D~&{��=^U��s�hV���Ґ.v�ϣn���\Xлc���9�t�}�+l%�fL��j�R˗���u�8��D�[������<wr����b��}*�EI��0�#�]w"�]��\ݿ)��HE!�~d��W�vt�DV8��z�vσ1ɘ��^2��5(�پ�N$G�{�?�A-"4�2��`�i3ێ��	��ȊB�B{�Ƭޠ�"0�4�?Ww9`�!y��Mo�qV%Iݻ����-#""2S����6�#�2����ӷ;���o��v�2�j��8/8wnh��w���⽑��19��~��1L�AH��Za������Z!�I b�x�.�? �\ :���cJ5�s~w��q���gӽ���{�V��=:��S�s���H�C�E��� դ)H5r��i��Z�A:x��̦����;�M��آ/b����3Xa1��j^�^�fn]���Ǟ��t=�(�v���|�]�:�����Do��r\B�,L�s2l��Q�\�����ޔx���)W1h0�NcC&�T㾡U1^=g��dZ~�h�~���b�#L �O<�7nf�"(D����|hzj�K����:�̳1�m�ļō�#\��ۃu��^�`�1����a�p'�"(W�Ĺyy����E����ob��e5;�-w;�������Os7%=������}|E٠G�'rH�Mʰ��K�Ѽ�!�������_}��"A:�e���C&�s�Y��ᙙd��WiB�]2�@�^roy}>,�� �{�~^�?-C�w�a�(�4� W ����oP����v�����}��)z]�}\��ϴ��Tܻ�S+�oŐ�.�����6��B�y��L'%�J}wm����ײ&�i����O�M��* �0�n�[�k޸G�@�{+<�Y �-�� 7%"ǆ�*���Q����Ժ�a(R����!�x�� =�r˰x`y�`��9�400�l2ǭ�v\��0����>N���*m�pѸ����=�0�����Հxﻬ�6<�=d�M�/h���c�7wr�Q��!������g�
�DԈ�3�3�^}j�0��ȱ��{�b��(���UC��S��A?$�K�t��ß��Ʊ
Q��G�K�J�Eܨ�0U�nm�37s$�ʩ]��h�P ��vUt�NL�������ڹ^?=XD�/\ѻd�AI&;����g�;���>'F����]j�uZ4cl��	g����0z�C�ۛ��)�le�ܻ<��^�ۤ�i�d��Ͳ����7Zݎ9���K��q�(�j���;C��t�>�6�[���X~���@��gev����h�\��3�Ǘ�9m�:�c]�n�"�*�pb��Wg!�{jG�f#pi�V_�9��]n��N�!��8��x���[�k�B�jbL�^��̢�9�o=V2ǲ���v������Um���8j>���Y���w<��"���L��u]��IOd��	��ΚΩ.�m�{s�Tc�Z�#�fsD�;��V�^�X�3�C��_�Iu5�%�w�\$ I���?���]��1�v�F{��0�q{��௾}x4�{�|�nEw�o���\�Y�Em�_}�0�8�9��#;ޚ<ߦ���i�|:=����cys3LT�?0�fz��8&�R~ �y���k�}y��W�y�H�l��g*�P�@,��
�˳���W�$M�=��2�r�K�V[y��~��lh{��Z(�1yfl�k�4�I�Bv��߾�Q�z�k9:P =�8ЭC���TQp����*V������@6�d��G�ܾ�ۑ_�C����kz�N���Lp�Dvi��Bx}hz�"�WN��ր���2���ĞD�׋g<^yD���p�`�lx[�[��q]��=6�V읙�pqsq��:��_�~���A���,�ڌ����(�7�̥��h�n o���{v�b)�\|����@��m��Rh�GE�4�蛇3k7)+��W����.0�zUԥtK��	p���͎��P,x��~ka�K�sc*�n�@^rkj�\�c�`�m�KY���']�,VKUVs5ʫ��o�.�z��!�������7���*���T�aǿ�rfH˗��zH�p}=7�O�w�D�]ٝ;]���^F�v���r�X��pDh��Qz/��H�r�m:�9��e������y��uU�}���t��~ӵ=coٯ�)z��N�+j�,OvO_�{jz�7$JDW���02aa��R���v�� ������ԗ�.�:_�X���f��ko��
3m��W��yW�Z�Gw����*�D?U�nQ������"�7O<;S��w��^6-�ɞѫIn.7��-����ƾL�~�j`�D�	������|��-������c����G���[��AZ��U��������B�e9/0afs��x_U: ��n}�s��}���т���=U�5�z3g-�]�څ��;�G����%�1G#l�#���Vӓ��(���@z��|�p���_Rx�"�G.�P�CDƨfzJ5�⬅A|�u�!�ww	���[�Y��)\;�w>t�tT>�/(����Op9J���DN�����,�B��=]��%u�����Ġa��N\���6�����^��T��[�X�l���=}\�x�������Z�Þ�`�n���#C�
�^\���R$�7X>�`,R{ܱ��#d��;pq�nw���VX�A�ɻ����N��wb�N�]QY�@�[�w{ޠ|"9ݗN�u�#�fZrI�W���;&Mb�g��n1͡7K���6^�?���K2�2~��Y�7�}�}iڕ��p�u5�q�٘�W'�z��j�u����At�����`���E�;m����S���䣮�0T+���TX*�o+�<*���`��	��>��V]�ɹ� �?~���$��H��7!��=��rܬ��ڷu�£�%��[�b��j��^��2k�`�HqoN���ha��=�:��З$%��m��ւ��n� +��1�{\
��S�W��3 ����e�^�")掠�=*��X�����@����[v�<� ��w.�u�#����I�_`��Ώ��m�KuG��[Ar��V�M�C{/��

_�
��|�ax2�Ym�e��[�ڱ~�:Wh�yPw��5vܮ�{ʅ�ӆ�����Z�eݻ���`SU��C���{/l�j&K�!"@�HL�拲�Ю;,��=�{�]�u��ǶJ�i9�n��Ya��%5��o]1d�;j������U��-os\��"����f����+E���Æ\h"Tf㤊f�:��5���z�|��=�	�����He#��9pO������zv�7�3�7F��l)R�-	qL��8kNЅW���Ҡ���G�����|2����77�&�K�|�jg�d�&h-�'�(�B`�!�Ӈ����N����K�a��f_��ީ�7.fb�)��Y��}|k��z/z�y��	�~u��8���"���[��SS��r�����B�}��	��r��i�ɢ�s=�*�X|����c��#�vR�+��G�ک��Gry���hE}�Ӗ����y���#�5��Mz�R�������j��-%�G��wi��R�g9�{6N�	dR�@���I�Mۍ�=��+q[y�{v����(��2?�2A�f"�87,��&������7m��ьms���Z�î������م9�0�[�К�;O/��#��l�Y�įZN9�b�c�<��iۜ7���l�l�{k <�OIҘ랇�t�xW�;{%�Uإ6�K�fx�_l�t�cmH��u	��Q��m�m ��XU��uɸnm�78�����7ix1�E�:lMt��i��S]]j{��ѰYl�!�ƈ�$t�_������������H���mѯn����e�Z��hx�n�$�"�7�"ӌ�Љ�ؕ�Fߚ0��[ڲ���{q��8\�@�}M[s��X*21O[�Gw�'�{yxH�{,xhMF`-��l��f��5=#�ak�e"C�u����~>�T}�h`"�y���Pڡ�o�a�|1mn��˼�{��{�}�uԜi��Wf�:"����~C����U_Z&?s�+�[�K(��_D1>���+��2�Wn��r��@���[��lzgf�T:l*�9�.;u�	�ϳ������;�{{n��~��HY2#����2�%��L�xգQ˞���i��O����=k��H�bڎPp��
'�ov�������`�z�	�:߃?(`��<��IW'����LXu��Rr�p�Jr�V���@Q�B�E�-&�c����r��ѹ��۴���[��q��Ý��v��ް�.���uA�:�GX���)�n�gE��1`�����gZ��"S2i�x�_��.�HP�T/�/ؔ��ּ�<☀�當��H)�$,c|�L�Z��ӂ������:�5���/�"����N��:`;�.��>_h$��s�P�d�~���9����{li���L�"�j)r��?�~ϗ��չ7��qNZ��K'�d����/S�N�8k9n_\�5��ߴ�a�c"<�2'�8���}$e�7 uQ�$V��~ס��v��ah:��w��B�}0�{f��ڥ�#һ0t��+AA���t����"�H�H���Vy��yX���^���H���'<yI���:=tl�()�$>ʍ�v�o_A[a��y�RK�b��o՞��o��z3�JZss�d:p����F�����Sp:�Q0֎�D7��Z��N�)LU0���n�Ԍ[K���tաb�3��[ªOJ���H� �sI�j0b��1�Ԋ��y"{�����B"�����o+�W�Z�Wn\������S��j��]�E#زvm���9o+@��i;7�{��G�S��x��7��\G��;����������-�>�r�G�Ol���ER��2�08�1H����W:���e�T�V�#)�^��:*���V���WZ�0b�$��Ȟc��Z��>�#�u������y{��w����9\b��t��/y̴�C�$��2�4�Wu]mxb�B4��0�VK��!qb�?1��y�
�{J�}x�U�D 0*�����(���nI�s.;b��� ��;;v:��o#��+.7�r������M~��X�$O�k"l��+�y�*�0b{G���ԝ����Ms ���?X���p6%�3E�yu�}�	�o�z�Ba��/3���]�R��Mb��g+��//�Rf�!��g
Q�⍔�M��L��L~��v�_�b����"<���qsF�M4��~^���,cyi��a��e�̱٣��F�em��PZ�jW������;w�+�3û*�};���绯>d�~���\���Iq��%�-��UJ�sP��Ҹz15�������t���[�;�؀����/LE��O� �'"����N�9u�]��8V�f��6�>�m�_�X~]���1��Ÿ}p<3��s�<��	�$[K������;+��h��֮��V��0<�nOG��� R8�@`�Ix~�|��+)��EM�R������}{1p��*��{�k�z�ʾA֯Z��/�-2�.\!�c�%:v�%wmG�g|g;2�Wx�nL�|��}������r1�؝�+���i�����y�_�b<��F�Re�H4���������\%k?`m�-㙖�e��
�{ֲL2�J9�)�V�<7�X�3[Aj��,$�D�y��`u��^x&wE5��$�У@i�}�N��Γ[��e�Rs���Wj�vc=�L�}�w��6A[���D* �7����םw��*V��b�k�ս:�H���"C��o��)"�2���[��v%@R��z�3���c���ba/.)�$�z�
��1ݐSי�uc��Fvx��V"�����n���A��>�8ͽr"������v6�e�Ӂn,�J�Os#}�3Vn��h
��c$�ȝ-��&G�Flaڂ{�G���[ָ|Vc:�M�V��mMk):��*��ࢷ�[�vj�2��nc9��nȾ��q��WABf�(Қ)`)#1b��>��i���u˝��&��76��ӱ���󮼮��w7���	n�6.R<�����mˮ�i� gw!��uyP�X�OȦ�_�s��o4�f��֮��`.�Ɯ�j�ju����x��{�s��H����:�0�jMđ1c8h��88},mL���T�z�����L�N�.��E/Ԁ߲Źpd׾�6I��[���+���>����)²�K/V�j����-���3)�te�ڥ\�[Mu4��r�K�I��#y{��LP�ϋ4e�w�>˷N����OX�st�b��J׃v�R,T	���n������\
�ڢ��M&N�-�WF�k��*V+�.��e�+�/�X�U�Tfh�XB�+M{�Q�򐝓���.��x�P\�͸r�z����鞛7l�VS�>)��쓘�4.i2�on�.u/Foq�i$�0yӖ4�<q�7�;s��_�Fz]������
Ţ�[OM�t��+����̺�W��eۅ����2��N���p7�2��{7��t2�~�X{b�z�x�.�J�II"�FM�D�v5:����`�n��S�Z��p�!��^+2ٔ+ p�)AT�N�	�`���1բ�"�epl(��!����װ�&�W\@Pn���z�S�O�ە��L�G`ۈ���<�\\A��y0�M��6H1�������6�كoMA���{fT#��B�գv��-֫Vۮ�z74w7V�$$�17ec6��v���&�۶�^����0��]�o%�z��x-<��wg���5�n.�i;5��qG9�F�hc�i�[����<>-�8sؖ<�s��[n��mW2�^�1�8�f�u��wP����m�yx�>����K�=V|.	{>�õ��6���o@n��ck�ɯzۍ�;66�[(���W�rd�n+]�wgge^�Y���1�5�
�m�.�Lg�u�m�rm<k;�-�Yvg�� q���w��eh������]�8�,�<�og0�6眹�3�����Y��1�q���A�M��n��ta�ۑۆpp�w=N����0���=q�'������R����nj6D.�+%�g%=��ǭ��nB��O-vv;	�]�˫��h�9��-R�dp�������=��pyy�&�m�dНc���f�G\Jv;;��k�v�������<XՆj<��s���R�汭�ڹ��O]�{Z�b�83ƍ�+m�k�x��ݛ�n�;�eɇ\�Tq�w1���Ξ�ö��a�[c����Q�v-�͖ӻ+Ѹ��9�Z�Qrt��7Z��q����v�E��8�c�pYy���Ϝ.��f���t�ۍ��*xK�հg�&�ێ��sټ=�v��ɹ�&8�a99ڸ�#mƦ�xnܒ�zL����;�r�g��g���޲]s��<E�L��b�.u��ˢ���\d��[	���q';zH��ɍ�m��˔�Dk��[ڂ��␺�_/8���u�+�ݜ�f������9�f�.��ku�q6����U��]�n�5i:{-�;G�t���D�v6��0��9SԦ��T�j�ӯgR�p�J�v7i��q��^����쫧�t����k5�w=�/l-c���ka�����ᢧ��L��ܾ��mM���r-�=v�;p��Y�7R���WZɫN2�5cn��8��n�8�]���:������焷]�e�_]r�m����ls�����#ԝ��݈C����N�{N��_g6�-�$�C�
uһxI�V'<������`���0ٷ��D�s�F��Q��$�w����u��O]��:~�݀�.�n��f�b��X��7Ym>�3FsU}�d��g[����������f��Żo3/¤)��"��mv�˖q���y+�c�:wz�'sVxR��W��w٫t���1��A����>���.L��	��D�9��k���(W��HUn��k�ʇm�E��vF����r����{��S�;�<�B�ᗍ�w����Y�C�}�%a[y�,z
��4��"��ϥ�� b��z��S��|g+�n�~W]�7�P�gQo�A��HQ�O�93�"��
��v:�_,"���]�+G"��XC8k�'+��:�E[���Z�g����)?��9j��3�w<nȕ�RÂ�e��0��8]Y,��b\
1#!��#PT��2��kѾ8v�g���0�]{g�[{x��K5��-V:�9
�G_���=;����QC$0�S�>���"�'d�yZ}��N���ȂC��Mw�zR��\
���O�
����Rֹ�s�ۚ�7��;	���:�?�]�jX�����;��}��k�v�W 6���w����yˮ �R��0K��@QN4 )�y��X"�}ݕ+�M×TW��#�o���|<ح�7�A�������+핎"�oK�<���m(SJB37�=�q�U��yPY:?v
��PS[����{�f�Y�L�5���5'�,����2r�y�<b!0�.6CN;$��(Q]���Z�r(_=m�ʒO9��������1��� ��	c�W^�_��/����$����#��:k��k�59z��=��\��V�0�k���v���,+��S�M�"$�=�>��oo�V�{e`�(��>�ݗ2]}�y����=�z������u�*��q�q7��q��&G��(i$3��g{���e������*���&�}y��Ϋ>]~=��FV�UGL��N}gr�;oM��{X�]�*jTKK��B#�wm�݃j^򶜇�j��Z����2�Y���˰8��"ZH�r��.�HD�4��%����ܶn�'���hA���9TI>ZA������!Z+� �٧��3���}�;�ǽ�*-a�.@�q&�獏+O��������	��[�8���Ɛ������uag��%�{Ջ,⛡�h��|�Q#�R��E:������Y�f(�1{�M���:�)}s��v�5em�xV��sg;=ˏo�T�:�ءv\I}�1w�:���Wg3��*u�z�n��[���;�g�7mr_�Mfk30r��6��|�.O���>�*��*���;�ˣ�{�X�q=��V���kol��Q>�Z�V-Ƅm�#��3a��/�^�ۢ{ENK�t;�æ=j���o'yy��G"��
�Q�pVq�����P�3�2�a�Y��I���n )êvT�$B�ཅ;����J���e-�͢T�wd���x��˞
`�.�7E�%� X� ��.X�����̝��g�"1���S��Y�iΘ� �eG����GO���=t�N9Xbm���z�o�Kd+��۳w�b�C/��Kf��ܭ<>v73Z�v�L�����ri�3�Kg�h�j�|�)�T✛�����ܪ�c�f�٦3�V>VηL����<P�ﻖ����>�%�a��� ��Jǂ�J��� ��ӯ.N%�}[��c ��s��g�[�Ns<(�_���
&;��96o<�\�=ׂ�n6X�޾�{[^���e�c��i��Q~�8u��%R/��3A����:�7���<=��ޑ�
J1]لy��G��0]�{�頠cqK��Zw��
��1{�^�{ݞP�I��3
��R
7������+�;�C�tVK>���[z�z8F�G���Ÿ¥}��2d0�ILI�m�2�^�#�ǂR���1Vv��\\mO_S̝~�G�;�uw�Tu�t�����G=���pi�I���A�~	Q-c/�{.�N3��\�%ݎ�������n����G�(���CnҺf^�t��[S���o��m���t�e+y�ژ��`z�PY�,�^�0ȷ�s&u�#�r�D�6>[����ۣh����
E$���U�M)q��;v��^ы��7�x1�-���Y��<��u��|H�o\��n�+�*���j�v�`��g'd��nKd#�h�Cv�G��sG@F����|t��c;V��;D��u����/IWk���uIg��l��_lus�-��I�����4i3,p���qa���%�ṟ3.�{g�����Akm����u@��&ըݺ۬��d���9�2mr�oe�}��{�N�^۔b:��mls��k�3Mq	�*2O=\7A���8\>oiF�  �R��dX-ž��W�%���Q	p�^�&q���zl�䴗�$�l�CL94"���K�i����ȵx��[����Biypz����1�دuXͽ�A�
���Q��9�07R2�����yPh6B1vq�9`�w9�6!�|*�_؟Ms|:�q����b��Uy��h���H�-� �f}e��*�?o^���5c��w��z[�g.���OG��o�@)6F�^{x��ו}��OM7������V]�X����X�iON\-��%	]/Ƹ�OM�����s��?,�������m�7{s�/�M�: 6�X�H�Ey�n��q�68���N��)����V��r��;n�g4dc�8�m���Hg+�lܽb��}���YtF���W�f�	;�h�s���c�M�����F ��t���PUȎ;_��4䒚>�V����շ��Z$Y�;>N����~WsV����6c!���U��k�.�
D���Փ5�f�}���&On_��*��x.fWB-zI�e����#��{j��v��=�_�8q�-�@��l�g.kf�B��{�偬��ܳR�uC�^�p4��
5��a��.(����n�D�B���-�<���4��{��BwxM	����*x����2q*8� ��� K:M� !3+/�o�����A/P}��=�>Σ`���|�g���&!
.���+؇+&���Wvt��ק׶��������6����u�]˹�Wix��/"�̿�Y�G�9{��oָ�O=��OL۹B�<���ïݟ{t�����m������ȝCTD�"
R*�����,w-��ks&\ -�23|siOAX%/M�Y��6�l��3�>�W��:!������x� I�@���S
�N0��e_��(�������Sf�(�_L+`d'K;�ōB�:���J�c(S�B.;�u�N�vޚ�,b�+F��"'oWd:��*ejub��֧��M.]���ߖl&��[+��E#��M誧�#��:��׾z��H��fN����A��R��>���o)]�k!�.�8t�;�Iv6���!�("��S�ސ:&��K�i�����f1��fMe2I�o����2H�z&R�w���$t��^,��("��E%H�N���nδ�;��j�0h��rEuBQ��j�yf��� �i6����8����fVfr��-r�W���[.r+oV�x�S��*g�9Usك{X����L[!@SE!	��yq
�..�+��I9��F���>:�:-ovvd�&p�4���R�{ҳ/D�`o�h���PQ�$!6d�ٌ7Gg��<��@טu�Mƶs���jN���Um�WuIV)�h��Ӭ�B	��Le����e�`0ⴷ�62�O��jgM���x_1��[sg�E͸
�|u��w~hR���됬{"p��>[o�i��t�!̥6����Q�堲�f���;�:o0n�$ݮ��u�H��$~H�
I;~������Etb8q�l��������_��c��y���to'
�w�+�?	��O'�ۺ��C�ɡ�=yOzM01�xC_2a+�D�.7���`�ᮛZ�N{>͒.;=�6.��1[��9��ݐ8a����C1Ź��*�z�ɂ���Ă P���Ĺ��O�y�p��ǻ�#n��L�!����/04��Z*���A�:.�D>^s=�a��7����-�6E=�~޶Ee������HU�G~E~� i�JN�q����C�Eߠ�{h���,`S���^�]�z��%1(T	w�
WD�2.��~G���%�Ð�"�
/���sPI���&�����t�Om�pF�Qf���0s튟�y��=���3�8R1���I`�qI[���eVw?��Ku�g`yuo9o�P?��6����C��3đT�u0#9oX狻t�-:�X��bz%,���������]��/�N� �gr[4(�ې��y���Rν81Qf��	gU��Oq$���]�(v�E��jA�rȹ}��'r��6t�ϧ=q�ϱ���;].�b�dJx�e����<��s�eEx�������$;��	ty���qK�S���nA7oV�������N4��ۗt��s�{&�Tv����u�wT�En�Ӓ�܋u�6��V�l�sh}���p�8�`�b[p\� ��-0�ņ7�+l��p�7���m��]�<��;�s�����*iF��ç���cY7��z��㧫6�S�F��*��2�-�v�`���~���c�|1v=i�Z)�t��y*�������\w��=1�����&[ 秽0ـ��#�S�Ao �SN���0���u�n^{���=����X�s>b�wZ�7Y�u��7pz���u
�2�Q7��c�l^��d+�VE�U�֡O�S�͋�)��뱇FJ�ְ�P�c����O�I6
�R`�+7����i�/®}����:��c�x,hJ#M��[�J��=$�~k�g6?WG��pS=|��!�4le�c�H�|�?�PAJ���؂8�X�p�����Wy��5�A�kێϳ�с�p�ǈ����q�^�����mu��;;�nǞ�ݗDd2�t%�^NoF|G�#	��n$#�f9e�:�gq�������9[���~�:ᓆ�����Kro��+zk��]A�L�,�f�yߩ	��N>�j���H���X}��f��h���em�n�h��Ьo0c���	/)��ݰ�O2Y��%l��[}���4F��άn���w:�f����CD�v��%�}�jM��{�����˺��%��iXJB-ɜ&��Ś�.�Xl�p�Z�r�{��[�>��M�u�8߁{^bs��x~&��A
~Eg6�!���(�L[�����1+1�V@�v��>ti��ܿ��}��4p�n���9Y=�=�?f�p��h�`0A q9&[��ݗJ��Ȱ���uRS�܇��9�ǥA���k�������3cj�]Dm�*�'�Ee��$P���R�n�&g�d��#/�.�ڣH�i']94�14�F}#�r��u.�}���
�m{�:��ɱ=u~�=�j�hhFW�t�I��0����O*��I� �;�Rv��ǰzoM�w�Vd^��+޴2]i=�A���ۅB��Z�;��f!��>�}�Ӥ�<�P�#"Pt�	:�,y��z+���U&�\lI�/|��n7�:���[�T�X���#=���S�]�V	h�;��Zl,bV�϶$(ly�f�RQ��G���̤#�Uf�6��aW^eY��DMY&��põ��]���ɮ�P��XWZ��N;���'�|����h�����31�~ �T)�o�EY��תBw��=�V��%5
r�M�H����W�&�&j��4F:�l��t�L䫹5�M�ԃ�u��wZ�5ם9؊	h�4�4񮹷ƷCb�����wke�Y*�
a�a��f:�OF)!�'�����m��T���]��:�c4�R����:��r��g��b�d%��@��R�5��n��� `�ܝ3�)M�[��fc�*f@h�q�f�ec2;�Z����U�b��uX�E�S�<[�`ي��J��%��P-���{�P�.��o��~��7O����,����JS��PPdW`}���l=��v����Nr�2�ty,���27���.^΂�V�Z���7����Z�c���.H�i�[���kО[[�]S�����&��7���d�m8�ۘS�%���W�v�&��j�a��|�׀M�j+
���>�zq��+/��[��2q���Bl��9���h�d�r�e����:v<�Sa�h�Z�8�ֽGl8(q�9O�ԥV���YcmM�wK�')yk�G�����aF���~���8K���uʹ�S<�ZL��7���F�V��+�?�H����Y矧D�+���Ay�����>z����F�*�?M��1+n���;[��ߕ0�4CE0ې�!̡�~R��&pʴ`V;����H�g��;��hc�S����]}�g��.�ݯܝ���ٻ�.ع���wed���y6�����ҁ�$Ú۱5-����d29"ͥ��K�r��C��ųF�E=֯}�-�����
��-v.��l݊J�f�'�n�����ST�m�$�y��Gn������cxY���ڑ��V�N�p��Ͻ騜�wKe�a����ޱ@k��r�ګ�p"c-/���H)�y���kk��\%�뮧-d,�֩ږ�1�2wN}Z%s��xr�#�SԏhH�	I�a�:��Gz.觽@ޞį+���{�(k�O��.;��+�T�w��.�f�~�Mo���|й�l���K%r4��t�B�d)CS"����ɮ�ܭ;s���ke�v�x�)��U�EXO�K�bQn;�ݻ��M�?n�B;���=�p%:-������ʏ� �b�]��U��:�:���W�)��.�h��۟V5�����g9���!�^f\ˑ�\ƲG/ �3��7�ʌ��}��d�7r#��i�}և��o�u^��%�z�ML�/�<�Ʃ�|�1�PQĤ�۸�։��3�W˽�_i|/8�d�s�wE`G����H�O�]�m��2wn�[��Ǟ�wS��̬�,o$�f:���#s޶���uk�Y��Ṵo�-�|�g�od�J�x�Y}ǳq� MHw��K5!��d�-�YC�����ѭd�7;���@9�@c��U��=B 7iG[�gn�畇�"���`H6Y��r<�z�V���n�(���F�g�K=�uΦ�����S��o�^������z�����Z4��^k3Z�EN��j�"��oyF{:I��:u/�gL����aї�jA��/P��im]?|4:wyrń�׀�fF	��q�8�Ī���72������
�$̍KV�;ny���6�I���e�l�5����y9`��;�\&շ�㓆��a��M��ӛ=Kk��gi���MU��76n����sy��眕���۵ۃ-�ɹ���X^��Z;V����s �f���WVy���-/����l�'t6"�ػ���ي43)����6��mv��XLn@�ܘ8�n�y����פ��ls���v��,tf6	h& �j��S������b���y�,�婢o'X]�g�_�zw����龓*�֍;�x�p)Ih�������9C&{��� h��\�Ι3�ۗ5h�������rb�]}R"����c��Q|Љ�Y�ժ��l9ֶ�
����̉z��vޯu@/������+�:�˱��W$CT�(DK���aoC����vl��EUr�B����/�<�
/�����f���v����|��G��طV��P�E��3n<�w�%\���=~��cJ,��=�ڜ�ӆi�>��`�0�6���^�R��dJeĩ�8��-�`5�ktqo����O��=�D�E���i�O�Wn���V7i�Q�yaZ�����������EX���S�W���E���窥p3ii�&��yv�/*���T�7��,St�i���t����ԧX�q�Ctf{	���M�gqIgo_=�].@�,�P�T�Ə$29N�����q�c ���fK7|�0ͱku�O"#����,�b᛹8�˶+5�[����G~PV~(�b��WsFE	Q ��y���UqA��=o�E��yԲ�����['�.2pƟ{9���t���q}�Ǉ�ƪ��e� ����ѧÜ��ۗZvW4��̷:0���y���Z��=�٤zX�O��z��{��^^,���h���!$�!!�#�91��pK�c�6�l�W�*J�J�=���;����D'��y��-�G+-cn�p_+%>�v�.�����P��d��EՄX���r�>Zc�=��l�m�1280�	���k�y:&{�c>�ƍ�d��&3(`w���/|uL���j������X~���!�0�3񅨁H4oX�vJ��S&�Z9k.���X��!=ҥw��ǰȲ"�F���^;}�	LD������Y�	i��(�����w~���f��a��2r{ٵ`|�g^���!�]�� �'m�N"���Y��}V:�WbP�.;���q�aEuٶ��S��������x�L���	�|N��]s:p��=��T>9��u&݊�U��"`q��62��y �|vYZ�Nѹ���>��Ǽ��x
�Rp�c�����{{O_�y�J��%	���%#�������3�%��\����[�缚��0��m�e�v-ۈ.>��ie@x��6�������Rn�Sz��==;Y�|�ʼ�[^�r�q�s�68E K����B�9�v\Gѐ�������^���z'�ʂ�����f���x�z�D"�v.4ҍ(DA���Q�O�+�u�=��u޽��؎���}���ΰ֡��Ot��{^$�$&�X�K�g*$$����l�D"�6�"yf���޿e�N�6�:�Oǻ�������Ա��j�c��R�=�O��P�!�1����ڝ�-}`D����}k���K�z�7B凋lOz�i彟U{/EpW̆�ۀ�ᐚ�)�Yʎ��YӜX*�I~z:v���g���]��<o^�+X)^}��J�WtIҌe���sW�k�2slϙ��DE)O_��a��-�by��;V���um+t�<"�S{�zث��x�S"W%�'�Ҝ�y�;+yW����H�mz��Cs����˺�	��;T7,	8"����J"�#rO�7ar�u�����q���ߦ�k�m�K�܉Հ.���&p���Z~�jy�6�mqe�SE�Jl坶�}蕊)�3���\��&��گ�ht�{�v�Q�P]�d�3GKo:
��~zV��^�DH4|ARH��f� ,
��=�,��Hnj���b��]�9[�'��}k;�/J��\�$�p'>��N:ǜ&���O��ܞ~�k�_.�łm�{>��a�҇}i���.���W}b�ģ1�e7c����<��*׽[y���~a�"h3��
���]�p��'/bP\�g5�������z��L��#�`�y�ޚbr��Mwm���m�Y����uN�>���}x}V��G t����amA�N#AM�*���B�H���t<�{gU��0򽧶�̆���>G�n�c�����=X���Ǉ�Ԝ�vzkv�ѵf�e���6�3�n�
6�m���g��t�@+۫�7= ��6P��:�6r*�Λ�v����:�gw��s�;s�ۉK��3v41�֎�:�����-�X3�.m`����{m̢�dݧ9�CcZ��sA���8�q؝�]�x�V���-v�dBHz�,/^�{l7+#�ݮ��-ԠCW��j��m�]�r�8w���+ ��s�91[�+[�I�e;'����J�����\�G���Y��|^���Y�~��;"ۭ�S�b�ژ����y�U�z���i%�[����#� iײnW������O�a ِd�*�� B?y�Xm�4�_��Z-��`O�閵ߡ}{��M�>�4Q��=�2��7�(:孤p�"D��9=��ܢⴥ���=�u{�ھp�_z�c��6H�=^N�d�~y]Y�8�%�n�uuL��)��M��S���O�ns����g2��g����VNء<�%wL�1m�}�g/�r�1�'+������\�'������&dk�̱[�����nm�db:m���o�w��p��փk��f�-��^\���[����}�3}�羅خ]��`���n}u�DU'O �Wȭ�͢e��>��n��&�]��ˬQ���t�p_��$���y�5ڲ*cmk��9i,�X�zx\�HZo��+=�^,mֵI�I���̄[6���L0��=��u��"����u�}F5�����"ݾ&��Y�ޔz��=��)��Tqe�����F/��5?:Y���n��I���"�,�u������]����qi��r�P d�}�[�ܣ}}�YzS���>����w�^Ӽ�r���u��_<�PN��op�V:�6�Kh>T(e&�(<�C��Ҟ�Qn"�i�.�Y�ʜo���}���N�6���znd\UQ��$Ǐ`����ϳp�N���^l:�K�F�5��k7��aq8�@�" T���z=bǮu֝�d$M��k��~rn�p7�u�}��M�����K6��^&'�	��22X-���Jno_��߆_C7�.y�(�V�ͯ/C�N"\�`m���wt������w��2Fم�"NC�ޚ�wϽ��xE��O˳)R|\=/��[���vq����,���V����E5"��!f8���]��x�Z�[�*!��Jl��i:�_ܯ"�e;��%�aC<�����ȱ碄)+m:tE*i4ۚ�V=/ j�/x�ђiew\�0��X�ޫ�U���z�'zs�9A>KsS�=qVk��BM���|�n��큨��̼h}��48�^4�!���#�L����r��wy�b5���nc$�%���[<�DB�fs�G8`]^n�ݴ�C��Ұ�9�&e�TK��仵n�����7�澜��`�F�����=;��v�v�0n����T2�zP��� }���r".H��8n�ӛ�wl�|'�'������ܷ��_)Z��V�c]8���f�5㗵��յo���xE� w�L��.BH2Ii��̙�~�=gq���M��3�=��@��p�>C<�^����/9�\]i*�4I�CtM����]��d��.�7�@�~��5Pj�{^*u�����;3��"+g>�ܶe�Ioޞ{�y� ��f�P{�4�E�^鮈c�`έ��<Y��{A�ޭ���
V����{M�����	�7po���*'�2I�3l��2�kC���V�g�R��>._?Et�^�����P�V�ޖ3�bYY�w!7�/nn�J�	0j�ŷ(p�7i��G:U��c&N.��5�x.<v�(Rq��A8Q�.�ե��7��x�|��]J�{��v�Ҿ`#�m��[vxy��ޭ�o��(I+�[��-����J�t��7/���7�O v�B3�rИ����^��E�,����{[ڇ~��r�}���I����TQ�:�����t�W�����F�/L�0���|���k�w"&��ƻ�a�0�ђ!�B��Uv<#�tE����}+��|��._�E�/ޒ� �����s��lwI����@�X\"�!#j8�e`�nN�wy�6���w�XX����q�nua��U2��|rɃ�����jdԅ��c T7{�z���f�{�l=��Y=E-��qp\#����u5��f�K�53�uݱc�hw�˽�5[}�֟�3{$V�vV=]Ӵu����|L+of���;nIW�]s*@���#CnJ���=f@<|��b�	̹��G�v�C���so��K���ۼ��/\JN�����CN�D��J�+��B���{{�V�i�� 8on
]ٛ����l3UB���f�K ��B�+��V��weN���b�bV]t+!�c(S�<�Z]i�y�v�m��}�M�:��Gr>U;a���2��z�e5n��&ӄNCj����c`��m��Ժ�#���Q�xH/$]s�ޣO!����25��:��ǫf�c7�E�rЖY�#�\/�W6���[Wټ��_Vcw`.�x�kHx�G-�rv"�hU���o�0�
5-.�9�n�_5��ݹ��ҽ��~�x�^�e����O����:��������Z䷹�qo���J�;N��ǻ3���fu�ٔ��+ý�"|!�.�W=|{���Q�����$etY��K���n�ۤ��Ѡ�Y�{�EPz���P�C��W�f�W����}t6O��ݰ��v�X�tL�7�g#���20rـ�����R�r���|�v�cǵ���oi�y��r\h+4�=1V����D�(+�S��:Gj$\�9ug�w@;I�x`�oK�����9w�wu��^G-��4ķ*[���'
���J�f;FS��熒�"��@��;2D@�UUUUUR��RP��l*����P�tv�'��v���)��6�]mAň�gc����#������p[̎Ybɋv"�˼2+7=n�<�؎ܽ4l�.91��G,D��vm�5�1�eDz�:v�xћ��.C���Z�����`Ճ���/Ky4nu;�3jEm��9���ۥ�ec�/��i+u;���R��WH�B�M��Y�ۛ�pas�w�V
���&�0��9�bA�-0n�¥�\/i�s��o	�CnۍՔ{F݆�G��b5Lgs�8���lZ�m�nLn���n��+���6�Ey���g�O����ckZC�G���j���`v�8��-̏0I�Uwy��T J$ٸ�ek����p�8V2�r�p����s���)��ĺ�v��B��sͫ�w�m�%p�����GqN�܏[)��-�x^͇O@�Q�Y#�NK^�j;,p�^$�V!m�Y�[�����уu��;����<ݱ�v��z�!'��#o\!��F�{��cV�܉��u��/V0��z��Z�pqc��|c�=�.��NJ^��w5�sǗ��Hꧮ�w\n��I�=;�9(��9�#oZ^�ۜg�[����k�k�]aF�������]����r��j��n4�;of5��9���Y����]��6]�[s���qn��
�+�;p-���Zۛ�p��Kb7/1�m"ˆT�-q.�pc�s�kK�<�nq�����������X�]�����knN7���"nqi{+g���c��k�ӯWnw9�ȗ@v����瓵�����=t[���|��� ��Żyy�4�ļ��5���AV�uXs���;�};N�d�8�*	=YU�ƺ��n�>�M�5is�Ԟ��29�q��Β8���5�L�:�=7��X]���y�8�\�$�#�u���2�B݌��P(���0��'5��]�]T=�b�2= ��b�j
U�l�#�n�L�Խ�"��Es����9�tqŎdn���J��u�nnh�c�[&s'n�m����A��R�:@��Wn1s��u�����@�Y.��V�Y�r�c��Ft�uOsv�6��q�7[��rnꕘ�ZM���ZWOY2��t��U+j�F����"�Ş8����k:��g�N�B^���s���/m0h��ќ�����6b��iϫ���a�����Gj��2F㺝�=�m��<�tq���/9^N�nsB���i~S��`������5
��8�ye���.�V����`��|��S�T�'>B!��7ݸu��H�O��qD����y<�˜���S	�u���BU���4k��D�*|�l�Yo'q2˧��߇����/{.�5���ϖ�g������b)}=��⭭���O�B�`��.H��ziz��
l�����9=�*��zR��ǨTi�8yU���~�j�O����hz�9Vo�Qm6�;=��VC0��1W�����W%��K��I6��#̹�\���K��/�d�f^U�h�V%㤻s�d�wc�tp�m˓��������R%� ��zn��&�8�z_q��lR�
�t�>S�C���b�iɒ�G+_�ɵ@�+�p�H�2�D�@�d_	���\��C��ߕ���xm���@}y�M!�"Uy����Y��H�R;�_5�,�Y��$nC2�03�=����M��p7�SVSyX�d[�gV$T��{�kǊ��; �k�/�<G#�C28q4"R+�;���g}�����{s��B�R��#�T��u�5�q�*�U���cd�R0I�J�f<��^��W�0�>�w%gvPK�ԨF�c��U�3|��J�ڑ�M�8�߹f�#1�@vH�	Rp�d���1Gm.��e`h��t��:�{�m߇�I���	�&Mi��
���Շ��{NwgX?��&zA�x��j���&�8��o3c�s�{{��k�^������nƖ��U�ԥ�hC����(5���X��Z��'���^���~n6�Etw8e�Yu�ጳ#i��!I����f{����Cإ\×5Ƥ޽|3\r����ȫn�o+��������f'i4�|L�p&�n&#�%��i�mdU��v������O>��������L=H������**����g���0�˧�7U7�^�����jdч���d�5��cV���7ے�?Xf��-@��i���,�T���ڻ:�(�}�+��Y=��I�ݢ"���7-覈�U{�4D�~�˒���ʂD���y���`��N9��"�y�wb���k�~}���R|5���~u�m1z��������.vH,����*B]�av9�#�{vc�V.�w9�7G�U��l���X���Msh%FYq�������K�( ����qc�8j{��n��7ha�2���g��׹c�#��K� eț����[xۉ��B�C�2��Mt����*v�U��/TrXyq�˼�+�o�����|W�G��NB�A)K�{,��|��k�O.�~'�G�iNKv}�7�+ֵߜ�}���O�Ȼy I��BM�Xs+��g�e����ՌJ|_tA/��Z��1sX��~�Z�HF��v��a�ZkwK3e��o�VY�v�|7�����v��a�3d����n�J�v�sb�����b�7E�o]�C����鳯��2dɬ�t�#i�����kQ�A��VK��ί<U��^W�C�h��������s;������q=(��l4�#�b���dq��8�Iu�n�|e�y��[�R��rî����2�rᶲ@�?E�w�;o3/���ÔB��¹�ì�O>�5LL�(�[��D�8�U�gϊ�1^	Wuw�Z��u�j�z�Ǘ��_\�_��ۨ��euI�� f2A�L�z�۪�-җy<���Ʀ_���e��~e���Xݬ�^�5oX�	�G#Q�Sq�k�wq�{���ݿOt[>��m�;��F�;��Lo&�o^���O]-���l�����cG[%q�B�g"�­�����#��%Z�;��׳�Y��II���;]�r��u�`��kw��i:$.������k�X��y4����ƍ.{����7�V�+��T!��I*wao�k^w�;�c/,��qe���.]��Rk5��1�^5��]̀��ޛLot�s\[�7kbx��ټ�6�v䙸�v��yq�ގ�-�H�ںv,g�\쩍��j۞�2ո3��7ʦ3�;<�7C���Ƭ� pP�pZ�&�����0n�a��C�z�
yyG��ۣ�*f�˳��ŷG㌇[�Krf��r��v;�g��9훌X�T�եrm��x�現�R��0�yI�� �;t�vp�!t��n�KD��Y�b,HBb�DI!�'���mNw��x.�|1e$���?z���h��4'��kU�Ӌ�B\)��%�0`͎��E�/\V;��e� zwX���C�e{�5�����i\���{��GZ���r�;�bi��h�nCN�p��-��tv�hܤ{0J'�G5�A�!�����J��5�9�VX�� S�-ӧ�l�LRM�v�����gۆK���e��v�M�k"~g�rˀ�O.*��ⶤɵS6P�@xr=���HZ��9`�n�������h�}}2�*���%y�O�Rg���-��a:��^����U`�C�I#��� ����;�!���ڵt�:�4�z����G\U%�Q%&�F��mm'z* wqq���H:_fG�+u&N�eGρ��o����7=j�e-�>cj:7C�	�i0(��j`�(�S��3e%�����'٬��u+���]��.�1f+�@fS��N��僉�sZκ�� �m��(7N틽��+E5���Wj�ʻ�!�޴|��G�;��m�~<}���@g��P���\��3�+s+��{�{�Y�l�=��$!�ߧa�dY�{������w<ә�S�-t����Bh���$�v�S}��3��9t�yH�f�쨰l-b�U�}���G�슸b�xb��[�x�4�W�2R� �u����u�Y��͸5�קI��nr�ݹ���$��@إbe��i^X�W��?nV��d��L$z�(B�(�0w�H���ݹ�	�<�g�{':7:9�x���Ӱ6-�i�M��:8�c��+�ޞ�:JSGy��8�vh�N�]'��֩�&�o����Hi0�
G#ۗ�Qs|�}[�ۘ)@_�G�����x�)����JԚq�ff5B�P�}O��em��f��&An9$(��p�UgMѝ�T◄�~���;��1��v���W�=�	5�̳� ��<�nsO�8�n��l�5����'�oi5�y�cc:�s�\gQ����K���q��kr��qHB�q$d�$xSqΩ��,��e�Y�0I�ҭ��N�TzϮ	�<C��Z��zIJWv/�;���4C%�����y�D�t*zWx3ί�XDs���evmv���ض:�x�+�[���!kE>w���N���E��$r�0��on,�;6ԝ��we[�ku��N5u���Ƶ	�W/U� &�[J��ތ�^��IB޺�Ëj��;=�Sq~;�Ƙq�	��d�2�ά�N�rl���E�ar+7U��5���'�x�Ӓ��)�+��et��k����S[�K9z߅�Y:�!����FM�L��Ln(�N�w����Ha�#܎�ܶ'dvp�l����nb�f�%wc4��Y-E�o0d�����܆a������^��A]�F0r��n�*NA�3�+����,����PCn�%u�j���-���d�WPr��Ժ���5VI�I�4�Kׇ1=yB	���L�*�-/M�,�����4�j`Y�n{�9�QR�b�����I�Z�9K��϶�G�/z[��^j�������yȣ@�R$��h�T�:a/n�����ez�-��m��.�q�W+yy˫)���pD�I�!���:"B�v�`� {;���ۥ9>q�u-u2o#+/��n����y(�l�"�����u����̝{0m?��Bl��Fs2��®vq�.'��3�
U�*�F/��̪"��M-9Q4̎=��f��j��8=�8yy�r�׎\
�;��U������DW�{�: [I77�^�O+��K�ox6ձ�r��g���է˻ٻhz�@;��{��Ou�.VPӞ��l�����Ǿ(g_k�lź��s�|�[7OκS7���ó�W����VS�
	�����غ�uB�[w�}�g1b�.Q����~c	�dv*���N��m��c�%���@Q��ms\;�u�G�m���:�S�.^�li%r����盭pt�{p�����*ۇsI���u�����a�n�i�q�]�D�<�#���+����m�)�pv�h���9�ϒ�6�(8���n��}�ݦ.�1�cF��<��r��z<k�{xT1�#/V|��g��k��<7a�CXt��������N��ײ8����m1������k��q&�Og���[dKm������c�38��N�m�C���E���J7�ځ��g�2�OC���\�YjA�~�Pn�W���L�##
o�ܺ=�[�ُ	4���}�c����}j�+�����-�$�oM2wU�����M�^�^��ؖ�U����#M>�*��ɵ�w3���}���Ɣ�D��� �6�h&�k2�IFn��<>�)yy[{9bfv z\��ۮ�C۵��Sûۗw&���:x+-Z��k,�ӭÁ�ߠ(>-�S�Z��],��ř�[G:Z>������l|e��=A�MM�@�[,�i� 	���֝�_�,��hr��ioG黗9��i���m��C�'�2�f��ݽCx��m����0Cn3!	D�m��xx�k�3�.�GG@8�M�f�9r�룮�q�.�4n���+ǝڶW��v���͘\{�;غ@�ߓT�׹t�gNje%{�"|� �����+6ʀv�<�����Өӿk�P>��fo�X�{v�ᩬ��d��O�����&�۷��!�f�9��7V�H�(�tV��+����yLp�?t6��|-�]�t�)E
e�eM�r+��	{<��e�YY�j�u���u�ar@��DH��:�ƴ�6swY�'�l�m�{ӽ۷PfT[8�u'���{��Y�kwV��67Zth"8��5#H�]�!�t�+�k3�)���W�^��w�V��\O�/�|��c+�N��tx��;�����G,5��>��T2)&�Ϥ���f���ܯ>�Իz�
c"�r��=����Wm���C��xV1��uC���}Wǩ���̸�ۑ0�"���fX��2N#jJ��r\��ڧ�<G+��6��7[b{\�9���WIY�qu�Ǧ�;9o�e2���\��ᮼ�Z�=n�����e�6��X9�"'�3�s��AA{����+e���S��Ҝ_��uwQ:*�u���K�&GՕ�%n��Q�i����$umQOs�-̬���r��g<V�e��c]�_%�v��H`�W�j]e��r^�F����E�-NM�w��#P��d�{^M���S+�!�g��%��&-�}��p�gP��؝h�]J��`�*�`<��=�l�H=���Y"º�v��$
�[����	,z�>��#7^�����a�9\+s:�Sl&�a�g��:N�r�Gu�nZ�*|�h����w���2CyV��z�>׆��Wp�j�q�r�k�Z4��v�^�B��]Qo�-�Εv���b�;�E&�r��"�w<˸Kܔq@��P���봴fɊ^��(^�חx��"�u��w_:��P��E+��r:n��e�f�mY<ܾv�Wa�y��|n����̺5��UBa]�m��g�֕�-�]�3�R.���r�[ٔ�i$	�3@��`������<�����-�˿/(�!��2?1Oc��*Ҥ��?{�v�1�+%����<�]��H*-}7]�/JN�vP��qQ��kZh�`��k:Iܐ�f��Ւ3�D2�8��3��hzC��n^����c�s���g��ڐ�&����LGsa*����={ߔK�r�x�(�7:�i��ELDQ��;��YP���mmn�x�.�m^�5�"���ڙn��I;�j��tJ�s
�x^���IX��V��k������62�C70�%�i��kNm�ƌv�s�XTI�_a�rP�"��r��z�����`Џ���)�%�wr��Q�ne�*�t�:�M9c��w�}���`�w�e^P��*\�"�H�����w�=λ�J��`�ǉq������t��_S�,h�"ڷ�d�^���zh�Ҭ�W�W��q��ZM�`�i-���M�󽝰k�����-}R�Ww���J�m��z�Μk a�^ݾ~�pB�$'�$aH��żkg��m���ɌnM-`uɤ�ǀy�^#��dH���JC��z���]�n�x���}�,��/�oc6�<]�d���;I<~�W�ȵ��Er�E"�Q�a��~&�d]�=6W���G����l��1-뜱��h��<<�5�3Cfh%�����|�E$�4��w;g?R��M}n��O��֊�+D�s�k˯�v e�y1�3SI���L�D�R���r;Њ��k��Y�԰��Y�q:�h���yc���7�#��M(�fQ7���V/K�ֲIJڝ+7U�:�u^T��9%�`c-�J�{u��F��Ꝣ�Ɣ��vG���6�tYʮ�͔8��C��ֹ̓<�����}�7O�=��XP���p_�m4��/^��}�hY]���!>�K�F�0�0��J�axp�\�m���q� �W��q�]��7[���\�^-�[�$�X���}9�ݹu�3;���&��u�@����#��?*n�[۔�f���c�.a3/ow>��>�g���'e=�sm�GC�x�_q�B�a���}�t�;�.^�øT�έ��S���F�:2�!�	mŏ!���+����]�X��
��"�-�T�ĉ�꾱�`]̀U04Ȥ��2J����z�c���B�����??-�}�����s;e���f��Z*�^?Y�W<{�G�)	�)"	H76Ћ-�w-���G����7'�Ǌ���n)���P��[إ�i��'�ƹh�;���rY�5�s9خ��m�E@�l�#����F�U@5Zk45�������`��]>S�8���p��.�M�'<���h�;�Q0IF�J6�%(�:j��Dǭ���tv�|ORb=Ktu��)�i�nm���P�#pcľ�2q�ҌrcN)�4:A��tA<t�B��.��܎8������ە��ݡa�����$����+ �=����*���7{UXw===ve7�#'</��V�u�i�3q:��7�i���Ox7#�ͷ�ۮ=s1'u��Şǣ]`�o�����vJ�W:3j�b2U��E��g'.n�����&����\��h�䓩����}���o�~����ݣs�P��a
U�u�+�;n�����z�O;r��PU�\=��\-�A�a�꾧Ƴ����y�}]�N�ηS#����ݑ�fc�}��{��Yr_��2�q��R
�v�SD�E�˄*>�r�Z0K�LS��=��� b��/_uy`��ÌF@�N&Č��0�N粌���XZw�'/�oG�` %���;3������1�z겻8X����]�Zh%�&�H�I�Xļ�7�_sY����ʗ�QsDd��Z{�i{��G�U������r�ޘd��!�Z�Pm�n�κ6{���8��[��4VxR��m��Bl!��Fܛ��&S�;K��/*��gT;�x��"J�#��ߴ�{<m���C���\��#2&IM�ɜ���,���.���0X��ۢK�.��f������0���a�	��;�܄��Q���E)��mf�{ıF��MY1^1'3���v���{��it[׼��n�m�(]��#J/,O�T�6�jA���]�P/~��t�$���W*ztU�˻�+�u={�F�h�^�|�E�@H��`�m��xn.��>�j����{�H���Yu��>����s�Dz�w��o9�|n�%�)�È����Lqa�N�{9�B�C��V����;�X�r������j�7�`���K���Y�-�L��wue�2v��ӆ燈P�u8<p��N+Uq���s��Ϝ� �p�
9ov��y�d;�����{Qd�����^�~��s�v�F�Se2 6w�V�Bt|�ogs��{3qo���~���h���'�
��ݻ��P���Ř.���l��L6��eke�;o�>��Z�>~^�pY����/>�Wӯ)ܥ7��:ں��%$o��J�̢��c�v4����C�ce����`���A�~�c��_��Ո���ct�Bdj&)ɫs��()i�X����:Y�en=����O ��	�$���f��ZH>!(�e�;�-�գ�ټd/r[������u�>��a�z��;����T���X�pɵ:�:�؆(H��Q�|�����kt۞�<�S�C��u�ŵA�9Ʒ���l\S��Q��v�V��g���ؕ첻݆���9�p�݃m�y���ks71Ow�n�Y) C�&���C(�>y��E��/O�͞T3/�6�ԋ�+w'��b��O�x9�������!����1��HH��K3a^�vh�;�7��V��7b)����N��O7�Ro�l��a��K�N'ԓ
�m�!f'Zw��t�d�4�g����^��-Q��]�ij�<�۞��ӕ��׫t�;
q%�d_g��.R�b-�9e_ewf��1�J2+��iTQP���w�+PK�os���N��
��ѥ�8Sq����ddF�����w]Lᢆ��::f�c^]l��e�f5����w�����u��w�M����7�����L�1[�Ķ��;��y[�=�];9�$�sw\�j)�\L+$:D���u��{8z!�}.n�a��}N�ݜ�h./d�W��_��y秹�rz.��f\��������mט�>��>����Х�HTk;�U�#��^����*�s��	^�U=�~+�W!��#t5%7��܏A�~�d]W�*�2j��7�u;	{Pd�/��tȍ������1����-������*��E���yv��ޡ��=����n E������y�����U�v�� �a�JX2�%/x�H���2��^��6�c���I)ک��j+���<IWEV��EP�Q�5��77@�1Y����J���m�2{�d�w�r{}Z9E�m%(Z�9L���f�ёsm]J��iz���3I�m���N$�)O�&�R��=���PON�;�och���uC�l��n��<�lV����]��sG%�����cB���v5m�����x�m�1B��ˬ��cv`�q�qd���Go.�pq�n:�#��κ@6��� &�OWa�ƍ'=Z'[��m���<�'���*1�۫�����U�Vx<����nۜ宄�� d�Cd���\�=rv���kN��:ױ����Vw�B�1q�n:��s=��b�M���ث�DRq��l1Q�����?KYegwc���۫��T�ܱ�{6k� ��|�_�{ܖia�v]���-�Ҍ!B#�����ӻ�g�ζ�C^Y�(�Wڵu+�]�0����Ejd��+��
���7C�SuiU�jZ��~�Cy,��ʒ��2Ӛ���+է��X����Č�ӌ�#	B�of�>
���S�9�m��/u���5��sy���`��sE��W���K6�<�	̮�*�L��A�D���]�Z���v=cv�+ٽ�GW��z��y����o}�nX�v(���}[~cK]9�>̻�o�c%����3$��yxݦab���R�c��z;a��]�Lt��ky�	�f8����G�{O]�ԆV}P���Z-\���8Kٯ7-����KSw��	�`�����M%nF���v�J����YyG�#��v2�ٕ��%7B�K��hcF�S,�}�qn\6v���)!]-�Vg$E��$x����#���ɾ@RHj��Unw;�T�ʶ$޿1J���e%��1���A��{��g�^��/ch�\��rE��M紉[�|���z��9�u�e�x_X����xڛ��ll�_T��"Hｚ|'� �U�ۖ�S;�yA�񘼽o�&�[`�aFe�RU���~s������2�C$�3$���3c���Azm��l��zrV���r��g�R"�U����%1��@[HB�e��ڷ�S���B�Ts�⮗ŝɮ8��M���F�jKq� f9𵯩�Qz?u��6��~ׄwV}���;�}ke��85��"/m�*�
(�\ש������5J�(�3챙��<{w�g���?����>�Uq�%1^��ݒ�W�*�H`k�a���l��m�Q���A��+�A�Oh]�̧ʴ��_��']`9q�&3YD�`ej/2�5FHkwvr���J�y��c�*r�,Q�/��A7i�e����l.�
39^��@ ���w|���8�A�.$�:=K<���������ɮ���b�k]i��ٝe�;���{�b-�YiVX|�5y�zfr���thwsM&A���%cxv/���~{s��D+��LEӔ�<zs��R����1w[��a��\�;k�J�7D�^�^�&�Mػ'vj����F���e�{I�i�̾�w4�0�Z+~N�g|߯�+ȟN�x.�����w�]��-�/A�,��Ƕ��1ԢL�h�I�	��YS���j�&J�Iq�٘�T�֐r���a�����!�6>�T��M���т�>n6�m#$!	�*�-;�/�v���8�9�*�D��[�}��S�~U�v0�.�6�b�J�4�a��|[�]w�OtվI�3ܲA�u˹�,k�{"�y�h�OJ��̉�׎��$m�}wt�J���	��#T/F���lN�R�������q��<��͛�嵍��V5�ސ^�����{o��Tl8�m2b0�9��C��x�aV;C^�Ș�x{%������78���v]�f�4�LF�e���%C�x�e�m�cx)�xd�/Zy�9�)����F��/d��u'h�<�H�A�$�7�^���H�o���;p:�6�.�����zT</��\o���sU*��W�L�rnf���� �yJ>�j�U���-p��ٵѫ�..��{�+�r�(�d1^f���!��G
(I�4�ug2�Q����5��Tn#H�0S�1wc����v,w�yn�f1����(���I��l)���~������6cώz҃o��|�������3��O���/�}���'�K�XEM�ɬ9��g����*Ԭ�ȵ�)�R�����u���L����7���QY����hU�6�օ�z
y��w�c��R/�nk�uu�~}�Lk�����7g9��{�Y�ޥ�Źu�"�޻J��S+&X�s;d[���ϩC{V�����;)<��P\y�c�'E��Z��(L̄P���m��	��5궀��odu�����,YA5�{,�Z���՚����[����2�fW�21n�=�rw&*p_N�;���S���R�"�)�!D�К������7��*ֶo��Rt�v���̜*��\�m�k"��;^^S@0gn�{�"�B�*>���ݪ�;y\Z�zv��1rΗ����^�Jۉ�f��a��^,�Ug��Lh�"8l^�Z��W�_���!��=�Q[ktq�ig�SwZZ�֚�11������&Ĕ�b��Ǝr�!��a�y��>�S^g[�K^���`�2�y��J�}:<�ݸ����Kz5���I.��4�Λ�N����%k�;�o�{i9onK֝�k�f��甀�х�VR�R�6�A&Q�V�j/���V���7��z ��WX9�ϕYm�ɇ�_;�΁����|�譬������]����1�d�f�����p= Ӛg nΊF݅ϲ�Ëji��͎���Qh��;�!�;�Au�{���(P�K܎�eջ�z��٭h��[��Ba��ޗ��7�͹v:ݎ l�C*�Z�)�Lr�8���瘻�2h��ܥs_�,߽Y�mHNl	L��-&˻ce��-
��YE�U��S{0:�ɣj%����@v1��UUURDғhx���;�ھ��=�ECf�G����c�u���z�Mcl@8�q�d�� ڶ`�r��̑1�d�	�H8fSyj�v0��cnc%�j1� �W��7���b#�I���1n�䳠�^�3i�v�|0�J/Z��F[K�p�7#�n�[q���շ��
vS������4VX�n̝�y�+�봾ۑW�4��Xۣy�4kQ��&q���cct�#qYp�].�˒䕺�;���pMG"[��D��a��{m�n��v��ԇ.��n�V�)�����ݎ-��%v�{Zy�>�M��9�/jnM����nM��r]�8ө�u�6̆�=���u��F՜���X�:�ӷ<�{L��e��۩�z�vŷN�ڽ���ǫ���ccz�՝nmx+Q=a�Cc�z�x��TN�.y���W��\��:L����vg��N�\k��ț���8:���u�v��'�]̼mу�G��h|rq�������nt=��n6��u�;��٪^۶5��}�	��Q�غ:�Fy\�s��|����˻w=@\�Y�']U�/kv�6Î7@���:�n�1r��c��1�g��OD��c�WL�n�hm������C��\+��e-v�=���K�F�6�ݔ<�[yѸ��P2��U���ɮ��b�L{3㮻%m�W!\����fsȯ����6vɴ �.,�gs#���/eM�	��5 ��XN��1�v9���]�yx��:w�5�k�����Sv��x�>L�is��@�-�.sv,磎���,>xw	ؼ��{Z=�V���ݵ;��<g�ͱ�v�]�����m�;�f
%�l�%ے10[������m�2']����'<zV�Höb��۴ѡn%�M� ������N�bt�P���b�a�h�1�w���.A�cW��%�!vݦ(����Kv��V;uV�<n�'%�]a�Wu�Y�{�m˭�e�K��ݬϤ�sPs�4ۗ�q�b��@��d��k�b��[VJ�lx��^CR6�L���
x���R㩦��ջtc3`���XH㤋\��x���unȾ�j,��n��E�����l���$ǲb��*G	��b���e��Zn�Z)ǲ<Zq+�k�cQ=����'��i�rѶ��s.�A8"ו56X��x�<h�۫��ۨ�[E���#�\P;y�<t�ё��p�rK`�9f׍��J=�=����@�Pc����
�`C��!�y�ߩs�ڟ�5��������;D�yދ��A��_ڦ�ZjyZ��R�3�p�Sf6�'$1\y<��K�Bv8͉�aNr��^�`z��)�ˋـ�q���_�|���tsݪ3�R0���AZ�	�J�)�eK+��0:��iGqot����o�ɴEofd�A	�tmU�1�⾴Ö��x�	��B�LCt&��U�}�Xuׅ����K=xso�IƇ�X�e��\��X��~�ƼDHbf(�)z}�:�]��̨PLqL9�Z�H��y��5�q��ʽ;׃}�G<$ڜ�}�2M��y��q�r��8���;o5r�q��q�J8}�nk�����b�wU��~ �`>���F��2�^~�d�M����m5��%�*���g��{q�̵x�1�v�L%��R"����MH���fǹir(����t˸��Ԗl��}��e@��Uhb5Ӹ�IhTR_Pg�==Y���w��Z�����x�<�1�|�&���`���p9=ݯ9��7�����h��t��z�ݻ��Q�CC!ID#M�r:5{QW�o�+������]���m��f?c���9H��\;�B�M�F�m1�+��YY}��Ak]����=Yv{�؄N_)wt���/2����o1>��1�CmF�j�NA�S���K� �}%:á�WtkN�Sʱ��U꾄ܹ�j�ɇ4g���c�@u/�[.q�c17h�ݹ��z.(�BֲZ�b6��07WKnmS���=z��f��9ާ�cƆ�u���=۔�x=�(��Dtu��#� {V�dE�d�$���*''u��T��ӆ�ts<�%�a�O/��Yμ����C������^����S?s�F����W�fK��֫��Wm<�����/����c,w+5�Řд3A}~�*^m%����3�&oLK��{�	rG�"WW��#�to��2]�E�L��)f*��a�3:tl����L�m�y�p6�0�e�ٳ���c/�'��X�nx��{(�gyf]T�m�,���+��!�~�h{^{��2�k��1���(��-��׈��3S�b���j�AuAv{����T#D���쳳ov�@��Õ6��4�ߒA)	��%�wE2�}<�X�9M6\v1K���˰\q�y퇠�%0�(Б����x�ǌ+��#�y~�$����L�zW�R߶�Z�ם��a���]p����� �-FeX�o����m�����DtOWu�px�z���P������wXp�T�&��b��"F�P�d�"��߼��\��_��J㬩��^�������yjm�.q�S��+OQ�K �|�&�iI#ɶ0����K�=�ڪ,���5Y��O�1�.���
#�i;k�ܖ��]�p˧��{�)�����#�<\�2���i���1�0�a�,�
w��G�Zp#�V�{V�;6ڗN�zW�<��e7I�NK���9��m�+'������t�VLё��Ze�y^�x�J�{�����l>����{�6�����p�"�����:E891�:)�nŢwK[��%�\n�Ǳͷ,?8�H"!��rJǾ���wk�[j��<�
�K��d���פz���-WG�<;7tkDR�՘V�_�n*)�~�01Kg����Χ-����f�+mI�N�nǔ5������h�`�>���$β���r����h��-�I��G�hZ��2�j^����ލ��32��ՈϗnA�9��m�2��X�E
�O`�5M��Q�[��lf?���l�l̒Ѓ!����+�L�/�{Hh�۝�wݖ�4�=�;���u��7.6����h��i�}��ˌ@��6vZ�{�cǭK٦SSݎ�Έ'Ou���I+��K�U��Mn&�����[���@�B�+.z<f%�;C�6������FZ�0�Qsr�ڹ<4��󵖝�Ғ�҅P���t1�箫F��hՑ��N#�[s��r�W#�r\^1�Ĳ�r)/����C$���<���p��\alp[Iظ�m�m���,�6N��Wۜ�#$��󎶺�d㝝Ō�c�����Cŀ�\�XC�8=�ٲɰ�/c1r�]�6v.M4�bV���v�Z��}��v���P)�	�m�F6ȫ��dޝ�ss�S�lp=�N�#��ķ+p������L�����Nսs��5�PtS��x�7?ۮ�1W�߄�g-�����y͛M�Y�O�����Χ�4=�1l��u���Ax=���7��r��NJ<�>�y<%ϑ��܄]w\�d��"b��}�B�Rr#��&�_�>˱��!]D�M�����c��+=o��Ǖ$/�܆��o�;��Ńg��Oǐ��{�Bc��x���b��=VA�"��4Jr]���oq�|��]髝q��2P��fy
�w�'Eػ�^^���Þ�w��2X�[
�e�c��ܯ����[k�����H�
o\�m�f�X����t�u�(����}w��0�xB&X]��3-.�=�Ӷ��^20�1ghC���zSr�\ܷ]qÂ�I٦v��>�&���1����:��Y�	���H;6ng��'����;-d���b	A�h�i��h`�}���dltDπ�켚s�wb�`Ν��1�Uc���W�]\!A}�r��'�6�����2�\T�*pU}�[�K�+��������(�������o�2�yn�'S�_US��Ow����ɤL���f����=�AM�NYͤ<xi?1��S��l���w���A�]2�-�q X��\�b�2�;�XQh��zG[�����U�r#��ʂ�}��s�� 0|����Ϡt�]�e���lw�6ZRH��fI��織�yg�k;�Ωk�m8�u�K0�u�=T��+|��SKH�(�7�EA1��W�d�ֲb��F8k���f9��/L�q����a���/�$rN�F�P}}k+��v�<G�|ޮ\61}w�|��r��3|��p�#����[R��$��A��v_1m�䥩Ox��{y��#��25t�K��_-�b�ҏ�b�^4��>�����"�g��
i��棈��ޡKɴ���}fw;ݬ�s�z*7�.�_v�N�q*��Z�D��ck����'Wn9����=������u,亴������Q��8�*=�UC!���K�e���&�{yׯ6�E��m0S�%#ʃ3M�Ǡ��˓Zf�\��X\���}4w]���7Z�����\��F���gK��G$�6�V��d�zs{�Z;��C�{"����aT�;z?�,�v��^�lV0Nr���C$h$���ڝv���	^�9W��x��;��m����f��s$��8T2Gʶo+��f�"���ܯ��P�gu���J?\�[�����/|��������#!'��%6�Uù^�z�Ħ����V�{^�T��٭;�hķ��IFv�
�y#�4�����ǻğz#��$�8"�B�����!�����"V�%��n�WY����w���:y��6��{�0�W�3�,y5Ѡ�j�͹8y�T�*�>�Ѫȯ�������m
���hKٮ��^�K7YY���0L�֟e=Ӏn7}f8��B�B�N2Lt5O�#Ur��a����ѳ�ja�|�@V�w��"���yVuV�Z����6#o���G����d�%�%/X&&���Y�@���*��c6S�k�|�X�2ԩ�DlkXR�K��k��T�>Ŝ3�{���㞀,3T��u;vE����9u�mTf��l��frFQ�ݭӵD�p�d�qYt�ڥө�����L;�)�x���r��Kx�h�;3+=�l��R�g:7�T��bݑ $N�A�3sq_.5�l��8��7��2�'Q�����v���w�,_����r�֝w*#���9h����#�ISM�o�3HRU)��4�喽���49���D��s���+ى!�u�d�1fO�L���"ID�,���J��G�X}����X� �ܮ^��v���K��SU��v�\�µ�J��p��d�1�!q8�ꚶ����U�6��ֵ粝��o�z[*"��yh�t@�����ǁf�Ι�=b*ך�����s�iV��sbw|�yo�Whi��;y��u�O7(m(��Zr�Z�������=�*3�i�@��ڜ��:��:��Om�����ƚ:m<�Dg�"�ls)�j��rs���nrݫی�j���v��l��������Y0n�B�	v�s��I�cLo��{D�J��s]<���Lvr��l�ۙ����\]��^�v��\��*�8�M\v��;��,U��I=n[��]��乤�^��ǭ;(��!`'�J�N#��<�J�#o\G�ak����<�Y]]�s �r�f�(Xl�����p�.�1)x���1���s�����Ou�˻��2��G.HQ���KOO;���x�_g.��HI/��W�x�w�� q�)ꮙw��>�޾��N^�0���c#H��o啦m]�c���}�~t6{�IK������bX]Y�~�x�gR�H���
�a���!D6�x{��ӈ���!��Mhfu���	7�r;|n��w�\��	��"���u��Ѭ�R����'ٗvIk2����u�e���v�e;��~��1���C��Y�M�ڱ���o;/S�8���L�������W}wf�D��P�j{[n:��S���i,�Zz*�#���`Vro�`���%��f�v&�nڟo ��^��b�'�^CE�7gB�5P�mu��p��oi>!�i�E��L�r{�k7��f;�A��r�����\ͥZ@�O�E��kSn�I���/'
9.C,=܂g���=ϰo%�G�f��U�fn�P�{�ٲH������pt�yX�̞��v�7��Z:��fO���RAaN1�v�+F��/%�;�#��D=2{Ǩ"6�߻(��iAy[�hF�dƢR ��7�Iʢ~i8�*����w��/�&��M��u2*�ݚ�z�z/V�k��M�da�s�$��K��O^�s(�4	s}<�.B��H{�t������y�Ҋ���+B�´u�=�>�]o(}	p"AP4�����['��ܦⷵ�Wdx�y2���4�\,�BF�nO���:��lѓO��΍�ީ�n����S=���׫o��3A����n�.M����i���'�=:��n�O{-�y�Ó��`����э5y�R'��r�o9V��"�QM='�(�i��!��y�\����1�B���-[{�����iWw�=��+r8$^;= �c�)=�Z9m�<���4�*�ZY�6ᣲbx��F��U��f��)�}6��$օ���,&z��ͬ�i������[�^{'�w�������Vlس�n�:��6$�u�Z�U�W���x�%�Y� E44,�	�ȕ�Ȇ*s&"~�iWn�9�TYq�t��+.�w�S��^}�)��,=h��ث��8������G�P�\�$[�1��5+N��Kr������]�7j����ֱ%��1�|�Ӈl\)�yu��Iz5qU��Sh�6`��aP�~������Z+}��g�;Ee���G(ot�؂a�yV�e�^�6�\JՆ�z���SLE�Ѥ�m� �z���w��j&fs���R��u�\ՙ2B�ୱ��1�nѿ���ϼ�S�X^�NC����ߞ\k.�K�.Љ�]NUΚ]��m�W��n��)py�c]#4�9����KOc!]N@#�h Nna����װvα��M}N���� ��͕1��[H��s��)��^�tr�b�.�v<D�D���T������y3.m�m�kY�H;������=���\�n����z��lt�r�9�3DQ��ʻ�1v�H�j�k�&dx)�.��� ���k
W���i��ؼ[�܇�/ċ�u�ASs���:����߲�Q�����S��;�\����,�KP5W:avp�}U�G땱 u��*���Ƹ�>��Mx�|���Dq��������1۷Ec���K����i�_}7~�'�>t��"�79 ��.�/w�OZy�����~�Y�S�{��#H����^o�-�c"���&+�:xP	b�.H��j[��w��Ȟ��b�[�;K{��4#h$�AQ���`:E��ƴ�<��<�Ӟ���(��ahw�v���ul�\E���8ϻy����J������gB�\-�+0�'��tiLa�B���o�e���E�g�;�ܛ�>! ��yL=^�O<'��Ԩ�ӫun�{}l?�s�W���:��^���`�xFB����m�X��wN$Y�㼮Ɨ��_+˩CW����y팴�[����T`Y�c&�*Iy���֞yp��wP�Ɋ��%>��+�v�1XU�&���X�e�3��Gn�`k�n����1�J����[��&J`;������;w니a�2;���1��S1���!{�xH�?M,�Ξ�t�??�(T	����h�Ϝ"��J��T�^k�5��w����t�{��Eή�b�1�)�o�-�$R1��TY�w��C�Yn1�����8�.ڃu������r˩�� W�.,�f���~Cu������.��(�yV�Nn����W�W�t���/XO=���U�@Oϙ�%��k��e���cvz��9vb�(�-�z�y׵p9fq��}L�$�]�^��������o4�(���)� �*����Y�o�d��{t���$&��s!��x',�|2�2��gkj�S�ȕ�3cF�oM{������^R�K�N���b�w���iЮ��C7KԾ��P���`�{�t��!~w���_K�S"k�k���ƳW͠��?~W�2H��4b�_֖X,|E`�1��~�j��L<~A�`��k��n~�,�s�O�"�A��c7u}��P+�O�^��*�  ��߶�u����k�yZ��O*d����Q���s3�a�z�0�چ)��񡺑�˦��v�umλfvwt�/���R��na����ZP�"��"�kg)ή��S��i�mWm����4��z�n0��\�W1�:����/A۞��(�8r�Avi97Z�Z.m׬����=�<����\n}�n��n�k��q��
s�a7�_q������b�:�gv��Ň�φɒ�D�#������=tpEج^85�W���qN��ѻDm�v�ŬIϵ! ��]��M���!�]�n|��&�g�ͺ���Q�[���rI��_���9���;�����N���x�%j����ex�O�!^AH?_�ʇt�{uG�퉟��;?\����D�؇걬�"������/3X�z6�s�m�y���8�~2�l`ds}>��B^��D�א�=I�O���R��|Ï��!yL�4?~�Mh���Ew�ﮌ�~��B|����J��b��K˻�����H�`��[�ߵ�u� }8�������:����Gm&�w�4-��)y+���Y�vW2�c�o�6~��2��G1əz:�ԑ�Уs�}xY'��O�ԡ����K��P�C�Iմ�q�)Y��`����CWɚ�[����ڤS�xk��&^*�hCEf7���x����HD��#��
?��]V]�"�,�!��|�=z* �W9�׺���nW��^�Z�� C}�_���H�����}����h�d
w�pi��Ƒ������]D�1���0W�]n��jx����)�w:y
�9ضٳ�,]Si&��Փ&�5fuA��w��G�,�Rڀ�MwOԨf�����j8Z���ţ�� V3}�J���{�n��?w�J��5q`���J���u|�<��6�ݸ�f+/e�8']�0�����W�@�-��K�������7W7l`�Ș�+yb�*���d}@�Z�[57q��v�=�3x���.X,�6�V�{[W����]6hD�ҙ�����~~�_׾�h��c5�fY��g]w�i_�������?�2���1,gX���f�6�f��� �""�f9�'���x��gD�������-���9ͺ��+��,����^˧h����-�J�0����~n��B���7���_�$Ή
�$rf�"�VDՙ�}5pu���y���3= �0�/�g{U�h��� ���Vǿ�k��~c� �f�߮O�����$F�C��4B�.�@���a���97I;i~�
�?W��AC5}B�K��Lm��q����!_�`�KH���ϿJ~�4��*"t��W,x�5}�n�#�����c8��2bV�V���_wɹ1�uB�u�n�Rq�g������%ۓ i�dFC?�PAJ���,�?���˿�����ҁ��x+$�����w�|I�\E9�ܯ҇q��E��	iCS�;���f�dli�C�ire���^e���q�I�4�9��~��̴�?w��\+�/�
����~���G��LXE~ي���xԑfȗ�ߝO3�iy}||��ݭ��~]v؞l�h��H��������	*#F~���#,h�$<*m��Z�ng�et���.�~x�;W��S�"D���m�p�J(����"]IoX�H����������_���f��~��0�4=�1P�_����
?G��W�r��삘�8����	��eɒLə7�<�K�����6eOE&���Ԩ~9��,��>�u�?:��,�{����ï�AǈX�_�ק�z���#�n�u!E�Qdt���4����' ���8*��g~����gu��~?>ܰ���=����솓�z2�?~T3����n�RhA^~�n�#p�������ǽH��شZ�J/�P\Hձ�:t��ێ5h�u��EW^\(�]e��@�pFL��#�#�}����B�����\�ƿa��I���9�U7� ����(Z�EF6�N���O=��j���s9�+�/%s�;l�g������i���M�0Ȯ���ŝ.WV3�T�/w�?L�},0nfᔰ�²������ϸW��W� B�߿(^��R�ʝ��:wZ(���\
ݾ���i6Á���4�Th��Z��w�*Ɲ(��]����|�Y.u]'��|xzp~��^Ү$V
0��El�ߌ��>�7���jCµ_C���m�,��F�z8���ς��?���V�����.�#횪ó[~�u~�3�O�����w��͟*[{~M����ۃ*�>��X=3�˴����?h4���<WR�s�d˭L?�5�j���W����oVGi(޶�S��H�p"���]�����@��*�9�9��>a3&\mrܙ�ï]+^ѣ���h��4�b��
ѵ��>���V�;�~��)ۿԁ�]?f?X��X���?/����T,��b����W1m~����9=Ɠ,�%��Yw0c8��rnz� ��K�6�L`��ܢk`��JL�CG.��-���ͿG#�����o��ϼy����o�8MG�ߠ�|��*5���`�����OA��n����b#�qcE�G�۸n���V��X<e��ǌ����&d���;��n/��1dOʿnU��F���{�O���m>�R_���U��*�s͝ �����0�~�.Ɵ�ƑE�u��V�w�6h���97l$?~��7�C�!��]{�nL��&ɘ䙘o��#��0��WO�Ɯ;�7���piq�����=��t��5!2�W�1??	��8v�B$�c�~��j���'��P�"�^�??����^&Eˆ^e��H��t�E���֊.�_���<"�: ��/��诎�0�u3Em���~�x����V+�.1���P�?{}֐8��X��q�z�Z�s��.�G�pU�2�lx�ט`��ܳDEV��R����N�ɨgi�է��ڃ���Tޮ���~��n1�1�.0v�g�߳P���"j���8����F�D�O����!�kMHUZ�Q�,�3l0GA��u�z5�m��4}&V ���4,��Umg�:99�n���!�F�8����UUS�n�n��؈����R=������v��U�؍�O5�JZ��Vlq��7,��f\:�83�X�sa�'<�u���ld !=�]� ��3��[�Y1��!���55q�]Z�p�����l��p�e�ӻzuϞz�6ۛas�y��'V�ۭ)glnz��s�'V���Z��
V�+w6*�𸥒EV����q\.�.�#���qU�ύ���9y���5��i34(��.z�++6qt�Kvv틱��ۦ�B�Ire���}�&��i�[&���p�����N~����-o�Mu�!w�j����:�~'�^#��};��CZY/�ߕ�A�{���b}���3Y�a��2(�m��o�DS�8�����Y�����.�=c���('۪�}ھ��H��U��ʕ�Y"�F�@�1�j�_�*ΐ����o���ڳ�wQ�~�+���gY>��q�[�>�9s_v�1<�{^X�,[AA����h��ߕ��V����mܲx7f���@�&�6(�׻��(���x����Z���d���$�[y�32�y��Hgx_���}��ȥy}�3�!Z0�B��t��J��������� �f~6(�(]��;����_���:���~�_9�A �N����Q�_��c�2�	$�E"���ܔE�94w7&u��W��L���}c���Y���#<�q���5�J55��׮��-^jGsFIC����^(�)hJv>��d�뒢����߷��Y0n�u��b9A�����&����� �F��`t��О�s�¦X��1K��{��E�>`��?g�~��μf4����c�~�Y(w4ѣ��hI߳M���+۰�8m[^�<{�2L-�0����X�S����&�*��ԐE?�¢I(i�\��}���8G�Y��B�f�oX�;+���}���gQ���DFEk8��1��n)s��WC����;�Z[�Sy���^I�����p��+���3�f�W�~�Fa�6�����~��aв@�L4������Ŵh�l�G�����"HԊ���߽�;����]r��odM�& T����F�#��톆'S��P��^�{�{M��1����7��?���?_�tt����GA͢)�����%���nSDh��a��ȃm�2G_g��ނ�����~������G�߮vI�`�h�Qy�G�+�ʳ�#��(0�aY����*�z��Z��A�#?f�hiv���Z�������yl&[2�c/�^��V�ɑ�$���y�i'!��:K�C��ߜr�Z�^?!�q�0lf��ժ�5�:�r����#/o��Ց��`�E>xh���K���vo�2�N�pH�d��Nx���3�G+zラ� ��nӧ��5����J8:�v�N��������Ĥ#U����v(�pĆ������P�d����2�G�k��lj���}��.#3z�g#�,��g=T4���_l���kt���cnd�2��m���@������lY��;�_*�Ӻ���E@���U?G�R���m�4PXv w���ugG[F�}<��eϔ��.�j��V3�e�o��?�3F�/���1n���N����
�I�_�n����r)��u�)x�;�h?1�q"����+~��~�����xyo�Q=�_}�湲�WҏeM���m�VE��ǻz�j�[CH����=qL�X��_:¦�Vh /2�N���w ������u;gl��A�i|����1sr�2�fa�+� �D@�A�[���fX����|�~y�a6U�I:��(0_w�ZM��iei��BP��U��K����p0h]�|�K����R[���U,#�r�a�;#/1��O�~{�lȸ�̵��L�f��G�|�>��랑t��݁b���g�p�qg��T�A�P�r~f$k&\T��k����&���$�v]~u��0�m�uh/R ����mO"}��T����%���p��3.�+v��Mv���u�Fruλj�P��iy8�kv ��p��#m ,�t	D e~��0a��GW��i���֨-_kY���D��}�ף{�xE�����[�����R&*E��"� P�lh#	 ����7����s�K%�N�r]vJ�)�a�sv����ƽDR��3��O�?���)�ü�b�b�^��=^�+��ɒmo������~O4/�o��?B���dsS�߁ ���'�(�D��+�?ȝH�g$Mݼ_�b���
W�?���[�U2���R�J�D.���٫�&mv��/��G�Ò"�&N׳M���JH�A�~�ڋOٔn!5���`�E������"��}�N��eB���?1�@i��������@ń)Z��F��U'���*���pI�u\�����F~���uQ(i�����o^ _]��52��m�q�x�����L�%�l�mٸ[���b�2�1�ٚ��0
�gL�g{�ot6Vu�&���S�%�|����G�>�������?e�F�r��Z�_e�	�{��:���������$W���C���f������/�����_���u3�SAZ��]��yIjF$��$�"�_�������.1�e$�bەyw�����c͓̻���t��z�,`��n���殮-����s/30������v�c�s�'6�׿�7H;��%����wd�<������A:��Y�U񳙝�[n>=�!���h!U�H��7��*ϊ2�$3��&�~u���K�sn�fY�~��I��t�0����?�9'�߻�q�$�#�z`���X'��d C �D���.���4��A�3�+5 H+E�~��x�
:��S���E���.�LVf^��d�r\b=y�,;"�������־�����b�j���g�x]�@)~=';���y5P~W}�8��хENo��V�씫]�{%,{s�
{]��ot�)�A��-/dͶ���=��3�r^G$2ff�JzG�ܳ%�y<^=ߤ^c��ܐ�Q'����'�ʷ����AMI��^~�ݚ�(w���v�䉹�����!������#鍇gn"��-Nf�;� --s���z'-IKJw�%��9"���s�칣2c.�L3%��K�!6����P�B�Z7 �ܸO~�fE�N�DH� ��J}��'}������w�d3��FV��}�G��m���'!�d�⨊���rQA�Pq�(��Pd�PzErJ(?PELb����(=��袃�(��(�ԔPq�(9Eb�袃�QA�PkP����)���r����0(�� H ��1�|�g*�.��V�l��;[���ٙ��\���-)p�:ѣ��gm� ٻ���*����xMy���+�]�` iJt
����T��E��5Cl�E�ق�UB J�	U
IWL��U%A%
t�J�J Z�}_       ��s�J��ٗ�sU^��mv���SkWf��s�2 U*@�Z`   � ��   ��y{� =C!���������袅���lQ�V�DE���/y�����-��vp6�v�=ơ٢px�y�W�]vܛ�:�Kek�Zz�PV�]�k�Sݒs�-�[�=�J��R�%(USf��o{y^�[�\�[{�V���uw��w�{=��{M������砠�����<;Ǟ�3Y]]�]�T��w������8�X��w��V�{޷���[���u��;hz��^����ݷ����^x$���a�P�UTշ�����y�6j��޽����%�;C��M�T���7T�oz���ݹ����Շ���^�K���m���{�n���ڻ{��wmz��޽�s���n��x��l�mޙ�/6�=��v�����R��R�QIU*��o^ު�ݩ��^��k���)n�W�^��S����I�l�Z��knd�k��[k��y��.ՇuM룠)u��m�ݡݜ��n�y�m�m�ow7W{Rw��g{޵�^��w�뛻oM��nҔ�)��HB��D����vԯw;{��w��ٷ�rʽ[��z��a������ڵz�{s׳��v����<{��6թֽ�F��kҽ�e׬�s��=�g�y�=ׯkw�˽�Vy�v��=��D�}6�;��m��QR��/g�駛��^�^��z��]��ڼꩻ�=��Y��������N�MU���wNvr�w���n��y�s۷[j�o��]ީ�S۽�p<�w;����V�{���F}����&v��U�}�u�[2�{n�w�������5�c%��m�g��ޚ���w�={[���Ԕ۷j͋�jג�����{�{�����n�K�����������[��d��[����������T�*�QB��f�qw������w�{�v���^p�]�[�ޛ��=��z����׮u�{����v���B�l������������v�]��^�{=��׽�KiUJ�)P�"�%]�W��a�z��ʳַorټ�ڢ/ni]���ǅ����^ڗ�n�w��-���:��[��w��z;������W^m�K�n�����n�=��5�J%�U�$D�ٮ�Mv����m���x��M��ۺ�;���r+��a׫�f��h�wvR�����ۻ̡݉�l�s����5��k��u�[���{���u�͌�̪����S��mLُ ")�&ҥT � S��$��@ 4 ����Sj���   E?��  � �������z�`�	4�$����=5z�6S��������������˙/v;Xe��E��r���y����z���	 I0������$	 I;����$	 I?�@���?� @��B�$����$��@$�$�b�q ~@YAE�
BE�X �b*0YQQ�"0U������i �"���
Y �����w��R,dAV �*��Z�oU��5�i��I�s(��c6�3��=�){�t´+zEz�ؐ�z�3z��kT���IDQUV"���QU�@FM����C����w�g���������)�j��)n�U}�¤T��O�K�]��k�*@K���d8��8�J��7���ow=��27`"t"u͒j��a�,嬝]i��'O.�<�9�[��3_S��Iًhܵ�
J����V�j��!�*�Tn�HT7>���V
�J�r$X=4�&>ڊ�/�4�-Nj����^�չ�6��~;)����w�֟��'Ι�>�\[ϕd���>�Yf��j��F��C_RBؐ�rR�_���VfeVM����Z�c�~�,hW�Mv��]Z�`�6-WP@��X�O�1+:�q�Y�q�kC�ˣcB��mQu���*�(1[uo#5P�N�|�fT��m~�8�ɹ�yk?w[�1�9�O��+�l�N~t*�]̨��̬T��o/[h�ч� ��`�Ci�W�qެ�Em��F*�V �2�W�!�?�t����Dj�I�5�!F�>���{!��y}*�<i����>�/]TN��b�R�]g��z�g1��Ʒ�ɡW�y�WMحX|����F
��/���LP�n�P��uӎK�k:h�������m��W���.僯�u��Gvl����� ���i�z��ں8ti��E��F�sS5��GN�I�v���f�����#�%�nSjS���T�x�$�P[3�K�L��ᙇJ$Wuq�L�U�Y�
��_��]�0KT6r?>[����k x�^T�uvi��Uc>0S�I��I�$F�c�a���{�����`��dQ7��sMY��+Dʩ�ſ}�3���]f5[Y�5Ij����P��Ee:�T��)�E�Y%U�ũ��I�����
�[��;�V�IJ@�wU����6����{�M2E�,X��ϳ\�֟s2�FAI�(�����gn��ӝռ�W�5�ݷ�/y����;���wp0CI2Ij�q���Hu�}k�$0}��+2��PfQ��Ղ�UE���6��k�;�ÜﳧO>pw�m��|���x�x��o<��8��b�<����	�p<8����e�a3�d�y���D��u#���m$��r0�5V]͚V��<j�;X����ЫL������m���(�m�/��H�2
 1U�ETu����Z�;�{]�}`����)�����-�cZ4&ڕ{��	����`��~|E�
��t�
��nS���`��	\S0�ΚI&���Uc:8_a�Lv�<߉R�S�m�ى)�嶲b�F��-/k��W_�]��&�ӥ��щ,u<������=7H�����xW�)�a �,�4R�Lҷ1�N8��S��*�6���`�tw-c` 4�	�WGF+�.`N�������m]�� �jA�4�5M⚜ʶ""EDPD=�����в|�Ԩ��5�Vv� �U� u��-F��(#�,㳔�H-�u�j@Da��ꪼ�ĺ�V՚��N�i!P�E�Ϲ�5�o��k�;o�uݹ}��_Mo���v�}�vPJ U𼸷m��f� Q.�{yl+&�ilL�8`�A��-��cW9Rfo>枳;�ot��Nfw~�3	�b*��X�b�X�� ��PP`�"���gsW:���F���̤��M��8��n�Ke�(���¬�v۵{�=[��21��l���ѐ��0�ѩ�]

���Q([�
H�`�2�@ݩ�nd�uLx-�5�ekX�Su�&��k�3uV�C��)0�)"�X)PEH����QR�b+4@P�H�*��#QT�`���EX�*��"�(�,AA�
")Dc*��Q`�A�b��+�TX+E��1��Ł�y��f��޸�)bh��B�iT*�`(����i&)�c-ԉ׭��CvT��ܳXn��9�
��Hx���XH�Q���ֵ *�٦짡4�]����c�{v���{Ksl˭vD`���UAg$f\��P������fڧb��V���	�^w��kYMYP���x�a��ӇEZ�wm��5JYvE�����kk]���j�
�r���x�Y�.��J���N7%�]=��{{�T@ҍ�co	��7P��^3�]ì��դ7m��X.�*mCq]Em��h��
w$r����#u�G7,"�1"��F��9�)�e��r��{D���`��='K�����uCV���+F��_��Z� !��3�X��MC1k_��:�+Fx.�<�3�h�,K���#����ZN2��+R%��,�*)��f�z��Y�E�,n�A��[0l[�����Q��
�b��Ko.㰅^hi�N�tu]�
1�V�*�V�Փ�uM,2pG�2��HQ�R,�	��t)�n�F3�-�r�9h�j�1'2��Am��K�s`ţ^j���x�*Lj�0\(�e�"v~HLv3N�P�2����r%�Tu��ܼ�^7a��a�xh�,��\Q+W{e�� �Y����]+��?O��[oum�,S�ʖ2�X_���\#^H_���S�"��˴$8�i����"���Z)i�C��q�Iֈ-j�M��,�,xԋ���"�h�Z�X����U&�c��q:�T9I� �yM�K%��QD��L��#v��S4��2�Ae��%�);��7W�1 ӻ�a	�JtJ��Q���u���Μ���L��ݕ2V��J�*��؅���O%�E�F�BV��H����lMnٴ(�ݫHH�J��j;�:u����)mb
���W"���a݋��1bF�L.�/o,���m
*����:RP"ě@�`S+ Yu�&j	�����9w��������T������Y'L�����&�aq���X)��A�X�%-�2��3��`�1�S�sD�������6���T,<GkV�Jk�.���<��o��i��oD�0H+>�̙�Jy7�P����JeD�Lo0XK���,L ���X�3lV�ǯp)���zU=W�q�Z6�B�(8�T�J��F�,����V+��Y2�������HU��Gw9WY�̭��jqdX�Eue�{�^5��嬈M�(�˘�]��m�ߐ��YeK��k�������>��͙�`T'^���y!�1�M$��{��(���o�r�Tp�'��H��@Ћm�$a�w��zs�ߵ�{�ڨT�h#��b����EIP<¢�!�J���+��ޕq�%#�+$���F�e��,��ıe\�ᰶ���xV����ܐ�4 B�(X��uK�,ڴ%�L�	b�Y�^�7j�(����{������7�z�ĥ�@�����I�B���MZKܛ fQzC�ˀ9U�z�S��Y�62/a���м0=O@$~��
Ch��
�j*��U��b)Ĩ��b�*����m�R���%gUj�e�<ʓl�4��F>B���b/)V	iU���CI!R���gRd;�C��6�dĆ�:�y!��q!�C�*Hi��Xivڕ�]ox�S��Nn��������l[(��EQ��HgRQ7i�k#�C��
�Hr�
]�(���(�:��Hy�N��y�c��f[Ԃ�T�J�8��d`������x��feiX¯U��$jݓ�c@����Bke׳4Gh���������:���kw��}z�!�qb�L�.�ER�R
3L��>�u�8�ƥ����([�����Vu]%�^Ď����t���ƳY㹻d�*�^f�ѐ���U��ܽ�Dȳq�6l�8�:9��җP�gc��\��`i�e�bC���j絮PTi�6�VѦ���A7{��L��2Ɲ����o])�oh̊��2��`�VR[B�)B�)�V$aشς�B�,�h�B�+Q�`{����P�U"�,X�\�"�5g�������LӍ�oz�³0(MܛܛD2�ײ)e���T-�J1��4�+"i/��4[51�t����%'r
�ƕ��y��ݓ~����lTr��ѵ#����м��Q�c�*3fUB�lA�.�1yWW��vi�Pm`z�X�y�Um�<��� [Pb�?~d �$~"���b�Mc?��
v��ޒirħ����Vn6�=T�E�3M����9,2�/���ae�2���m4�Wt���N}��p�5�[�d�B޷�,Ksu�e訶�����.��$IJd9��cc��w�Mw�;F���͐K��lʻB��J��5��
�oT ���42]n<��۩F�S�N�$�M ��5)n��(����b&�9�E9f�ݘͽ�N�(�Q�#����F��]���(]�5a6��"k
UAS��f�a�����m�l�ɭ͔��2�م�%��Oo353��
U�d-�l�N�uP)h��/,\�Ȏ�����H�E˦�(iJ�_Y��W2�3g4|�
�ط$�@�y��]*<M<3FZ`R$��V �m�0��݈F���7̽�܄бUU�	Q@X1R
*1b�E"񒨊���DTT��""��G7�o6縻�臭���h0�=Uy�//?YC�)f/��ͩOoO�2Lt�yt�+5��R&�9n��@���d��8��or�h�@<se���u��ff�R���1��y��"���m�1قΛN�]�7AYyS�FhL�fA`ԢF8%�</0n��'m�X�(�ii'J⥛
IGb�P��w��1�i����og7�o���٨��VKE;�eYX$��n3z��(6�����Q����nLn�1(�8Um
U�r�J,���:��:C@�h�i�7�z���!��W�H�<r�3�)�%KX���50l�*��V3�u��Ŵ��SB��Lpν��6�yn�Y����0�����z�h�pVcL�U�;l�[l�B��Fc6v�d[J�QҳCokU{7d�r�[^��n~@B?;H ��6�ւ���2�UJsӜ�CMb���tY�+/��%;��ĵ��Z�"Ni�L'j��+Y��re)���pYPQtq��&�3d�@[.�էN����uC[�k�R�ͳW ���MQ�'�A��?m
n�;��l��_�BM��Xk7@�A3�m���ǥ�R�T Z	ک��Qb_���4�pY��qm�X\�	��	��u�ĕ�%=6Q�Ddy���w�{9�:�>޲�'XՐ�4����8�Y$1��ݰ��bm+ y��Ci��D8���V"A`w\ә��ޝo/����y�P̇XHu��C��aR��$�*H$4��C��W��{g;�bq6��EP�œM�f��*�㱯k���m�m�kH�cB�x�ͬ�����T4/�?��:�l��m��I6�j�o�p�	��%��l0K�[I&�m�Yi��m���]$�m��--$�m�II�m�I��m��m�D��I2I|�6�m��m�[m�K��i$�-��HJ$��I�L�H��Ki6C��Qh��H���]6�A��i'D��t�m�m�4�I0�I��H�Ҧ�d���n&�i��M���)N�l[`4��m$�m��D"�I�l��%��I3�]��n�x���Vp}sH.���Rc�9}[��}��C�:����XE^Vո���s�+n��'oGu��1u>�F��v�l�`e��B"��2��Rঙ� G��v��ì���v/�Jќ��q�Ǡ�D�S�=B�]�c�����p;��r��aџ��vu5�*�P��8/T5�o3p��	]:�O��]��-y�
U�2�7]�V�
��BG�zuEz�)��{�82�[���_Ј���0kY��V� �D���� �W�z�����]��H�J�wyP���\m$+���F5���,�/�*����f���"ţ�MX��gn��Ⱥ��i3��i� #:�"�{'F�ޔ���f_��-���K����n�x�=�����`9�]��+��:�����t��#�؂��woc�����f���Q�]6Wm�b���ظk��d��yb�f;w՝D�������`c00h1lԣ���i�b���v֫(Sm	���92G8�_b���	k3�wM��|��p�6n[����<������`��כ��(�u��H�'�uyDEy�(PyӺ����p��P�3iQ�U����&�s�K��n>řʳy�x���`�\݊s�`���S��*�N�(�m,X�6'*�	��y�j��s��r����ME:��P�c��r�HN�F�2�H�n����J����*I�CW��*7����#�Uą�+��2�k���Y���(h�k�{�l�|�^�Z�Vkl�XĠ5}\!��H{���C��Ր<�	쎸��<YE�҆��Y��ΐ����E]�&��K�'��Ìd�S�;B�7Ů״sr��'\�G�)��[C)C](�-I%MB:畃���0��\ue#6Ƌ��[k����-�|�5��<f�d[`	�fo6���6a�WP�t�<��7W˭��P�ks,=�L�uyz�[����ʾ�g�t1Y��rf��N橙�����Jm��ǷF�qPh(�r���b�w/���]j����F�q�L��Sjd�7@*���A�ȩ3L��4r�fR�ɹ�;�6��ú�_eW=6��*���Q��l��k��6a�x{me{�W4]�Ny�a��C#��+{6�ftX���S`�������>E!�+�mm�%�F�Y�i}u/��gv��s+�R��\��]p/m��G\"Rþ�V�"n� bȖ�VLcI4���[cD�im�<i��s�^�S�]���i>���+��](jpގ���8-C��R�\����`����,�爂FT����y�Xxv�Oy�yLC�ʴ]=V��	���z{N�Y9�����İZo��cmi�([�C�j
H8[甘�}�t�u��ʼ1����J�@NK�>��6^d�2+]�s�˭2pV��r�˩賣Czr���5���7l=��)$̵�q���*��]�=:��w��X�-x�1����7��ɴVFy��]�U���cZC��)�!�Xt�(Yo*��&�n�%Y���e�oUڨC�ȦK�lw�R�Uѻ<m�`�b�a���oi�n����Q�p#c�Q3g�AI��l�Ļ��m�L=�9�9R�)'E\�TJ���-�W�
�����O<aˏ�\���:"3��#w#9����]Y2�����������)]o���4X(
wiv�As[9]�I���ɭ�e�]@��:َG�@�]���Lv��?�X��rN�1�n��[m��u�u����D�.�/%{gz:1!\����-沼N�Բ,��]S��U�$�T#�1��cJYw���E ���cqR�:\�e��:��FG��I&3h�k������q�% 6r�Δ� ��f1dS�p�Y��η����3E���qaz?b����]��mֶe_[1sݩD�2`�2�e�e�V:4
������ɹk ��������H���������-9��L���,>�l�J�U{4jʙ���TUmc2&K����bx3\�CX�.�!.�Ѡ�CW���j���GI�"n4e��8��Ʃ�t��a�bF�at������.pPa���5����4����4�"f���O�����;}|9�A�C�9�'����ӛI��ud�u����a:b���a�"˽Mݢ?NY���i� ��.`<�'��@k]�w���"pm�vNC&3��e�D�mvt��+Ehd�3��CK���t�Ó��7�1��Ft|%�q67/�Y��p�%���X���b�z�1C m��܁i2Wmۥ,]j��.ܩ���w�m�E��.�	�T����q�n����!GhPJ�6��w�oq���/wND%�:b:Y�Ҹ�;\AJ�n�42�=\j��	)J�t%�ۜ�3�Yp��-��e��Nq猭!�i�m䳖�t��k�:4P�ID��A`�or��ws�Ps�0�(�o��p�ʶz-7H+;^��tL�^�dũ!���������`�����˜u-�nP�����r� ��5�ï���4[c]w�:U�����=���#[��B\�(Rbe�'	�$(fd��;�SޝA�Ҙ�5eҾ�nj�$�p읹�A��@K��b� ��(�E��ѫ�69�щ�����ȡ��m*&q�-��\�k;��4��!ܻC���M���@����xm���B>�=U��,/�h8���"-UQe!.g`�WU�~@�4�7u�uoQ��w1N�����lw�W"��ShѥY*��avw._���ݦ,!���, ����3����7�@�	��gJ�����.��v_κ�iVs�E�[�Tݱ�)Pt�J�0��J�V��G�+k�*��s5�Ւ\ݡ��i(�V*�t>6� �N���X嗚h���X�P����"�{ߘ�]�'J���3z:]�%7�s�Ք|��fᙑ�X��:Q�$W������ܼ�Iʽ�F�kj��sF=�MGLV]� I"Ƅ�
<;k Ht��W͞s��N�`*��'v�n�튰u�K.z$o�>F�qR�P5�]v�Tхts�#P�W��+v�d�z�D�PA�5���g��X{�s��{h�+7|t]����Y"���S�e�1v. L�}vK`��
);�]�����9\>�"�����n�	����T(�	a�M}�G���!ȼTa���% �g;{LU��2%Ɩu��)]օ�W�L6w1[҅K˟�Pi�n�tl���U�C(�!Ut(m�]�)�@����lWjME�	��F��%���RWٶ�8W:�WƸ`H��u.�z�;�G��t����nf�ķ-�F����-d�F��k�_��)S{��y]J2��qY��=>U7���*����q� ��*�y�:z��@w�XQ䂱���{�kgR�`q���!J��2���*pfO$F����oV���TM1���+���.uNx��]�7Cvd��G0�K:��8n���MY�;[�m�rl�9�_+O�Eqd4��䣣X��s��FA$Å%D��օ��2Y��G;�Ǎ��
}m��cM/�L��Hu*�R�N=��8����Cx��*�iы�ot$�0r��|���C��M��z�s�F��<�3���WQ����F [J$˧�:W��2i�/�m���x�u��GU�«MСV��Zd���h���`y��ox��ǐ�Z�khLW��[��9��-���v�nu�N�@ѥ�^C�L����f�boj�֪�[ci��.�Z@[��m-9�:�RW*��{��[y}+0��'����yԹF��os��fd�KBdR�Kj�:��ݸ�WVI-X�+����mӗ9�F7�ٻl'˩���hh��;|2f�~&�2+�w:JM����s��Y���m�b�[��<�ga��˖8�%$�f�Z�3w#�ֈr�F����㝅��b(󛱝�:kB��^$�J+)���b-���̌fӕǧW�Ă��9r�l6����h:}�k�a他���B_w������:���V�Iu*�]�Fm[���^^��k���V��_t��|60N�m���r������yF ���g�[\ ��;o�m��/����=�iv��@�#� �MZ �47��k�W���m�-@��t�kkvjFF������up3�Q��[�t�j�9��ke`f���˔�����u��.ZJCw29�j���K���S��y]�������
v����e31v`.-��k�;�q[�܏�V�Ǌ�.�7�ݑ��&�/k��dVuՌo�!1_n���e�]ܮ�p�S��l�C�Y;2A��>�DOhG%�ݓ8�Bn��qK�e�j��Tv-��ohu��u�%w��g���҅�n�o.|r����^<��L}b<����KC��Cӊ�s:��^g��
��_�[��v��aVc2����<��t���X��}�W�0� �Q�e�11T7�Z��K-�U��sj�{�,��duɢ9׼�j�]u�!���iWe ������B���x�+]���,�hj��T�0h��;J�-�+M�fV���|OT�D����@ȫ���P�w�+Y�XZ ���7Ǖ�t��[�����P[�*�8)�e��o`쥕�L��)�η��{|�8��&o\�+P�@�7-��(�)]��Ұ�6ug+��v��:Ζ�hԷ,���@�w�����d��1��1�Â�WRyJ啭7�8�����`�����TMm�k��m�j��𱭇�9��4�2��ir�\juݖGX�G[����n�o���-�z'B#y�6��w�mq�~=5l;ۄ"o�h'+]Z�Q�����΀qj�h;��ҹ�؟:ۦe�fe�1c-kZ{J&U����(,�P,}�^SR��='ouS����~B�����rFN��{�����ӯ\�we9x�>ޫ�ܾ�h���|�Y�W�Mq��I��KPݧ��4`�i�΍�͹0�Ն�f�ޫ$[T�˹Y�yM�j,��B�oZ���+6����v���5ݏ�&��rB��U���\�Cy/�&�}��\*��}b+�n�sYlom�Q� ��%��nTjQ������P)Y���$F,4�$��*�3:�qoV��b��x�[��m���PZ��ZK<�m�R즈���:�P���7�Ʊt�9����4q(v�Ջ��H�&i�Ը+�:��u�ub7���)@�DlT[c�C�I�@7�^�}Ӯ4�]K-�F����
n��M�ب+��m]�%mt��S�7��������Uކ��cz¬]�"ʱx�<��"<��VT�a�(!A-]i��"}�[�w
b)��a��U�%Z	��ic�w&i �W��&�G��{b�x3d����enuC"��J��UAm�&��fq�<��KpYb`�ʼ�gaɁJjL�<����b:���VVkb��v����)�]�[�PMp�B�2�Pd����I�f"����^]}5�m	��%��pH?j%d}ux�F�
%ˮ���p.�+r�DM�P]tҭ��!wW��D�
�C�ȳqHvzv\��X��#�٠�R�җT�,��j=uc1�6�v_��<7�r�3��f��z��36�.Pv�@�vN�/�№�L��Ɍ�t'AwK.����:��!�\�7�v#������
�^Ӗ{�nL��I�v�9S���ܥs���RlW��U7Gu#؆k�h��9u}}���*�V���k�HӶ,@��p�.���H�-|����b�v����ς���RN����M�Yk�j��{Ő�K#�}ڸo��X�E٩/w�S�AʶҫȻ�D6X#Z��l釬nKλ������xD�Ǧ����W^�0!y�ݯr����l��a4���2�5�2�l��d�U����eoo,"�Ub�\m��tEe	��T�25���6	Pj���mh=���Ğd��K�]B���;~s cr,���yي� 9Ie\{�>���Gթ����T������9�%w���J��]�Ơa��J�ޤ��R���=uoz]�x�<���K�`'9[����E��{U�4B#䲆�L��y�+("��W��Ku�}C��3w����+��S����.� ���H�W�EK�9=�:�;�rk{����<%+'lM�t���#b��G��gs4{,��R�N_(�u�*�_f�ǝ:�S���̡t5Te���5�]��QAܦ-����j����p�E�D��<3�lj��A�)�mGy�z�����#���w�e�lq����%\s{6�:��W �|2eA;�4�f�1�X�3J�8�(?�(����3�u�+hv�u��Uŏq����˒ J�tehC� -��X�6�Ѩ9c�t�)�S��J˛�׆����D0F@y{ө�/jI�;$�6ڼu�e�j�R���e^�g&�.{��9�XU�|Յ؋��|�<�I)Z㧍��bv0̜P>��m�[�ݗ�-!^đhL�*�T]1Q51��^��&�q�g3�	Y�۵��5Ee��擘uE�������;�u:����{���A��S�m㣣�Q��*�u�d���>�U�P����Co"Ʃ-5��B/,E,�ǵ2W/�l5���%�Ά��V��+�e���^�������p�$	'�`������Ca �@��H ~@�B��'�I ��vH,�!X��$�1CBI!(��c �� ���2BHw,	=�,��BV0 s�$�hBViB�� �H-�@� I+�!�Y n�$�VBgl����XC�G, ,���&$(�=��}��,$,�� |��{I�`d9�st�@4�T���@RH��e,RB�I�M�*, �C�s���>�c��o���`(C�ή`�)��1���VH��h�'XaĞ� q�/(�!��
@�i<��4��#���ܰ&0 ��@�'���M��|�	����ɘPP�ICZ�O$�$��7�3�L`m T�d��L2,�d��$YP�1 ��<�	�JȱI T��:�g�	����d��&!kb��tHqhCZ�7l�J�i����;��,�`��Q$<¤�]�6�
�9dQv�0�{�����C|�ڦ�Y$�d�`�����)�.������(����'�CI��5����B��`kVM!֌����e�r��}��(ECl*G�S*lB���.RbIY�AAf��YXm
������"@������P���:��Q]P�&'�r��hdP��g.���Qa�uC�kVm&٦��P���Ir�!3VB�
�d��q�Rc8�3�0$�}a7��>�=�u&١�q&�PPOY��"�vq��*�'̆v�
���yIX^���v�٘����d>C2��p�s7y�3��0�XT�׈72&��.��8��N4H���� p�2:��ַ�}lb��H|�M�����F�Ɍ�J�ut���L.��/xa�4�d��:[-����M�o!�
VAuZJ�^ٴ41(Vy���A���#��!��yC֗��t3��̣iP�c1�߯�k���0�N30����2]Ӿ�SM8��/�����S>J�h�`�%ՅE��t�^P�7��hE����%�-�iW��w�z�t�fDw֙��{�4(i����wk�y��ScR&{$����y�CGd�i����l\�GW�dq6�<��Hu�޳�s�먌������)�U�^�&��]�f�a��,��wY�Yǿv���lC��*���_nÌ�~�IG�;aR��;ۦs�\��^5u�vj�>�Y�iP�[L�S"`��ںAR�D[ZL�C$�d@S!�B�{h*z�of;j��)P�[�Fi���]��,m���I��G�4���\�@ u��/W΀�h�h[��\JԄ�@D�G�K��l*6'�(A ����VEKk�+�JTf��
R����iJ,�Bӹ��q�8����6�� � �m�E��I�Z��|+�ΥH�l�{/��TpG%�T�N�Ѥ1b�Ѕ�P�E;��\ͳ�������@�3mԫg$l�V�I|~ýڀ�:a&��&a��e�K����ű";�al"S�b�QA�$�T9e� H�ˑ���tǖe�f�H�T�0-Y�&�[ѡ�(|P�L�������%d���=4���x�y5S�X"����3i�uT�!��X�!�$�u
�ֹ,{��s^�o�g�V[��n��k0m:���d�ni���������`�"�i��e��mG8�鰈�*�IT��HcC�z��y��3���G��ڕ���(.��� �'k��)�uۭ{]�'�;�j���"��Щ �8L�� z����B�ĥ(�ز����"���dY�Ƹ"cO۶�h����@��IT�� ������ʹҩ|$�
�ExK��j�R��QݑSV�g���8�xK}�v�
�h��l���
��W|Ri��{��xU6¥	
��ي��X�g������N>���8Y.�h��1	,��ZT�jv)G�A��o��)��PX��Dڧ�3
�%[�K?�-<z�����R6,��jc^?�h�L�,aI���F� `G�~6��ɖ�!��^\x�h����x��L�����M�ꅒ�A�&���]�6�c8��@1�+�&���t����O�p�)?$�D���XLB�hp}Zc_}J���SD|�ƣ	gZf���H6i����*�(x��Q�Ul�1���H՜uM�	��+�(��!�k@��㛟$�����/�R\駦��n|��<s�ᵖ��{&�nwZ�>Y���v,���뫀���,4�EjVi�DL��n����*6�I���m)T��iA�e�Cij�W�{Lx���sK�5�{3�(���d�Q��,,|8AV=;[�-�"�NPT^��e��!\�H�	�o�73�K���ү3��T"�-��K��e�W�`qڣz�!4�qRciY�@²���XU�~ ���6�4uS?����. å-b�������ܫE�-1G�>��r,b�N#�j�)v�A�~"4(E����9<�B���8��]��:M%7����[b�0/k�U�%�D!"d�^4ڽˡ�3)��B�4A�'�6�{t`�^H������C"D1��JE�W�3B�J&�q��^���--b���f6DjJz,��$M�˲@���Ⱥ6p�
ΰ[ա��e�j���)��i�!~D�t&�x(QT��ڤ�T�F�M�0�b���A��e�r��p/�<���!!/�me���7�2������C�&e�7j��(jwc,ҧ�6����0��8��5u.��7�7C�^�.yWcB�QB
��Jyp7P�^�V�W��E�ҕ:�좳�E�
եU�� �l���N!��~_�J����f�?X���6��B�4F�ʙ���0�Cl���`��mVş����G�7�hDF�uz��	�_�r�"��Ɛ��уF�̆퀨,�i��-�H1T�.��Q`M3�
C,L4 �"��P�����W�f�6쀨���f~��c	Q�@YTѶ,
�R����1�`bZ8(���f���: ����%D�qFv�`�0YL��f�����F(�L�8@�j��wND!�#C.m�Ć�UU��".�I��D;�η?,�(�9/r�_�����;�%A١�f���ۻk6+*JsJ;�t�Րf7pZ�N<bmJx���y ���������?�����[��!�M&�(�	 ��	�$S��d)�-:Q�eU7�)�A/�K���������wχ��	�IW�MK�:�u� ���T2l��׃�?��8t52���\��vm�C�v�gvB 牍�z{��A:�n��k�_K�Ґ�r��*(�8��P��s�"�Vj�uRQk�H���Y���=�>�m�C�۽7{9Yui_>r�Ps�E݅�5}}�_r͢�;u"��x��cx2VS����c�g�#hb����LA*ƸF�+��w]fm�c3P f�2�ε(���ږ����T�4)|�qQ��7lm$��
[��li�y���P�~�T.]���v�v]��Xwh�ZEq���4�������WjdH|��(�g�@�������():ރ5�n�-�����a&.��bժ���٢��P�	�J��K}NNzV��v�F�xo�іm9�vl��a|o&S���q�7y9�,Q�-�<t�9k�vu�������76�M�2c�}���d�J�^3c��GCc<�z�|ܲ�����jU�)g.w����J�.9;֖û�#�+��f�B���-�RMt��4l�=#Wm-j�J!�R�wuڲ+�m�j��M�G5%��֍X<li����ۤ3[�eوұ�=Z­\���K역�EG��xk�Ft����uN���H��� ]������M�E�T�u��P�wH�-�y�����������/{�t�\/��Q�T�>ItM��������������=w��ٿ�I$!�w���y[�j�n$�}��wRk����)��i�ʘ��9b)�z1�Yc�*'���G;Dǲ�\JӮ��ٍ�Bs�����Xx�媾�Oh�v�u;���dy�G�Rg��\~�uo)~�}���m��`$$�	��Bd�8���4�	����IXC��:���C�&�r�I��L�� y�I�(C�}� �5���I�!�Bo�ΰ$�$4�/y�e�>�r�3|�7��|���((
#X�EV"����*"(�"*�QNRċ�EU��R*�Q�)�NZ* ���U�*ł:j��"�(���B�����(�2*�����" �*�JEX�(���q�X��>IX���5���UX�1��Eb��U"�F*��5�eTX<K"�*wW_�T���F+RR(�UV`����B�B",X�|}�Q���1EDb�PU�����QV
�EY��wgE
`*��*��5��X�Ȉ��Q��b%�U"�� "*���*1bŞ�"��D��V���Ȼ���Τ�UPX��UdEQ)Ub�" �Ȋ��F"�D���b�1QV���`�	#R �)ňԶϱA�ó����j����EQb�#��Eb�b"��T`��TEEX�((��X��d4�,�j���4�b�
�+4�Qb��ҢDT���c�PAUE*�"�AS-���V1v�QTb��U��U1��X"��Т��*�fb���,UX"��X.5���(+l��rՂ�* �1~j�PcUQQX�Ec�S��0*("�b��b��UF&4H�iTUYU���TF)�C���ۢ"�b�O�@�*�"��T
����}���~�m��ǵ�j��_�TX��AQ"�D@T�b핋��ִ�PU�"
~h�X,Q@D�ϵ�����A`�`�TX� �β������{1Gv�"��;h�ő�X(���+7�kJ1�"���1W�H�
����Z"��-aO�FQ��M�(���w��ȢŊ"�Yb"��(1wB�*�IDPX��V
���E1�m`�������uR�UVk���"��%�j�E�U"(�\����m�#��zw�}T�hH ��$�YQh���X�E�f��PQE�*bTQb1��փ��#�*�PX(��w�ߵ�c(������U��z��`�}B�~Jr��g�A������b��3�qE��Eq�ʪ* ��kF�X��"�ER}��}�
�TE9N+1����g�UU8�PY+7�����=��og:����&*��R�E`��Ϯ�hTb���+��ib���X/�#����Db1���H�v/�EEEG��1Q<�pX�Q>�fZ*��;���b�1^�$o0�UkQ�EQ>����'�(�����UG�E��DF*��Ua��}�����������o�y�`1�W�E�ܬX"�1ue�ߛǬȊ���z�B�����:���e((���
��)��'m2�>��mq(�)��^��a�X���^~�#]�Ub��)S����b�E��Q�U�������]����i�����OͩWMU��������V
�U�LEDX*���V(z�UP5E5��[MZ*�1N�Y�D�UE	��fGv�����q,u�y�>����P�F0D����DDY�ّAk)��"��k>���~��.#�Yu�䵓7q-��X 
�q Wd���}�mQD8�*��Toy�LQDD8s�K��U���&w��4��0l�JŜk�_�+�M��*�j�TX�$���,YR������9��#���N��.��ו��t�o;/=��DE���4�*����~J�U_W�f�*�g���R�b�=�1TH��,���i�.4A������.�{J!�5����V�b��AW��8^� 8ѡ�ڦ����:b@��=w�Q���أ3�:ۼ0ƌ�k��t�b7���Hj�Z0uJ�r�o��t��>��H���N��n\�o����:���%�g�V����V�ku�J����A�!IT���4��C�*q��^�LD\J"�*���DUWԫDݨ���kzUk

.��{F�UYYE:�Y?}�_����#;h�~h�����TcR�b�m�'��كU�޻���s�o3��c���Yğ01P~�hb�dO����رE�������|�R�/���z3tEO֌̢�S_�ڸ��(�*��>pWV�o��W��~�E�b=�1�TA=��B���v���N��3����k&o���aD�H,�H�o�,妋b,M\��&�j�(�[*���%g����3[���^YF*~g<�\,X����R���(y3*�Ǘ��M�1E���ֿ�Y����?Y+�w.[���	�������ד߭��6��u9ۤU|՚j�k'�:��N��4~��X�����K�Qe����O�9t9��T�U^&��*�����)�s{��0D�g��)~ �ɭN��^^�(a���g��C�/9솘�l��s��/�n���&�M{1yjs���]��UEQR��2~v�)T�o�_��PDO��;T�1^2��U�3�M"��Z���QG�L���%�{�##��š��B�|j��
,n�t�1~k�DO������kGp�2��=w��k�}:�mQ2[[*�"��_��]�T�:�~֏5q�Ɉ�?Ͱ�P ��E{Vz}C�pɘ-�^��pÙI\U�̯�4�$$Q�v���ډSg�y��^\U`�Okxy=���4�=lF&wδ�;j"�AU��?4]'r�~�3�Z�1-��3v�頧�ʁ�A��6�E�F��w�B�� O�H�g�i"��*���c�Љ���Y�Ɋ/�Q���S�b��/�77aX������k�P�f�UQ|f�f��S�E�����F�*,~k�(�v� ��[�[�[޺�y�\澴�<�'m���F���(�Ҷ�TS9��粈��ȶ���1F#"�5ݽ�m\��jUb��X��H`��������o�ԏ��H$�!K�Pބ��VW��͟k����wpbn�O}�>lY�T؞�4v���X����7�-�S�D4�������h,F(���S!mQ�-��*�QW�v�b�~���E޿wp�U�J V�z��`!1Q���UڔQ����LP�:�޷<�q��bΗ�8�ցt�Ak��-f`9�h�
�t�]r���s�T����usyu��Ĩ�9+PQ��i����� ΃Fs�5�r��p����(�F��U:{?s�c�3�k6��lQ=B�-�Tq���c��md��j��N�DƊ�;_}����V/Ţ��LG���ߞ��T�"�j��dϽ�*��jŪ��{f��5:V����?g��?r��k*��b%�(�����~�b�@��� �N���e��Y�U�J���Mcbq�[^���sj&��T.���7J	�Q�RA�Y��F�G��W
`�?�^�XH@�vį��O�
n1	'�V�����$���#�,��I��G���F')�����Ek�~��+1<��u���x`ǉT�wc�ϳ�Om�f�,���EV�p��;�0gT�T��n��g�҉�?d:���0g�QDY�S��l��<~-� ����q�b�(|��h �z������N�
Ǩ�w��<ӎ��~>�C��mDA��}�1X��u�Y�\�����!q*Fw���01�K�3�Y~���6���SM��?%�*'{��vmP�I$���<}�=�/<���'���~�8q���7��uD1���/��u~�u��\�q*4�<�%o�^�{�b������ٰ�*1a�)��Mޤ��L�ʿ�aF"�C��>��B�G�4��C"�|D�7ퟹbE����{���,Y��'�\_�\i��?}� ��,0��!SL5ҝLG/��8)�����j˕�}�H?QO�����7�67��"��ʊ|Z�~�|�|�F*}��Xjӹ�b�n�F������UMZ線����`)���~'f����'+&�X�|�uk+�W��>g�#�E��}|n�=l?w�����\�)����SY֋��K��A���Y�h}����u����#UUV��f:��u����~��۷��sPhx���m��.jZ#�i�����U��<}��Q��Ww�
�O�QM���r�?s1�5�S�S�*��S��fj�#�Ǽ|AD����os���O�T�dDg��k==�0��5�ԤD�#=��>ȗhbS/3���gfP5w<¯G����+�6U+A�ˢ�O8n �LN��G-�xNMc���1�'`��8F��5�����r��WA��C;R<2~Z~C�f��ǽ"F�0�Tb�YCm�Ǽ��B���������Q�����o{�(;o�OwYV�𿙴�lM� �H��׳W�)�?g�s����bq[�o�(���j�����B���}��w��lٴ��]�3��hT��hֵ�0�������I�G����#Ԝ�ϟ�L�lV|ۋ��D5�B��7���,���4���tv��D���CIK����6V��?0�ｚ�X����oB�m���QtkZl�Ym*H'�~�z�L딚>>��m��Lxx�u�wY�S�a����qSM�|{{��(�j�Xe�=[1~y�f���^qX�x�?;������欱��V���}W�ڋ��	FJ;ϔ���E��-!����p����_����ѥQݝ��}��[�&'�X$M�$Ro_��l��P;��i�J��,�&8�=�yﾯɷ�^t��Y�< f��o�����Tk�]�]��i�~�;��N!����ѤQ���SE�Q������;�g�~O�C��f�~D��M�k���T��Q���Bԃ�$����1����θ����I�>�b���WO�H�����I'�yjE�l�|6n=���X��,�	��0)���W�#���-P�D�Oٵ�F%��#��8��c䨠�_f)���}��6�CL�s1���U~Mbq{{�T7�99�8��U+g�?���3Y�&�P$�Ce���E�iB{�O��t�D�w�l����C�9`�,�\jD�m��?�B�5o�k{�+Vo�ob����`���g�����(Q&�?a9-5�S�u��.��Gɼn�xր�5H��t�X��+��Ԫq��_kb��=�����Q��P;��n�}�yf�m�]̙O��o��ذ��i��,��m���:8VO��]�jU��D���M\����݁t���N�[29C*�٠�akIϦ��j��P,��8Y7�:���rb2�79i�h� η+���\z�J���oP�0v�[�fNч���jC�`���ʀ3N�'u펬��QM`)D�&��D:��CR A�οw�S�E�[�q�&�ݞ��^S�Yם��w�kߩ�WT���L''6>�R_m��n��/;�+����n���4Ti�%	!}�ƣ���!0�2�_���.����@�>��++���
������;�"�w}E����Qw���	m������k-3��6;��Ur��j��f��d�h
6D
Q�؏B��_�V���*wGRv�+;P#�Z4(
˯��P+�e��0}�"��Nꆁa� 
�xW�F�U��O�@W�&B�|�8���S�b$2}��
G�sA>b	o� ����f�����/������C�{�~���3Nf6��4��$ij	���O��P�b�7;z�=l߯FЛ�#�� �n����i �䆤��M�QA(*�D~D��TFD&��u�}k6����1���M����$8p���g�!�;Vuq�e�}� 6�L_�c��}j1���6m1��J�҆�N�ȏ���ã|mo{XR����kǼ�{,����Z_� �,���=魱��� ����ضuL$ef�͂`���92"h̏��]���#XwT$��jL�\�"t�����#��EC����m�Eo,��0�����VyC[ 2 �@�'m�4T��"Ȣ�,
��.i��vI&�[�ʿe��_�|��֦�ֿ��0Y!f�Hm�*��c=�Wm Ï8,�ڵ2i��
~'_H�U���-۽��s��Y���s��ĒC������\�'�!	��� �� �2m �II �C����>a�@��'e�]�� ,���R@7iM�`u
!� q��@��5��y	* y�M�����|��HJ�bN0�:��|���Cﬀ� '�\��]g�ֿo���>�Əs���s`��'�d�g������s�LT�E��f�+�`鸅�s��2��&�iց�@��= Y�"ȨΏ~�tsp�5�*WG}�Gug�g:���n�	5��|�\��n现ך��`觺=&�"�M���ǐˇ�����F=��eNP��3��9���z����@�����~ �6���^���zק�ݒ�{�x���e���@�5�^ΕcƢ1�8(��a�ă}̔���˱�w��||�O����LR�<F���W�׾J��*��,N���R`D)8`��� �s�ҭ�Cw>j�R�~�?P�Ο��y���؋�+;|R�>f��e?4�z�}t~ S�}u;�:��{O�k�;�Ӻ�"u��i��W^�@0���H��$�����=T}tO�&����T�"U�;`���(�~ ��>�iJk�$-���CD�yχ@��V��U��U��*��H���0I�c�(�1H{n/{V�~���zQy r�P�~Y*��\)�!�B��DU���}A���j����n����.��?�ap��Q�ʗHw[��jد�G�81l%HL[i}���:1��p
^���_4@�����p�л7MЖ�S��n��B4��dyu!J�b|��@��l���7�b�|�*e!����1��ѡ��
��T�{;=nX �" M_��ڵx|��B�@��w��Cey h#�	Re��|�1)�~�,��- g�%E�i���"�pNj��iF����+����?���꺍�)�~���>|��I�Y�Y�$�!?1O�$6� s��1���΢�׺�B:~��9�׾�ٳlc�� ,m�$�E ���o�����w�7��^�$�%�{QLa}q���OfY7������{Իo��x���d�)�^�-~��-[�� 6u+5�Օ�G[i0&dv�i�rU�8'�~��y�nR����٢���(��6	?^��D�W�F�E>��(|qI�ڜ��������[�G�+Vց���J��׮J�H��dZ��CyLaY�}H��D�ď�!Dh�B���7�hP���A�Az��>�!�}����*b�0۱[��@�B�o�*�|���|w}��j�<"��ث�Bά�e�x����V���	L����cI]��z�4��I����R�TABB�=#�� �s�{��MW���7�@��̫�t���y#��4o�@���a�
N�d��7��0���͖��ƌ�����S�q3Cؖدg+S������^��ܪƱ^)�^3���ɻ�����&�.��)B^��}���	S�MN໬ʲ����b}c�**���+Z��6������>�����#��Z���:(�U�y��B�p.�S{�w��`uz���A�b1�'O��6!!��cW����Q����WKEY�i������<ʒa��&���4n��
LF�U��'�e}.�ڧw���B���L���c��+��Z;|W�՗��ޛ�QC�Ι���/*�ܯD�hD� 
 j��:BZ�$�R�K�G��~���_�za����޻/�~,T�W�+֣|�\I��K�\����\�Z��Ԡ,��v���ə�������M�P��D���m�q�{�U� +)�M����k��:5(MhBƞ��&�j��o�΋��$K�e��Sf�v���v�G|�lZ��B�,1)x��� ��Ɉ�HW���BAk��Yj�0O���BG9t�-�W����e旎\��B�1[�F_�2��a3yYR �"aXZ�+�d�X�#�f�ަí^��}�^�eE�Y	�f����T��J�_�:��s44=x�t��閾�R���&֨�P)e���Z�u ��M��.�n�{��s�oX�EY�sr�Jbw$4��ʔ!����C�"��,��-�
�.����#�Rt#iy��$J��芨n�����,x�`��P�^j�7n�/}>u��?��Qv�]�ˬX�>qBn�޺�[KEo����}����{�LK�!N�o]1b�����|�w�e�o�3�C���2Lf1��WR'`��A�NC�[\|�+D�3Q��o�q��R����Ϭ}l}U50s�i��61K8�b�8�z�{��o]k���k�+�@���6��Xw�y��'Z��'Y�=��w���:Y��L}�B���\���Q��R�Z�*��<�Vy\%`̣0�^w�P��{��PP�l��� V�]ФQR�d+��RĈ���,�ڤϽ+��2�k@�e�C��F��]���f5YGԇ2�B`܎��f�j�I��*m�.�S�j�V�֊3d��\j��.֋z`q�TNKW{X�������%��T�`����^��Y5��^1�d��ZM�Z�4ΜW)�F�AP��է0p����j�Y�$F~V�캔�2JUki%���p[@ä�����:�˴��� �>f�� �(H���)1M�
�i�S��-P�b���Mu�I�N��=H��=���d��/B]{<��T��$��`RP4�\ĝ��Ru�qAD����,�D��D�V�%�iԶ���qӬb��g<��N�@`v(�5̏��U?�1�=B䴆t=�2|+օ�4Ʀ���d�!<���Z1q�^\�Ƀ���/�ₓbδN��`~"��'2��YJH;>��x��ǆ�?[{^���7����WV��b�:�BxY�������U����;��k����g�ͧ��U]ׁ�N�8=�=��;�{���@K����R+�49�z����(��7lS��1v���z�x�Q~<AШq%��h���W���wʼ��(}��R6ZU�x=s��oV>�� ��^�AU���1֎/|�g�u�*�����1ゝq�A����ߗ�׹T�4�WE�����k"�i0�~c��\�x��W
�m�5�m�UT�w�8� n�Ӂ-�~ۊ�^CD�m�0�Xj�
&��S�-�o���%B��3�U�N�E����P0M,nW�܉���^��xz���j��O58���j�ZDU԰=CU��ō�+�j��6r㾜6to� �+��pit��w���3^H9ҳK
�^�.� �"��EP��3%yպ��e���t�� ��Y	�6�T�Ty���g��U�BWq�{y�w�����?Rx(  �h�9�05�`�1��x+^�G!f'��)J��_��=���`����2~>���b�a�%g@�"=�r�&��Tk�]��l)�˯@-$�q�*[���m
Έ ��> D|���5>��>{!�p�_?zr�@JU�wcuVk��;�b���D�y���h	| �۟�؝VN�B��o��}��.��.�^򎜻�O:!�1�p��U�uy/}�5�i��
ع�	�̿0��)����d���'벀`�NU#�S �C2�(�l؂2�4��<�� �wo&cc�Zߞ}�C�>���NF����_��axך��B����Q�Ҁu]vޞ1�sh��)�]\����c$M0��45 hi�����Ӗ�8:��\��n�S덛�}��D��jڔ���_N7�e�g�B�y�C����UH@�[��6����T�5�[(_��hB��fx�M;!�@��϶`�(p��>�x�݅�MR�u!zߔ]偲������<���>������dx	Ɓ�yƑc�> ��v�e� �^��[V��X��ܱt���#�xy����}��d�\�@�݇oH�5�	��ӭ�G����Q+��
��ob�)θ@��,��F�%���ƅ�3^����`�p*#e�M�j,����e��!��૫�)	���˫V�=w}ٺ*]vt�H
Qb����w+)4.�g=z,-p-�q�Qž�λ�1��gu6wW�&QD��{;��7��ܼF�-��7����]�j\\��p��z���b�눢��fv;�m�Y�-�\�L�����zxq���ý}�����0�����0�������G��s�U5�@Պ�怂��;��*�it��ѿ��u���z�[O�۩K�79�i\\z�m�^��2E&��]�*V&/��S9��kif@�����a�T�4�;VrE���X�qYS���8_:����_U�x��]�%��R�lK�)s���7+R|�Ρ 9�)/�N�z,�tBV��.�8V�ܫ{x�*�7�\��i�}h��$C��v��Q�Wz�]z�<�][�7V��zEIr���c��wW��M�U�[�� Xyj�����	ǡ�Ҹ.uث5L�5�5���j]+��U	1p�S8�wY�Ճ���ͺU�v7�eh[��j��3���jw˓�����SPуa��`����X�>۴�:Uɲq,��W���᫫)D˭�F�y3Ь���|*V"�wvK�RS�n[��N�DY7�EU���TڇuZs������0$�Bʢe��/r�ޚ�nq���ȳ��+5����ʾ��!��[,Y���o�7x�Сaor�Jv��g]t������WN7��)k_>�]wٵ���z���!`���=Ȍ꼾��(�ը�Y�1�{[��Lw��-2����I��ɹv��-��K�BΫņ�l#r�o�ޣW��2�3]"������x����4���M�V�=IQ�:����ܳ���4(k�o�V�<����s6.��i*
KQ�zz���;1�r`��D��[Y�	vΣ
��Ns�8T�B3��-�v��[�/�v������(9+�wں�ƧU�5`��E>jR��D1a�;k���3�s����@�岖�Ǿ�����q��Q�;��F0�$���-)��l����b��t��f��7W 0��|�����ݾ����4�\����/���{������;:r̸"����R���F�K"j��L �R糛� ���r�C���+l�9$n�Ӈ�����l�{$���2����.>���!�QP/�'�Mk`EyƮE3.����0��P�מ�߭H���6�+�ŕ�r���O�����8���c�_f��	���QV�X���z;YOEWd?�)�"6�7��G}�?*�җvhc0�>(��rTIZ/�� 9m�p�p}jrB:���,�y�������6a �W�d|bg.�GQrͭU�c~�J�
���Ml�c�?w�H�Yr5�+�8�dh"�dm,���&����)��S�e�� l.�j^��>���KŹ��Q���T�Y�Rk�xS�����}N����Hg[y�Hȗ&
:P,��
ʡFL�6h�
����R�M�^DGZ�N��s��u�b��C�-\�W��V	��2�!L7FaV�hY��V;(Ҹ)!�GN�:�����i`�9�3kB�^��HN�����&�!H.��skZa�w�_��X_�J�ߩ������i�C�A!�Iy�t���E�Eű	4'}�r+��׈���YV	�T[��v�Ij5J��>���G�\����WG�2/�P	W�s�޸b�.v����ۧ�p��kM\��<��pkI��*�
|;���ՙ	�vcu��!��'�"�"s����O?�q��c �$�ւ
ޭ7ua��|�65b@W��U�+S{k�.�mJ̗��&��7��VF.�nrP���|�K���U�KF��霊ع=YH��oG����o�^���u2�SxBK�����7�+���e?T�3܏�+�6�=��"n$��**l�n���}��t`��y�@���@��C6N�R�)�h��^n�:- �۫. ���4����#��o�>�H�ccU���Ż���z�����d֛�и�����Tm����w��?O�=&%��T���r���)^Rf�f�:y�U��Mr��Z�#��͔Q7�/I�/�s�"x�^ȶU��a��� KO�P���F]��XF��&�vE\����E(��jW1\ZQr+�Z�.'�0��o�R�LV�C���n�"��zs{Fq�9��yEp��z�x<�z}��D��{{��ZGe4~�1��xis�V��遗�b��G�΄̭�� �:z��C�jv��tFK���;>8h���~��༺ү���[�ÜК��I��7�]8Yc�eo�̮;�ʼ�O`��]��,&*ϵ����Z�1�ϵg
��ٙS<4��[R}��e7��J�G&�ϧ!�U��Ͼ���}�Cw���~y�}�І��Grݱ��0�HH똁d���ky����f�"� 3C��1Τ MYWnL�b��_yw�s�n�øRq0Cl�4c��u4E�3iVxWNQ�<5ӯ������o���@��	u���bw �M�^���>������eŦRSӪ�v����}�c���u9������ग़��&Of��{r�,aqj�E�=y��QaLΙ�T�jN�Mch��kH�F�.��-V�"U>`Q��6�p"T�[��P;��v�ѓ�GM��z�gp�u��+q@�����K.� ��򿿫C�u}�'�/������ZE�W9]s8�a�O�,���?)�ڇ�7�JVH1^�R���Fw2w2 ;����a��޸X1.<�	�Zl�c�VI�\�}l���I�5�����9F?}��h3�����5���+��4u˟�?n�ߒ�����ACX��#R�2��y�ׇ^CI��O�����D��_<�@�y��e�C}ʒ��)��@��^`D��[�Y(�	�����k���/�i�L!8��v*�v�V�<�>��S�vO��b��<�y� �(1�	�L4Dc}!>R�:h$i*(Ru^�i23�u�uK����fu�]���SL�S��ꦵj8r����+:��@���i�/|D�;Z�P:7L�{�h�}�B_��0��%y�]u}�ޥ�e��X�ԫ���W���a�G��z*�4*�����{��vBo�� ��ƣ�ruc�;�´]C#R�	n���J.�zꗟ��N/n/d�c���KAg�W>���j���uc��t���4�������_���~:	�6ĕ�2*ൕ�?�{�}TE?�r������q���v[�!��H�*%��N��ކ}�2/�2-�����9���>���cf/��&1��O�6��Y�l@bc�(9�C;2(N�Ged���j\/%^m��t�������wƑA/���-��A�������{�AGsZaۼ-�N:[��dhu�[Ke����1��3�b���GCEu�Q�y���M�;;�
Ծ6&Q��n��gZ������j�	�GuRW.]�ٝj�S���N^�ܡ�{N�81D7���ݨ`s �T������R�����u�H�}���4�)؎�^��+V[i�׻�'�����sJ=~o.�1����� ,�_ݛ,8v�]���-��iߦ&�їX�݉>S�y����]�1;ն��u����e�1��mN�Z��~թ� 3{�݇c }B{��������fP4s��� D#�}B���J���Wׁn�F��>�CH�06��nP�6Ɍ!�{�	�P��3��By	�b���8�w����1��ì&ϨoT&���HC_�	wd�	�8��`md�`^P��5̀~I� ���	^�w�_�S��]
z�< ��&�CO�1ߵ��
B��>��P�C	y��n����7C��,��E	�?`�Hi$��00���B?��f�q	�L<��EK�
� x{U�>{2=�y�:"ieV(��HU`T:�m��!�$����uۨP���C�,'Y�uaPP��q'��"��?g�h>`i��PP���b�P:��A@�>��P��4���/�ﬁ��@������q��Qo�M㬻Ϟ�S$��{��0�8� ��2C���� V�0���4��L'�~�l!�����1�gX�q�A`}��P<�������<�y�	��C�
��a���@$}G�<I TQ�}���
z�s����C�!P�'��3��~���d<�tOcN]�,��U'��}v;I���(��*��t����q�
�g��!���.�v��;�X������|�B��fdA���\�#���>�G񹏁���=c�ɻW�#V�^ ���(�{��hm�V	/��I�L�d.���s�����̤���l
�r����L�
��!AT��w�g�J��K��^g���W�-`|�Ŗ�D���[ڏ�v1q��O�Ei]�]a��&��$r� ����k5ƅG͡I5��\؅��^���6�����y{Iq���x��˂9Z/�֨�ʚ/����l5W�q�����N�̭ܺƣ:��g�*�~Rf��CƼ��^�9Y��ʮܲ��r�����u�^]������t�F�.�P��h<��ѫ���/.���s�ϦS5�ks�ך6#b�2H�1:3�D&�G��{����ꊷF��rT���m �c���CH��w����W������?%����\���oL����y*�_���З��u�n��sba�[}-��{�fK�P�7:(��h/�e���������<q.�M�{�-�Rlf	X��F�Q#�}�͇��+�6}<������6e�U� �>m~S��Nٸױ����u�5���O����}w��*޶����2L��s�z�T�]�B�>�5��z��=�b���p�̸eO7M1�ߐw͍��vu4&�4�\��zu���#�j!>믷S����
���'�ϛ�MF�˸�13��L����V�QR�H	��V	ı�܎/t���0F�b������Ι0�����vd�����@�ni����m���'��y�ؽ��o�!҂���1����9~wG��0鿣����٪��##+k&؁��X�+�`���w��b�+����aYҘ��}�Y�*Ը�թ�b�/�_P&e}���E��]~�gR��N����:2��Q>G��+�-e��	f�P޼]ӯ�e�����>�ә���Vw6C��l����C�ݜTʮ�X���Y�Yg5�	��W��t����5�uv��}]gw��y�K�AT}]�:��;�/��rWa�5eݮFet�ߎF���R��Y��Dl׽��X��,!A��N�� ;�N��D�d�/�=���r�T�V�8	�7*�V���������
]��z.R�'� wT���$kػڽ��
�4&b⹭��yw+M��q���6�?e6\�J�Ńj E�yLT���ݸ�M�����c����z�pJ(VA�;=S�u��ճ�5�2=	oxw�'5��75V{���i��.��(����=Y{�)!K���'�D\H�ޣEk�����:�~��6������K_{%��Yl��A<��],и{�Y�?K�ܥ%�=���g爷�������̽ʅM���{Z}'�U�+
T�Ġ�m[5Y���O��>��1��]y������b�7z�z��5��~v0O旿q����*��v��]�٤Gz��+�A�d���Ǯ�0s�z��U"6W���&��ܮcU�x��WA�a��<;��@'Z�����$�����g�j>]q�W@?z��/<9E��7�=�[j�y���3�~�tqB�ql���Y�+��:E��(��@��͠.�"8d�ߏ�Uf��k��M��C�%S�ktvzW���'s������Ѥ�c���}�i�%�˃�N�/6�����c-���~[LU�L)�D��J�g��{�n_�HH���x�s4!�ۥ�&�Ps/zQZD����$�
�.�����.��dY��n�� -�\˧B������� f�<c��J� 5wϻ�j���7�ɞ�｛��ڼ��z��r@�lӔ�m����f/���U�~��q���ϊ��/�},�d2\�ѷ"#��oej��1b�[NG�yѾ4w���q�Fm���W�HH�7�$�g��Z}D\�[To�N�t1,��*N{nj6�~��p;#���kM�f��b�;���7f�QT�A��f_\�����\�Ƽ*���5����4��ߡN��|�ñ�cT��e~>�M��]J}*�z�/Sm��K�RH���
����s�y5O
���F��c|��64ZC�ճО��s���䫟d�~eo��0�xՆ�F�Q��ۘ:[��Υ�?p�V��Aؑ��� �Ũ7k,�T3�ۻBk���H�	�jw�;��L�q"�Z̫-{3gf�D�4Dug]ݐX�&���}7ޯ�n����\HחJ�J���${=��ۋ���\K�}9n���%�:z���kpN�N�B�ًƘR�j�f:`=�oso�!V� xb��*��B�����W�����[[�����2�q#���US0`��{`S�AR����_��`���4n������ �}�V����1~i�8��V����ԥ��(�%��yKz�!�1\&Ks+0��O�����+�>+_�'C�%L��������x���sD^���4��}��n�m��o��$���/"�����m'�:�R���ٝ/M�$-�]Lۏk�Xח�#��"Yw��G���������5�]�U�f�N*����XݾV���k��r����,����;h�(,�t�X�3@��n�.�h�g)�-��3��;5�S�ݝ����G�SR�ײrK���+�u�|4"�v�;wB�Ȗ;����DV�g��	?r�%Y��vXN��1�{�U��>Q4$Z���Ͻ�p�:�W���j�-"Q i�5�(W�nn	ƓB�+5!�W�����E1�	�8����MD��za�zY�L��9B}�Zj�n��)�2{�]��#y~�3U(NO1W���!�M��c���Q�ՑJ��>���+:�ծ���bttA����-?M����RnW�P�7&���{��ۢ�"�:%�.�����g�V}���`k�֫:�ѣ6H��Uګ�,����Q��*<$����&��uݞ���&ľp-�&��v���W�	2(�#J\_AR�^Q�7M���`o�W~�h~�Ɏ䟪']A��F�Z8J����+a�;����V�x���~Ϋ�)�tU�
ǡrW�3k�oՏ��#��=�[�u�l��ѓak�p�<�S/������~L�C�a����H,��(è�Ⱦ��� vX:���^�R]ED�_8�h#�n�>]q��v1��W�{��R-��	�ye�g=��+H����rW�G�S�m��Z�"#B�&�(���V�P�T��^�ڤ�{+�;ʾB���v}��%n⹷���]ʥ�S�]�ܝv�<�m7��K�WEk�v>s����B�dR����W]��A˨ȹ���f�Lɜ�1��s���G ]ߛU`R��7j�Bu.���s���S��6��|6hu����up@�c��X=-ͥp_|�\JK�<��}Z���w���M���1
�&�[���>T��]H�X����0�)�*҄�A)��_�����i�>�@�����Κ��҂��q}���?x�Sk�jah:�6~,�\����Z���b��;�~pL����&R�����K<��s�)]䰔C}\������_ca�y�_:9�lT��#޺n�E�IP'�������n�� �)$�[!\*藙�j��3[����苂~q�J<�������AR�vVʱRċ���2b<ٌ��ѷʥ���6(����{���5B׫��'�2r��Ɲb\�ގ�ǰՕ^�p�\�6�.w������1YP��݁�r^
L?I衜�Ve(j��,mT>���fb�X��W������!��T~�E	����mA��:�7bg҉\'לs/�?�6�A��\R/��[n^w9���皥������렱o�2��됱T�'8��c��n?HK�]M��T��}�H/�(U����{�;u�[�o閠sL�:�]���c�b��u;1�2A4>�T%�I�6����}@�(v8�.�Y���G��T���M�~��e�i�C��{bd{\�����̭Q��[�/�޾��L�M�F+��?A��Π������%�a͂v�X�︧gr��N�vdZ���irm��#W]v���]��%󥠚s������`9,[�Y��C	�'^[�5�۬�D�����l���)O��b!���,�2TOy�]#��/eQ}�EJ�<�ӷ��P��\���ubZFs�X*"�t��_�y�Y{�XT��y���{������zx!�E���*�Q4�j�D!��kE�����1��{�׸������[|�#���Ǜ��h��E}U�j����m�߈׀A����Wu6	�N��5�8q��Yz����mu�=wI��Ϋ���Р�W�O���H꿟���X{�3M7ÄN���=}Iv���/���P#�='�;D�?��-�]�bz�é{�L���y�VcY2/_�<i����d��IBf����q��!�`pE�MC�ʩ��ɷ*�'��3����At.�^y
a�7�yY�׬?��GY���0��h�iQ��s^��2e�X�=b��g;f������^g��M�_i�l�}�{�p�/m��d�N�5E��Gr�r�V�^�ŉ�`�s�l1X=��Gή�wA��:���]=���Fw��[�k�7u���A�=K�g�݂�tֈ�ك9{Z���ǚwq�ކ�Z�B�Q�R�y�ONe�\wm��?y���1�D��*����͈]=�A{?BMOa��2�\ M�(����w��r��?�H�G+P�0ٱ�q�$&a2֫��(�\�.� é/�H��:�̒���uEZ�����B܇n�9�\c��fH;(�ʸt������Q�+W�P��E;�Me]��i�{�0����ۘ��SWZ�:`Zɏt��j�RD��.CwI"e]�-��;h�.�ͤ��rd��.J5�Ȃj���k�^���ý&cl�&4r�7Ou	�U�������]�_��,��,��б"�(1M�{c9�gX�`=�ҭ����}OH�S%<��S:��B��:�AK�M�y@p|�Gs����q��6�i-)C��{��u����;�َ��e����^�`Kk8��٭�����$_�u Ӭ~��-JVyckN�j+�D>s��=�E���A=�2��w�V��`�"�K�|�u���"ଢ�E`�����k��w$!y��.N�ޟ�뉲�Xʞ�凤�Շ��1E���f�
#�adȹ���:K\�V�&g�X��f��:���ù`NHwi���:�ŵiK�"*Sa�����r��&��f�]|��М�L�y���}Y�]q����W�VŸʲ]D��0;~՝��징��l��@�d����i�př�Vkˆ!�wM��(�l�!Uh�Kw���p���	���Uf]�q�cf*v�vH�z���j�4R���������9���Wׇ���I�*��aRa=�&$9�S���%��2�U�3����G�h^b�/��}��>�[�濚޶�EE�H�P
�����("P@�Q(6iҦ	T�Q���&�����NS˳�Y�}Vda5������8�ז��f��3�z�a���b�1��<,� 2�άU�&��ž���zm1d�0M��\է��Њ����s��S���5���v�-YPN���{�t�ѐ3F�*XҚq�\�M�s�iFDM�kcj�鹍*�Lv��_��3�=6��oU
Y�W��r���')eԳ���]��S�~帳Z���
��1f�;�)f�m-|[9A��[)+��b�%�9Wf��Wrg.��ᣀQ\9��3�����j�Y��x:��:���"�}���L#CR��ha�PB�'
 ��t�-+��T��|Oّp}x�(!�#�@3]�pt��͛QN�:�Rߦ�)
g1��N3�(ĺA�[�}�7p1�D�+C�h�X��]̤�R��3���Dq�t3G��	eؽk�$�G]J6of,C���ݡY���?=���،�%�ѧ2Ҙ�(�B�e��� �'c�܌���ˤ���'x�ݮ��ɮC�Ƃ������1�[��bM����Nʜ��!=��CYs1�*:le�K���l���q�7�,el�lN������:!|����h�M\e���=p�؟'W��?�ս��k���<���8ξ+
���r���ĮOq��g R�Ӻ`�<�p\�.c�iH����ݢ�"�V��1V�k�ⶮ ��7}wP�����:u����8��}����x����9lY��_�|�	�'7��^@�ﺋ��:��F �˷�&�#P(�vR)� a��OM4��g�Q���\�j�0-5�������_2�� ��]�5������;��љ���^�4��-�����qc��ܴ捘�P.�J&�W��v���N<]���r��~G������M��8�}��b��Li���'�������{ˠ:͜�,�u���҆�T��~��1�廱WW�Q5ԥ́1VK�g�T@W�{{�}ļ^&�챏fq.�L��
���elIx;�d����r��gԑ#��M_ϭ��)��>�f���-�Z���8߾a˰��]>����Z[ݱ�`u޷�c�x�C}����:��d� �{{;�;|C]~���_��$ I����XK�+v�n��K��Z���A�}OeX��xfe�t�o�_w�2D�:c��AM��~0G��� �}���Z�����\`�k�%�8�B�~���N��E�ǃ޿O�M?p�����8�t$��b%U�~̝�v�UaN��F~uh0�W��mc'<#�]=����Ʋ�e&��.�<���|�,�ᾙ�m�r !����'~Y\ǩU��s�>[E{���+ȱ��l�;��A���Ƣ�r�D�UH�,G�>,��"�<�ůp�D<�T\UVO��[׌�>�z~<�r2�K�2ng�3D��ۯ�֝�a��u��,7w4���?��l%ae㗻9c�޼���ql�J�:��;���i��uP�fi��_u$2���\[���p�5�gl��=y-J�Anך�/���?�a=��|m��{N�.L���Q.����_���$����}Z	��T�E㗕fN�����"��_SY�kb]�Q@`�Џ82�И��$�tUL4g���]m���-��[wqZB�=�,�)�[G��H56��c.��+{ҬWQWaIG�w��p���;kƃً���t�[�,GUx����(~9��'>]/�t~�g��]�6�wI�r��*���ٌ���'�u��{�*������;{�ί�{�����kg���X���~"\7t�+6����)T��c6�Y���v�b�=�1�Զ{f�U?]
��k8��гMz�J�ՆW�[����PI��~vI\�0j�MEj���H�5�,��v&i��R�'�L�_����i��o�	/�2!�e9��j�|l�~����|x�^�
3�0��M���WR�%z��c5�x#<�[�Mﭮ�R͙�s?3{�Uu힗4=�2ā7l��~��f�~�m�P���݅}��fM���oj.o��.��D�u}v�q��X�� \��x�B��s�T0/j�
���$8���dQ��k�3+��-���ԗx7D�u7LB�y�!X񥕃�*t�`J��V�rú4�������5��|v�^�Ev����`��k wu��@F$Mt�§�(w:�h�JLiӪ���S�嬭9>�Q�1Q]��;�pp�*rT�z��X!�8�J����U/����t��.���G�7A*�X,W���6 ��'k��Ή�d"�fr�{�ߨP��:�JS8ŔK�����@�k�폺�3o��1�"]\17�������t��}[��zH����XѠ��[;�j��y�nH�١���TO�Yʦ1�ѧ[7�����i�]O`��b�J�d��
z����c��%��kzj����w��P\�D��#���r.r��$M�m�E~����w��X���)�ؚR+�=]���t
��'7�b���,tO���*[�*��ϧ�r�]N������IܝT�%�:�P�g��h�?)��c�|��h��df�pYZ��}57�f+�d���x�F2���Ϻ�㿳E)�:v�*Ш%����-���\�J��*ql_��,SE 0�u����2�=�������n���%yY:��a=7�H��ܖ}k"�bAG��ka�k�v�t�y���U�;k�^�`���x���p�7�y���DLJrU�mk[A{�b����`�/�r�X�w�9_Iut*���]�EsN�� ��̈́�ǈ�Q3�s�,Tf���g^�xNX��%��s�3���Z�E�l�LM���r�@�aŐ�΃���X�0E���@ܻ[wԝ[?�	oV�[�̶�>�*`I]Lj$<ʕ�m���3W��Q�����O:���g%�z��x��+���v8{���!�����J��y\��b�Nu:�%��]u��)}$S�k�%����+�:�e����`�*޸����e�V��$A.��"���7 [��;�6�0�6�g�\cv���N�<�?�K��:�@��1.V!�o�43WAGJ��ô��}���f_��L\;R@ܨ�������uH��#n���J-<��[�d�������#���٩�I}��z�盾�1��o����P��l�QN�c7�j��2��S���~����r�~~+��]o�0���8���/z��m_�wmZ5~�eq�Q����ͽ��Q\�+:Ҏ'��}>qHCW�.|i�2��Ь���*���X�c���>H=9j"���������<d�3�]��ͦ�l�A�b�i#<k�%. �
>*j9�{9Jf�5����#u�5���&S�)n����Ț��0�6�<��r=Js���z���׬�5�<�6WL{ܙS�4S��0��r;8(7O?fd~�b�W{3�G�~�Ρ�}A���i����������[Q˶�ƙ�}B�0P�W��'�f�tm��Q:jy]=Ӏ#s8yHW5����+J�Ú�
�>��gr(�7���#�sB���/���������h�ˋ��ǯ��*Ӳ�$TL0�
�{������n�p�8cޭGw��($�	��5e	b��˻7b�]��of���R��������0J(�n D���U:�K�����ۓ"���e�9���ɪ�ɼv7����7���üM�oZ̕�x1�r�sO��J>��#]�K�u�b����6�O�o�e����գ�6�uT���T+�<*��9i�G�"j��\���jM�v3y�p�\�ˀ�_X�>�|��]*�gfiԅv�1�ꈀ;�8�|������>	����A��d��G�-�7N4d{g�0F�K���	��o��.�jj��u�=��_��"H�!7�I�=S�}����lXI�ov�b�V�R{��lzj�F�x%n}��r�_Z"*����"�!P{��]y����(�C�n�{���S�������5�7�ט�*���z�s��f�b���/����v��lfF�G�
�Yx��u�6�� �[G4��+Y���,cRI���9��\Wu��H}9!���,�{:�y�W�"��nʊرD_Oz��VA+۰��a9ӛ�M�90��~����!�W�xD�U�O���@W��N?�ҿ��7�;���>�*��mR�H�<����L�c\�M|:]�[���о��|��/��O�)�p��0<,�8�,��{[��uP��S<Ay�\�J���Ӻ0#�7d/!۶FZ��&��M��{Sf�Nq�*ղ��P�SqV��2rU|qWX9i��ë ֫ww?ֹ�q�å<����AY�� Y�[І�mTTI��T�=u�2��qvK����G;6����a;pu�������r-�o$�1���t�ҷ�a��ˈ]�7��W��v^��ú\a����AR��,c���$ě�A����
Y��ض��:*D�ery�L��Pqe˷2U�2"�wNVc�1��ތ��׮��q*���5�Iw ����_v��[	�����Om�y�0��Emt��\9��Js�}u����g��_�����ʿ�׉З=A��A8�x��g����H�G�+��w)��g��T�¢ y@����y>���Ƈ&��~c&�V/v�֣g/߿;���o5 �]{� ��n���^O���:��!mgz���cu�6"sΖ�oH�\���`�@��Ԛ�>�wVY�d�u�8�Eu�_ !{K�R7��A�7���VO����U�"�p��j�o��e|Mi)g�dH'B��~�~��u^����LT�x���6�Z�}���!]�V�'�k�ҟ �KOޒl�95g��pG����W�*��&��_m��#�9&��������b�������B/.�-*�عz�5E��Ddo�J��u�3��X{cmӾ�&�<�b��7C){���H^�;|qO7���+ةv��8��;o�SB�Ggd�?�m�ו����I-[���Kd�S��-wQ�ʤ4`p}T*B�d�5	�;��D�:����|7;��:}�F�Ty���w:՜�p������ox����)��mq�p^���[ߥA�H�,���%�v��uM���t�����r5���\���x��]�T˩�j���5��^��}�\6�.�=���x�f�Y���:�ui�t�}\�6��<ze���J'��T��K�Ү���dTI��fR��ޫ��u1��ky׾t��.��V�o�|`���c��tؿf<�l�\�;4P��&pܦ�]����������
WW��w�Fd���)�n�>YY��.9�^O��Z�O=�ϝ�:2s!��2c��hk��S�G؜x���d*C�(�6}����w��\�G�ÌL"�_�^��>��)�C��7�:����ް� g	�#��	��*׽k�{Z}��9��>K1u,�}�c���g�1�������R�T�Ѐ����Gqu��U�::�
��|l7��*��y1d��>�۸��R�w��f�q�}��x��z�������:�w���J��ֽa̭y�w�G��E���p�9�^|�≹'�<"��]��<���k��Z{y�Y���-R���9R�R�&�t�<���(>��6�G����.�]��) |�>kr���a~YB�[���R����E�VjQui\��7��9,"^5����7�)�[�0-H|l���O�v��|��V�+>���ǝN�\����s�$#�ո���6�+�G�w���Bbiif�ܹɁb����3/���ғx�qW>{�;�b�\k+V�����&�M���:��ȕ�66��{3�6^�����D�Z�&|*R{u�7�E�i�L#��YyY�v�r����*M^����_z�@`ư�A�}���aDуxǫ���b�w'��[l��M|@z�ugN�<XlP�]V�U^���!
81��^�G�
�_�#b�H1���^�o�SU=�=vo�f-&|�����7���]o$��[������@9�V�8�H�l���6�nT� 觙Bf<<��]��u���;����bbĈ7�S)�^���4��xe'��y2�%�PG��;`K�('�\up|��$/�U��؍�:�H���X�>�4���x��>#��z+�S]P�ޟ;�ߧYK{SȌkS����}��$���l�+���W�r��̧j<6�+,�0[>�az�^���)�[#�:��׈�h��5����֍7�޿k�+�3;��Qk{�������C+ �0.8�	�я���f=��.>��TMK���X��w�)���V�;�^�|Ef,�N�<��}�hd�#�}�s	��	���Ϻ�c��l�Pg@p�qN�θg��O��i�`����o�:���
���*A�y�`V����ˈ�o�}�L��J�+�|rr�Ŕ�K�ܶ��s�OEF���lU�b��T��II��y�����.D���&G��yY6��I$�@1����xr�]��j֖��qP�Ҫ��vXjb��v��g$�V$ǒ�",u��n��������ٹ��VUZ�����y����wh��m�E*J�8?h�hgt�%o��&�ݼ3�S��D�*
 �G��Q7���cԍS>�-�EQf�f,�)���L���M�V`xؓ6�S� EEċ����F9�<<��-�i��q܀B
{2�M�(a)�gۙj����A����,�S�U#I��4�V�/=ΐ3[(E��6��B\iz�{r��̟k|7�xL 2!��}_�ϱF:��\���k�pDNԞª��.>���І�*�<�g.����ѹ��v
��WK��w�Wq������e�\��J�Om�������V������b�*��]h=��j+�"�Q~(z_��&��zj�f%��t)���_%#e+�R��vng������D��n\�|�Qΐ�9�Ҽ�g���ҟL��w<��\j��{��Oe	1��f�Z�gax��G&�b`v�NrF:�弯��d��Z����0�`%n�^ �%�,��_/��_n�+�)���L8�;�SC9ߐ�j�W7���PO�t�H��B7�ѐN՝U־s\���eXQ��FH���g����z5l~w��p�ܧ�@;�;�j��~����~�k��#���/%p+R�M���FȊ��V��Y�M�h'[���A8O��׋7ټ���:��9\5���k�ʴ7��*�PSY�S7��{�����f��ԦR�����n�s�7�W;id� ]u�y���c��S��N0�n_�r[4��.>��8h#�G��wT萁��>��Ȗ�JV0�Zuqr2��u�@Y����:b�����M��ma�{����7��j���z�������Ź�z8��
$������:�d��	LW ���c�F[��k
�)=a;��DWX�&Uf�Ѭ�(���g�Z��Iޮ�d��uCrXb�+#���;F�o»�q�e�pH�a�
��{��]��w��E�"+�����Ύ��j�[[�cw`(Ư��N��xz𯻡�K�\��m���)���]K�N�zRi���oJ�`�%}wf�Ƚ�+ �qT�8z�U��lX�q���_&K#=�O�WSy)�DB6�2�X~(��ߐ�am���Ź-�*�ǂ��///���MAUc�"L|-аpv�Nj�U<�s_�u<np��J_9�s	�\{�.��2��f	8�����1�z� m6<��"����&u@俣^Ɏk�N(��}��ABV������U��w
�-�g�|����*dT	W�v���e˱w��;�W����m����kp��I��"ǎ���ݫ�`S'�nxF;'{�^��|(���pC�ԗ���A6a�v��/���,2� IJ�.�n�Vn�}�j!����tŴ '`���҆���f*�i�h�˩z+@�Xp	�h�r�h�w��ahu�żfu�i!���u�Q�7���mu���>K4KF��p`d� �=��jk�ǧo���3c�j]�����YGY�PӾ4ۺ't�My���5��$��"�w��n���P�3�V��u���L�L.��EM'��#pЙ�d����1s<N�l<��ۏZ���Nk����#V;�_����d�,G�v��Kt�s$�ĴM=b��怙G��}�1�u&�:�)e�yu�o��.!�ь!Gh��f]K�Ѣ�+Ʒ�y)J�0V�} �n�p�Om$i��u �,��as9d��oj\8��T�νhm�U��^��Iun��H��UʽU�\�����9pK�C�n
I��Xyws��OUi��.��`se�)WWa]��U���N�Vt��Kh	.R�ղ�a��A��w��.eX�5[��K�d��nf������;�(ٺ��k�f�R���}| ����A���Kr�غ�lC%�B�'�iV����v�����;�8aM<b���&�S,@w-[��+1%���jX��Ⱥ���*p":L�^.QV��Q��p#���i�*�I��w[%ƠW�;/��h4@gwa�|��q��s@���Q��׆�����
�Yu9�Z���z��Y����� 5(or�9�2V<�+7��<��
HѴ�����8�:<Hm����3�R�;�ugb�@��<2���w���P�u�$q�P�p24u,�����h
|�Aᕮ�t�u���~k�?'�h�S/��p�^1���fN3�y��u�̾h�P��H���dK8d�^+��l����:��l3
��PuAƳ��.�'vPX%+C9z�ͮ.��������P�OL3LxJ�������٥�)�6��i>�����h����Q._StR����Z�V��C�v�jΑ�|�ε���˜�49B�c��Q�7+mS&*��_|�m^杼E��F'@��tU ��[9���]!V�>�}�J�#ۺ�t�v�mJCvK�j��N�i�[��`#?B�RC�ь,��U��μ3�Pܴ�x�[��ꕛ��}�n����O&f�ۑ�_�TӼH\��ԣL8x�˹���쏦d�jʸ�F_<��{��+x�a��0(�C�FPۃPze�|�B�i�~�:��׮�Lq�s���r��H7lS\���n��TL�3��J���U}46�Q��&[��;-�5z%Y��k�-�Ο<��.b�ke�@��%��>9��Zr��Nk���a�cgLU�EXHARLV\g9"N�0�Wzѝ�nԸCe)���| �񭗖W������Oeǂ�EJe�Fun��>�֌H*�uX��Pw���B����sO]�qq-�ӱY��p�ȳ ��Ѽt��[	\m�<�	�iG\�"g�#_w��X�͇4<�ū�:<MДP�Q=>%���~�[v�5�+��.��P�V�G6����#�] VMzE7r���Փeu��@�-���~�PP�A�dnlLz�m>��u���f&=xlEB,GR�α'le��s�g�-ha���W�ϑw���JŪ�yË�0MFv�{�`IK:EW��	��+RS�gol0U����o�c��EV��xk�EK��*/��ʖ�*�K��%!NáK�#@��_��z�������݈�e>����X�|���� ��@Q��:���ƛ�i�7�{�O,���4S�~�����ٔ�𥕼���@��3<	�C��7R���h����}��T�oۛZ}�֠H�I|�n���O<.l,����n�+�#��/W��S�]E��b�����Q�K%�Gß��꛰s?��3?7�C�jx����P�>�q����{梼l�rcw��;=b]g�},W+��M�f�P��v�u�o4EV;�,A�^��g�n�z���*���n����N�5���<-�4��9����u�>�ք"����MVQ��d��j��kG|s�R�����K�f|
���Ɣ�k1n�c��6��p��*�`w�YӪܲ��l�ժ"gL�

N�Z�Ig�j��'������5RG�<'yJ�z�Z}j�S�Uy�w��YD�Չ�m�]��Y76.�O ~�xz���ǒa����M���ezF�6i�r�{|o��_��Wl�����f�m!rB�{}��=_9�,���l�,z���UC2��1T����Yw'ױ�U�����8�`a�z��;��%{Ԫg��N�=R{��A{�Q,e��K��*�q27��,��'����#N5i*&���Z��&	�7m�M)Q���T��������D�R��f�w���xV`��_�����3���0�����7ЕŽc/GP__Nޭ�m	i���m��r�D�}w]!��ѕ���Uo��b��,�!LL��+W�;M۳Qr7n��p���=��nw�Ǥ���3l���&^�D�K�m�P&t<-�H�X'�ZϮf�ř�1�Jӟ@���a�\��8�{�0l(B�&�Ƀ�|.�Ofrw��7؋�C�� �ة��kd��.hb>���3�Ь�4=���R�����9����W޽}@��7���m,������=W�+�z����W����ʾ.|�R@�熞�]}�z���v��e��#/b

g�7�7+�I�o�f��u��F�F<�A���,��pYqBM"6�֕����m �m|�$��Hd켊�aͰ+-p��VуUб�0^�G�Q�7��*��J��CQ;�v	�����XC�#s�e+��u�SঌڷN�{Q��j�uȤ+_V�6�L��ڕ��n�>��j׺���m-��fJ����O���lߩ(�h��k����k�LxSZ+g�.�����1'���T8���m��m)�y��~�s�V�7�	v%�}t�^�֮��_���܉����o�u~�cf�V`�ZupŜ��������2�����1�Q9;U^��!�A������HO�d�\���
��`�r�B�˶�ұS��~��ϸq���W+w�`��p���ٳd\��o�BYk3NtQB%�����⹍�UhWw�r<�I�w��#}雌�w�q���f_ռP5Yg��ƷA�X��嵉��ŚS�
ʎ�?��lr�_{��]�����3���.=�YC��N�4~Y�&<D2eg��������k��3��
]���ō���Wk����K���jG��?�䍥/�G�2���� �]������ہ�<p!{jz��|D�V5�F���rOh�baa�X�3�=8���흴i�o�^�Y������?S#-W��-��:�G�0��F@qNq�UljRy�BЃg��A�Y�SD9EM�> �y��3��Y��
z3H��t����k$`���N�����Bh�T-_fY�txNc����\���\�9���!����H4	��C��뱆���0W�B�J~~�\܍���K�|��:ʇ�Oj�$P�D��a�9��\���Y1̝��ǝ��Gs�?l)Y欄��'y�Δ3i�i�ʛu|��Ě��ٚ��������qwա>��繮�����{�k�����U$ʚ�߁���>����?˩	b2��o�4�}P��F2_�+0��bx�?o�3�Kk����E�5ޗ.7��v��0�k�wn:5����� Ԧi��2<��M�C��p� ʻ�s�1i��6�y�87�����W4��st�[_>a���F�L��z�Z��FE��.!	uQ��0���3��adm�'8�E�Kʽ����,Pm~6�^���٨t�=Ld�q3>ɇZF�!���������[��CP�c��2��Gx�\*`Y�ACp�F��-�7l?q�m�qj;]���Ӛ�E�6]/ZDj�NW,�߲`"����!����,J~M(Y��{���b�����d�J|��S}ᕥ��d\_�C��Z������b�DL�M�؜��y�j6��U��̊49᧫����E�?�YHW�����[ ��� i�x.�y*4v��mx��^�V���qW)�D"++u��e�[���i#I����:�U���V���������ȅ��v�aF�1#Q2��ْ#�*Q��e����j��B�MX����)��>�e�<T%-�hW�S)�|�~=eN�X(U�fQa!/�\�+C
abS�m%p@6�Q��'����`�V��[��K�(���a���������#�x�u�4FR�<���֪��䣒��=A��� �K�PA]��n�t&���SN�p�D�>ޤa��� �S�Կ|s��k�cW�tH�'C��V�l4���N�V�V*�Ԟ<�oY��Lv:j�$���Ju�|
;�7�����;���)t�V딬U����!�M�C��7���{yJN]��8Y��㽺���I�ĺ�DkSYO�X�[8�F�|P^(��%H-t�MRUp��Z]��
�6h�l~?������l������A*���Mx�9لaB�>��0`_}���XW�y��D�7K����j��c-{	��s�]6����IA�8z�:�?Q�S
����Q~x��!F�#z-E-�٤,�dT���I��,բ�.�X1j�ZM4P���f:�(���I��F��:���4A���L��p�B<�ϱE���N�sۂ����x�yQ)�U�L>X<"~n�-����`�=B�T)D���V��΃�4��p5f�؟z�������J���K��6L�חbP8.-���q�L(�T��9�e���U���Q;�&�2Z�W��@��̶:!1d2�61�ښ��R�}~��Xlz�����h5A{������X̤@+ʎ�W��P�B��看.�#��N�h'�GS�ܲ���#�	��`z+j��$�[�T��Q>2B#d.����I�L�`�2�.# �O���&�گR5\�I�Ε��|��e�YHo��嚊�N�ȼweO�������l��몰!x@���b�:Y���v���(��,�������(e�L�L���?�/������W��n���{�,U�F�����"T3s�{�X1����׶Vy3^TQ������vxB�<V��<Z�'m״�&p����xΪ˙u�����>5i�,�{�����C�~*�m��XL���������_I�4���+W��O����5sHdUn�υ��y����U�{���kD��}�tz7\�/Q���n�$�QA�H-$�P���g6���Y���Ԓe�#OLr���r65lt��ի{mT��<]�Q�`b�wcYw�Ezi/������f�9��n�(�����A꽮�ɋ��Ȃ4�:g�s	^���d[\�ܦ|z�\
�K,�CPT�ܭ��2�k&Zt�6�/a����`����!*���I�h�zT�E9c�Q���MWĪ.#��,��mF���\Fj.4ӽ���C0ō��Dpd��;�~$�
��f���ҭ�mqA���Q�Ѥ��k�k����ʼ�,r�F���1@���T�*!�(/jz�jZ�9⨸�E/��~�՛���b�a�)�j��}�у��ˏ�6HEz�����C��UtЅ�t�Ҫ:p�G�0�b����GV����{aE}21-�a�B�����P��7td4)2�&����\K�3KeqMq��ڭ���yA�E�k� n�jT�.���@W5=M�]��5����a��bg�2�Y�Z�d������[wBZ'�4�4|��ͦj���slY���l9�k�\��-�����1�Q�ɐ��Qj�R�î����Z����6m�L͘e娦L�m�s��ɯhRY@��N��z��Lf�M�91ы�67n�szS^-2�-p�q�#"��;2`�T���ڲ���$��z�byp/9�V�w�G
?�W�
P����d����[Nyl����F��\���!Z�=��	�G8z&��
Xu��@�篘�ER~>�Ұ�S��.!G�����L��� q*ͱH�}9��ɜ�H᫃��c��Qj��ai������j�ۨ<a�V���GO&�+��|RRo�i�Չ���A���wZ�5՞��������$|p*I��&�����_@�D�N��A]3��N5|F�q��6��d����	@Im�����Pu��Et*�����ʤ��x�Bz��n��B�0��	5�v��!��B7�6�h�;�ML������W��x��x�)2��h��Dθ�ЄT�4����S��OY�bဢ�4���J��I�9�:���.\O�� Mv���t�9h,�$�ۢ#:�U��_^���`�p��IQ@Y��\w]n��]*4�#'�.�V^'���AR�E&[]�95T�`��͖�W1���%yd�ȨF����,559W	V��������?)��f�Df7��E�]t��B��1�L�m����"�wPb���p��������VB�'�ګ�1���2>TRD{��,l,/5�Vw;�`�*�pp�z�Y|�	�{���IZ�&��F����aM�ï��7^n�͆>\U#�L������*_�_'V�)���=�y2@�JuA�ף�s�W�Skrb��*ZtȢ;��e"'MWT��ڪ^L܅f4���A��}D�a����W�	��H,�������!z+ԉ(�-U*(�;�au��k������W0ݱ%�B�;jM�j�U��LJ�9�.��:э�g\���<Ś��y~�VZU�nP4�;����;0p�b�	��D�",��������mn���F��3�n26;(�%gF���,1���_��z�5�΢�D(�%#8��b��ႃ��~׃-�:2Վ�1z�ʰ�9���'\��e�r����mmA�{�`y��k�sFp@��kMB�	�!پ3G��aMC��H p�"SY���YS�;�F:����!공x��v��jC��L-�7^�Y�|�Q��ƍ��/���+5e*N�5��_Ew�K�i�R0*N�@,�8��q�1&�:�N���C�]���7�rgj����N����z��a��Xu9�QS�n�R{��o��n����TS\w$)��{�O̮j+�ر�?G ���4iP��^�C���g�_�����I�q+�bf:څ�!���lQM�QG����)��޸��%��P�w��[���l�}K���������������F
�r�\�Gka���J�����z�{�<�zf�s x=���C��K�x�ϩ�&a��v�2;��~LqI��$_	(��Ї8U��-?��֢s�5�{tI�.��q�G��TXF��1����h��+�-L�k��y�L9"~5qֲ4��l7�����tW�}�Qgt �����	v!qAD�5J7A�5޽��m���(Zp��8�'М���^�]C=�_]�g��@\�^�Q��<�b�u�8W��qC��by�2���TE�s�rNe���r� ��Պ�*�bO����S���7ȅ��X����9��o{]O֣�8�R�����ӥ"��y�	��VF��+ж��EBC��p5ߋ��r�,O{���T׼�D��Skh33�d����~����C��ܹ��������^ە�<0A��>�PF`/^F��	��֢Bz6��`�=9��1,���P�Z���ٚ-�r��޳
ч��t��8��6î����d�G�v�U\鴲s�r4����]�q,��8�xJ�񗊟�����1K(�v�Ac{��PѬ��͍��Ũ�(gK{yIYX�Υ�v;��\�����ǹKJ����O�?}��⨊|nt�0�{���=�E53q�:���ҝktYGp%����wxG��2x-��c���}{6N��?�}��)��ͭos��vz�C��~��򈥒�%�N߮9�%N�m�ZMF
�Q{"�"a�1�[~^�_Q��<z*-l���9�{�0��s��X�=���:5��'ݵ��e���w=����X���1?Jh&l�^����0��ʺ�t��.�~i]��]S�߸Z�z*��ŋNq�x����⹨���-����a��:��m;Q�:�߶
���d\�;��Ĥo5�S��3p$�܋��k�񽜟$s���Y��Z��z�~S�jF�~�H��|������vjB��dLl}=�ݗ0���RT�b/���9K6�ZP,�2}-{ٌ[C�Q�z#{�K�īK�^y٪dE�4/X5=��ډ��WIB�6��`�1O6tA���P��a�徉.���<�>�k�Pf]O�ȼ{W�x2��Mӯ���e�b~".:;�,��B����5�b�մqT��n.�Kn�*	��>�g�g�o�u}D�Y����}�t�J��ϳ/�
�J"��gm3��T�~��N�f�gOvNJ�Z=)���.�i��nS��,�ח*`舱x�3y__�}7^�4��r�6.����.L�y�5�;��Pi�;M�
�O�I�顳-�S� ��JΡ�Z�GW:�m��/{ʡo"�)�-���T^'x�_\�3/P*��O����Ȥ�f�x�!LuY��J^���÷µ�����6��;*����I�ug�t*{#W��1��@��+9\k�T��U��|��x��~�"�8l{�w�׺h�x���}I�K[��E���p"{���G���C�'��ꇗy(���|��~���oQ�7���甆��Dx���^���"���c�t�~iIV�v�@r�K���������>�DiQ2�+V]q��Io�a~�6�w{�*��A�a�9%n�n5�/�~ ��^I0{#',{jwj�>��#�c��b�':�t�]o��ڠ�S]J%\�c���4���܆$�VƁ�fؖz�M���$ڔ�ˠD�¤��h�y�=���X��ϱ���
��tɇ�S4P��W˥��� n�8F��BW:�}��N��lF�"��&��ɽ~�U��.v��|���`TsAܶ� �	s����K���U�����U� �o�U&��J��ï�̽l��W���O�(7��ゾ��~O�M�"�vn�~���*aɼ�]��D
O-���݃�ۊGG�q�K-j��;ˇIk�ޖ�#o�X�`�eѥZ��e�j�-�Α=��Zս��lZ��M{�|	��Գ�K��;k4;�����˧v�/wL��v����j��na�	�u"sj�ZR��r�o��)��0�
<i�D[,��=�}Z��ajm�V{�޹6�Vyo*'Q�V����|˺;�����=)����t���z,gc�W���L��
�`���3>���N��J�5���N:�g�F�q�s`��s�*�u=FQR��n�:�xZ�k�y9A+�~�Ȅ� jlŪ��:ܙ'+���k煂l�>�Fp���o4Wev��(����o0��G�2�����Bu#���o^줄��^�oIR��gz�Zw$BV�Z�7vLo��]�u�U�+C��������2�_s�ޡ���v6�ު�iMv���9��g�-1E�O�ã�p�,TH��$-��Mk�����٭�y�}܁�V+]*wˍ�s��7;�J�anA����㗡�f�}t��O�:����3������8[��}��]BP}aga�o[�o���*��q7a~�1��;]X5���6�j�"���ý䤵�r;g�y�u}uW.w1��h]�5[�� �z6;��FXĹ�Z��Ѻ_����؅ժ�;mš����s����Sb��n,y�j.͸�]�z���IZT:Ǯ�7��+aX�����@�;P&%X�V��!�E=�-=UnْIt{�)oV��"6152��Wu�d+y��ܘ��"�k�t(�[m�%& D��m*a�I+�O��1B��MS_QE:lΛEf�s"}�g݀��]+%)d��V��M���K){�g�Y�<t��S?�"j[b	f�5�0e��Ȩu�댙��1V"�Z�c��	�Ie��(�7a��T{u���7�6�2N����6M,��Q9�[�s5otI���jy��]�� o�����'�=Ǚ?�+�<��������U�f
�H]�]���V���ݮ\$�]CUj䃈_^*#�@�9�Ԟ�\At�TZn�6�뱦��,��\ۂ�w����))V��,����u��j0�6��������8Kv�1�v>g�l
G
�gv-S�	�iLk!���*��4�a)�To,�P�OE���rב��v�	��3^�Zq��C�I�r�SlG��K�˼�[3miY��0+��oM�ΙO���6��S`��郫�Ղ�΢�K1�Le��Yt_���b��K�jX���E`�ͫ�]Qa��%e�{v_�����X�}ac'D���r�^�֋��v<�����˂�)��+o���1t���Kx���[���M[|�pe�ט'=��-̺0;DU�������E��cNLNĻWy��y�M,���Yp;$<5��J}ab����af؉(��M��D&�p�֨<�kw�ne�n� ��흣(j�L���6j���BVgSΔ/��o&w�Wv]7-P@ZiVdx	�}�I���b��v1���iM���W�UUo���A`K�ʞ�k����u����`�;|)�s(7*�`3V��*�kLg�Y��8�G+u\ea�v��O�U�2g.�i�o��V���֎=��J�<�*�U��'jZ���Pڶ|5g�z��O�~��rQ�;mv�==)�.�ϮB>���EEn�?J�m�nߌϽ�:v�E��ȏK1{��p3J�w4�Q�O�p���TG�7QPƛ�Y��Z>���X�1-�J�C�qzO�4%�d��$��q�u���S�wBb�]�5�y�yC��q�^n�5�Gz{��d�:�O�'3��rD� \u��ߦ���/,Z����L��\���ՙ9K��;�|Q^��H���[�K�_hal�)izi�٨)>G'2�5xRَ�z��s]9�<�y�S]�����WJ�>vw�{��=}nNzqg���wb��o�U���Գ�M��"<�^�F�#�W�<�v-v��I*Q��-�"�9��w ����лT���ptj��aa�e���������������׉�z�b�jU�.�"y���.��pR8����^U9�Hz�,���%Y�n螾����u]V!�=ɼ�Ş�����˟up=�h�k�s��t�T���5O��-��&k�����RA����bE��7= ߻�Oj���R�
8����
q9im�4�o���b��S;��ٶ�#hE˒]�f���b�0`��9
�W����=��`\����D��<��vu�wԺek;�+M�S{4$�Z�ҩ�-�yDk��W��7Ref3����x��g����X��(|��v�'c\��u�8�FWr�qSe������x���S8�)���N�y���:2����we�;o����Wy��Q%\��eu{^��~���~�>g����F���|�Į=�Rܶ���;�b���3x��I0x����q�#�g������d�2�ucnь�?#_�P�	���sA��ì�]�ɓ�1��G���dW^`VP�tB���}y�ʛP���f���|$�H�岛^������,xf�K4 ��x��v�8�	��J�4��g�Jv���kO5C�ɨ��ܸ���#�˺]��Xe�UFE�e笩[bN���-�K[,���vŷ�L��1��X��}�m9f'�����&!�˲"wcP˜�e)�!W��ő��^f��^�F�!�_@`�v��^}DB�8�\�1բ�&.���W�\MU�v՝���?	C�����T"�&\g��Y��tZs���S��
I�Ц�?x`e���߽��sɶns֪�^�������I�]��P�&]��4m�&��;��17x�q͈���\�e_2�sF �U7�ΩKx�;t���c��1Y)�A);�Yya�KpƑ�a\5k_J���Q�{g����wTD��u��jJ�� k����1��dW��$]��n)(B0�8�p��3�ou �=d?eD�ħu���4.�v��sb����8��g�]"Х�ݠ���7�T�Uc�,k"(9��^#�0�"�Eo��1>�i�.ڼwBj���L�S^�P���/�j�.�s{`k-�9�t�M�Ӿwn��C5������	P�t��$����������ጫ���χ�{�����FUQ�Ϡ�_�u@�1�¼ʺ��A�<kӶ�w^HFG��i�ȝ��@y�6���ʋ�c��fapxPTS3tb�!q�|}���u�w��Y���֮}#�
0d6�JNㇻ�F-��d�B���M���GH@�GT�}�Wdܩ}�Er��y�z���^�~�d��;f>y��SG}.�ȼ�6�#Ҝ�q�s���f��[�Q�p�{g�d�5���>�7Qn93��t����s�08��Yr٫bn�����7��ٰ#��v��(f<;�3�:���SQQV��t�>X�L��.�ވ��1�r�P�e��˷�'39]��Z;:t�Mz)�M7���p-�!x�>����,;�m�W�͆O�=��GNx��_����5��p��N�o1�;̓s�x��N�=��%�Y��9&��H��X|ۧ�P��˳�Q�ڵ�m���i������,��#C�$!�0�p�\9��v��Ij�K���a3'�JU�c��&��op��BùS��g�y3���_"s�O��."1��g���G�u�y�6�v�q/�0gF��S]"��~�^!C��>�}	�,�f[�c8W��֨C\�)�	��6xX���sJ�_U�M)j��:�F�1�,=2S�b�������*��_G��������o_�F�z��M���;�L�E�(31ʠG���"���>�S�F�Hɬ@Y�֗^XE�4_�]��v2;���G�h���au�B�̖���d���c�U�:�_4�&c���ӝ�j7qБ���{�J�c �p��:y�tψӸS�}1�57��뱟��Q8*nn�{)�5�E|*.67���VVP��WB��_lɽxl�������Oȅ�	|7��;4� �/�2L�KϮ�6��MD���l{�b�K�u��0Q�VA�E�=iχ��(n�:+ 6 m�)�U�
C�	��w֝��֨P'�'�7��N5��.r�4�xgc�r&��E����D�n�$����ʎ�|��R��WF`��8��!z��{D3�^�p&�5>'�����,��BoTP�=G]�}P�
���Fn��,T����F��A/�n��
#,�W��_�O�*�u����+h�l��#��ѓ� �J�p
�:�[���.�ϥ`����&I'�[�7Jbﺟ�֊p��묣	d��]��N�ά�͉�?nv�kuA21�%�
u3�-n���94m^.!T�]��S�uV.��#�{S�`�H����6�9�9v�o���7�Ҫ��H�W]U�o��.u��q�.�=��pՇ�3���A����n�js��n�����#����r
����c �6��~� ^���x��:3����}�U�e�ͅ?�S$xp��j�A{WF�a]f��>��chٞ�>��s�Vk6��ga˿~P�OY�3=5��@�)B�c}PW�z�L���rSs�����c��������\b�|u��R�+��]����N(�A��m%^�ϛCÉ�;���x����j��/�iN.��:C������s��S��ۣ}��	���w��3�V�I8��y^�]VF�TfTp}JeN�C�{�]+>[�^<��(ZS��^����E�������tZ��t���)k�$W.�:�^�k$�x[tX��1���{y��Í���9����熶� �ߢ�m](��N����}�a���ֺ�7����v�+p�ߪ�X�Z}Z����_�ߴ'�X�o>��9QKk=�v\V��etn�	�X���ܲ��QX��軖�LM	u9��ɼa�l��r_ _.��kv�n�_:�KTK48 %N�-F�\�r��is��Y.:w�󚮍��{^񡜫���B��pu���;��\�$f��NS�v�֢�����/�V=�y[��ϝ���[����l�{nt�9�2�Ն}I	��m��A�v��/�3�(_��}�w�O���2Z)Wt1�ݕk�'3�h=+tv���:#��v�񪋸p��hy^��dP�����7�o/Z��tz��B�f���v�Wb��{!���u�n#;��CǍ��[�A��6�\�3�ܕw%�8�G��&�q3D{@���˸�|Ð��3�k�}A{����V�}���{ޒ�d܀�N���آg��R��'��c��ƺ��\��l{x�3��![�k�¼1�3��O�uq�k.�4HÐp_�ڈ�'��xRw����uC�Z���(�B�拏�K��?��GFm�ȼ�Ϳ�or�1�9-�1�b��Z{ �T����l�Gn�_&f���E!�6ϑ�K�"��S�m}����{31SF�ʝ�ݷ�Q���z.�����,��۠��]�t���	�m�Z��������x�A�ʃ}�ex9��-�h���#Q=�V�ųׂV�ّgR{�d��p�;5����u�.�\�4���7��B�r��<��j����Bφ5��=gk�[�^��1�R�WnS�Kfu:�Z���G�t�VV�yz��͵�y�By�6�f.i�k�:Jk����3����f��2��On쵯��`7R���q���Y���{��cYKo2�����]D�\�g
#0s����;�{���W�7�_�E�D��dg�!���έ��]d��#�7ڻ\s��]����;�mm�f����Ŷ���;˽]An~�s���ǚ�tֶ�jCQ���J:����=t��u����F�:2��j~��{\2��z^J�^��^��B�^�y�7Lɬ8+8+:m
���6�^��/�?Nv̍�!��"�j�c�У�ߏ�c�ꙁ@����尖i$�+0�*���5P��G|lG�0��{��y1�牡~5<��޽�,�_V_L|�����1rƕ��g�^?;��d[񭜁��j�VG[6L��r�_چ�.����*��u�=OL�-����ҪY��1K�����
s�����ڱ��s�;;p�8�*�D��z�~��z��J��E��1dvUt�[�9�y_���'�B�� `�ݏL�*�g|]։��f$^�t�+�}7����]��YK=wO�Y�
��="�q���4���-�&�;����./g߷�҃��vT�U�zx�'�Lc�jY�쨏EKF]].�	Y��ez��+���g<Y�U][a�bW�^����Byם���I����=	�L�O;���p�N�벜/JV7�Ј�f�dۡ�{9��2�b��:�8�7�[s��e��N$.������(6�"!΄�\�\k�k�J�UD^=��r�U�3b�p�${��� �?Y���2��t�i\� i�S�y#w�ؐu��n��g���ho������q�P�U�e�YxC{�~/+��߫��=���~�Nu7� n�vJx��`g�+�|7�TZ��&ۋ-X/�iࠇc�7���>ؽ��Y��v2x���xlt��I;���\�������h���sDLME��� ���W���z�I9��ˉ#���5��V��/oc���s�q/xَ �	�1�ڞ��J(D�z�F��W�Bm�v��b��.Tc���Kd�ÝG� ���b�a9���	Pw�0'��������L�}0&�|��?K��Y���ԣ�W[��K�ٲ�ү.��z(��P�%�1���؏���y�#��ܱ��
����d"W�XZ�(]���Z�ϟA��lݗ%�#��N&���d�Ml�Q�CNKf/wҚSv��z���Y]� W{�����L�ϣ�2��;Z�]���u.4آ��s��s���ݬ��L�W�Gа��{1��YVYu�V��6��v��d}5Sn5"$�#��M7� �צ�-�M�4������̆��)�nU�Z�.���%��h�G$��p]����$�݌)�W����ƘŜ��,'oS}� �3	^u��ۤ����Z���� �Fs��[���r�n̵N��bv������¥�WΜ�hSu�Qkn�����.=wLe4g��9�U���#g���1q�V�^�g޼f����E�̌��/r��A�����ǯQ��i���-�Ƒי�I���?"`����=�:1G��'�����{�5�;���R6	ݩR�3�(�b~�_}6�p���G��}�Ɗ&��?9�q=����H��f�M/&pxg�_Wo��@J�nq���vk%��U��13̚�t���m�pݓ�c9�=CYε(�nbkPM*��hŻ��k�^�`��f�]>j}$���ٙ�s �;&�%��V',��}y�ڽI�˫7:�3�t3�4��6��p�R��������̖���Y1Z�8��iS���8}J-_XE1J�9�]��B.��Ʈyv�f����S�-���zM�g�mx�sk�gև�.�͝^>�+��3@w���(�l]�}-�m�UnS�?���XV�'۵h��͡c��K�����lJ|��nȬ4�1/�؞�Cqe�3�Lԥs�J\��8�P���,H���M~�ӥث�zI�}�K���b�?��TP
��B����En��.bZ�_ٯ���n��b�YW]NVٟ�󁫘��W�Y����8'߻��̮�"����צ=�Q^Ô#-�L��g��M��[����ڗ�g�qåï`�s��6f'k3Y��n�w��iE���.#qm�`�R)�'T�Gat8D��T�{ݗҦ��5,z������sȰ�e*4M��V8+���/**�t��F}&|��phOTx�uMY��OO�8ټ�����B��q����΍~���!��*~iƦ~�7�f��bB6�v,�4�dX��������iF��)�+�n�9��58,~��9�_V�'2KY�-���P�#�=���rǗ�_d]֚���f����c[���)�콵�ķ�د~�����`�7^�_{�Ǜ�^��O.�"�]�$����e��EE�b��k���ǿ�Ş�t菴�?��	🲹|,U�Q4�d`W���s�ۚe�>;�M>n�U>�x��������;A��쉺��9���_�����N���֘x2�?���h��ܖm�HJcY�݉w*�����rsb�zxCq|cmE�	)d{\�Z4�2`��+py鷿42���QIM^�\�����Q�<v]�����k�U�t�ы�>��NLޜg3��7���JE�O�7�n�Ny�u����,;%۫��b�\	��Ib�:�KՏ,��KW�G��+��!�fE��N�5W
��G -�a+�6x�{l�9W�
�]�vi[��U��"F��3:�٠��bل⷗wP�n�s��0+�X���`�N�5�� ;K�ӏnP�z�[��ڝ�]�s�J�Q�[kY�V�����åU��a���t��������>!T�.���C���N�a�r��i�<T���l��f�&���ak�G���&��� ��V�kN�nQ�n���;r��Tȥ{R��[wj���v,��|��Æ_�6P$�w�� +��$�y�~��CL*�V0{�)�ݒ�N�'����udĚu'e�%�C#l�gA#M"��:X���%\Y�ښ�]��o}�w�޺�G9�HI�ۭ��������0-�	&�t']v��C=N'r�R`>�{U'S��_�BO=����Uu�Ē/X�v�$�!�k1��O ���M+�4�)!�]n��t��{vF⒮of%'���}��^�io�i]۴�@�z������5��+�2cP�/�B��-B��&']UӀ���(/�3\>�}�,�J��?b�s�����)�G�3z2���6#�gjY(J�zg
��㻒o�7�+�;�H���o{��>�_k��o�gl��>�"����Y,�VM�<Ϊ��
�;�����6�D(7DIJ��jr +������8�Z�O�Hu�%�K��3���7߲����'[��$�y���I"�>d�!ϵ�]���l:�����~g��a�+���kk]��1�|�$��v���yN�}���Y�M<jN�!���8�n8�/�Q~@�����S�Q�f��]z�R���v���~�;��N��=�?]�:͸�+�J��� ��7s	�W'YO��4��^�)y �z�'ʛg�� G�f��)�o_�DZ��ic��R uʕev�iZ��N뼥i��C�2/Lcl�L`q$�2���/�`��l�/�>nv�HL��7x�Lt�/*)�xÑ�N4����W}��V�Q[���\)��\Q#�lB.�5*�mw3S�w�����!�G��+��#GN���q{�Jثs��"+�K�WYx���o1�Cb$������K۾�_[����}��eo]�i�t8[���WL|�CP�z�u��3u��Z�3�Che<W���:�s�h^����W
xv��t��ʬ�Wp�`�YՃ�-�r=������w�2b�O�n8�Ҥ*]�٨�)�z�n��M���K�=�5��Z�u�s��(���u���,�ؤ-��a~:�4#�Mד$:���o������˒�˯�o0����a#�ԭ��pU�E�ٛy��R�u��4�dX̛����)*ơa�{�K���v-�f�Er���c�I"�	b44�Q;w�pD�I�+_n�5�]��V�=�H�Py�'gL;-�7�ޓ�3�v���]9q�چ+B讍�ť�ު<$��PI�N�C��Y=�<����Օl����S��T��{F���b��=6�#OCTb����`��<;��ڔ�m�7n������(�j ,gQ���5��r�書�I�{�꯫��dW6sa�i��]�����'E�T#6�<%�J��`廓�(���zL���ady��o8�]�hk6��+u�',Rʱ_������{)�S�����qp����iϛ�.�o*|�����*�Q��l��]�V�!��fWޱI��v���0p���_&�T�rx-�j�Q{�k��LǬ9���F4�$nPܷw��D{X���ڿV���ϧJ�f���o�1�<)��,.�͛
&\y���=�7�A�?q���:���{�Ż;k�+Z�g�En��k'��7/p�Nl����.�Ÿl��>��^t�����و]��^+#�C��|�5{��^�I�^����Y������fۗo_#���}�g���Of���4!�����;)-�^��"=��g�:8�{/Q�ʾ�Dne@�;{�Evl*�W�g�j�/�����(�l�.6�;S|*������3����z�8�t�M3ZW��(ތ�|Nm@�xU*>n������.7�MOY���η;m��U3z%�i��~�ؙ�K���7Z�]T���&���q�:��Q�â��,��zi������Ӯ�PvMڴ=θO,|=Ჵ�fC_���
׊)F}�⊑��a������B{���y��Z�ƥ�I�C�&Y�t�\u���lA]���a�kC�;���Qוo���]��ro��l�ٻ'M]�t��k;f\Q_d�u�k�Δr��N��vs{E>n<��B�r.�Um������Ecr:b����e\G��sD <�QۮW��}1�*ܐ�Dý��^"]����JAp���5�'�L̘�+\�M�;���ܦ��,i��~;�7�<V��~U���5�_��sћ%�߳���m�c�����'�{۽�+����<�g��W�7T�/_yK���n7�{+}�m�̳n��|ߏe��S�6*�}�YK���Bz��`Q����*��]-P�Y�~02�۷wc$ӎ�w�SX�ğG�d&���9z�s��"�!0x�����+Ѽ'��]:W.�'C������mc�@!K�|��EΉlyT1��	�|x%n����$��<N�D���G�y�͞��i=�1 ~��j�/f����ف_W��swx�F�!�1p�4`�)��;�_q�W��A6n'n�)m]��*�p�}��wk%�̤����4�uN��N V~�o-�t���v�]1�׈�_�șW�Ӷ�թ�5o��+Ϸ�&�WZ���xfQ�>r���f�'l-��y}�xZ
�ciO=,�^J��=1T)��aJ�:8q#��.�pjEK���;�,�&V����7�ƶ9�҄nw������qj�r����2]�a{ΈǼ�VZE�D&R ����Ӥ�YL,�%[�n���Lѕ7z"�6��>F:Ъ�s[T��v���1d�塙OI���(����7؛Ήt����2���b*iH��"��,yN� ٺ�-�a��;��w�lv�nD�M�z]����ם��'�0�Rw�e�!�ɿ]�Gn�7���/3V�������NX�������k�M�yn��!�����D�T�������_���'�s���1ty~ʯ���n��E���#󂉖�վ���;ILn�v�b�5��6�i�&�E9��W{_b�D�hU��/�vAU���c�{;n���%؈뾌���B=D4�7yܭ"Vs3�w��"����յ��^d���.��O�y���,j�_����O���Ä4��ʂt6q�ё1���n�H�ۍ��y�|%����}e�y��0(.����{���w뗕c!�R��n�&"���F����ul�w�f��;s�GA@94��b{�v��r��W$�a�����.��#�S�� =�
�!@j����һM�j�>ͫX_��?H�^V�H���.�J�}|�U:�dp��0L}SK-�[��Ns�ps,��q���vv0:��jP�>�c7���Ց��_>�S� c���j��]j�I]x���o	 X�]k%�^�6ی�ˌQ=������:����a�űH�DwnJ��L�h�t�y��o��j�9�5X�Ό��1�	�rm��L��4`÷2��*~γ2a4�u���s���a�ӎS�����Nx.��|觑=�s�!���0D�J���Bޟ��fݧ�	��<o��o�bߕmg�0��ٛ�(��;��.oK���Q�"���R1�a)��Nڍn�u���M����vڨ�>;�hz���Q�,�r��j�a��³:��<�7c�i�=���j�/���QT۽�As�9�uO��t�j^�ֻ���'��~������8{+;׍^�ᔍ�/M�zh����FX��s�m@�#�~ܗ��yP��v�)�1�F��7�I��3�7�">�ב�N��'���D=�h�F�#���Ỏ�<�]��یë��]~i����|Wg��	)�(4�!%�,�����Y�nv̠|/&���XQ�>R�u��H�ɾ����z=i�p�W0�^�5�6
'�Li�R\{�={x�~�z.�&�}�����fydd{x�n^�w�7�*_��OJ<�xF{E�X����T��ڽLJ�:��Em[�7�Ǎ�y�����Oc�;N��w����4��69�R�sZj��V��l�wh8�E��}Kwܺa1�#�f~��M�_������rEI6v����ZV/ͼ��Ϫ�c�Ri�E@���RC��(�P�+�!ڙ5U��c��%c[��H��;*P�r�+�[״�64L����<�ŗ�DQf����8��堰eew7ֳ�&5�?���i������v�L����0u~��a�Uv�^ߤ~C�ͧ�>�_�|�Ѹ7T֧����&���;�\���tx9�=�t,D��š��d~��e��� �̰���F^m��	A�u�)"{���]؅�a�S�����	��q��I��C��AC����e��#<u�{�K�����w�#n�!�(�Qdy}��]2�<��>dU�Y�$�a��t7v��Q�O4p�KC_�9<y�Q&\Ւ��M��}L��ϼ�����=zw-�.ڵ���&3�������;+0��ԓ1Pg���b����Jp�]0i^�%�tEe��`zmQ!��ga?9�Q4]�:cio?%b�ν�.�']p�ء��w�{S�>��;3D������?�;�q^��g�0A_B���>���
Vo�<o�
�.�l.�q��H�^v9
�a[��ڬ�=���"8;G��u\z4^�����_���y�|;r�oԄck�v�=�r�3�\rLۋ�xH��w�
n�@����[������q�q纣��7hp�Zr�6E�m<t����jT}�T�ׯ��U�vGv:M0;��5�[:�Az���Wf��i��)�h�D��dU�T{}��n^��Jl��੼�����:ܒ4rS���HN�����FlVV��G��J;�][�V�y}�m�L��Y��;��/{§b�~�-���{=��N��.\[�$�X���T�Ε�wvA�q�dm��vLܱ��A3�-r�*�w�WCm�^�Wѽ���}�UM�}��W|�<�;�u�}~��3��,�H�(���#�Q����׆;
���+_~8�D�����a�1<��1��t0����~�4�^[�٢�7���;�q��ݦ��u�*�p�R}l��@���7��W�~��iﻲ*�D����۷(?W^qy3��/�)b�^C�3��K��G�f���:��
v����a�^�������m�G���β�PnB&�C[Q@��'S�V���y6(��-��L��"S8��K��V�8��ơ2��T�{��b�Y���2y*^1�U�k��EYC�o!<+5�p����&s���V,��'��(���XJ�)��}��x���{�9��`�p}mv��HD=:b&�M��~]�&�U�b��L�L�/T�pcw�u��Y
EH�(�#C�3�e\[�����ם���f��v�g�������>�5/����͓�7��vB�(T2���\~���X�ʏw���+F���$��"yN�]IӚ�j=Ov��� _v�M��W����DI�������\�[6o7X��ݳ�`Y�N}p5���y����*V-;ToE��h�͒V�²�Z.WJDv��&�d��Ņ����U�T�h�ô:�cw�=d�j�*�5�u��ۈ�B�=L�&��B�ۦM�H����I���p�Z��T��������eW�^���r7����	�=o/���P��s�.���D{�����zy�>�]w7{֧dz�j9F5�Ե�U��Ю��ѿ�^
j��2�Op���K�h}�����.�n<�yŨ��p�j��3�B����UR�E@�|��Ǧ�p���%�`�z�B5�C����V.�)[^�v}�J���s*3���i�.�*xB(�,cE�(���.�M�t��5��pC�j��j����4fQ[�ĺ՝<�a��ܯ0��vO��{�u���W��Nc�Svt��\V��W�	�u�2S��O�v|����Jwa���!���N`�;I.��w�����.jr�����Xs��v:Td\O��ޅ�F�7���/O�g��	�@b��@�(GG|�b�Z�t��G�0��=�<t��pkݳ���S����^�����u�cj׮Q}�t0m�ܡ���|˝�`x^�]�7W+)n�p]��O�[&�t�[+��Ϋ�f��{W���n�gi�䕞�mq"�����:�6>�5��06�.������ܱ���P��ق�.�:��9�o]d�8*4�S̢ڜ�E'K���b�a����d��������+>�-��>��<�J��;�48:�:��(U<�Rg0Dz6�+��)&�C�N��A�M�	{�6��U�d�C�c��d�w���.HN{Fv͚z�LٳPg�f���?9jT6p�Rۡ^>�#ѹ��9���%{����r�o}�W��y٘���<�y�OZ:��h�
�]Ջ�^�3�9�R�yh�|��.�؇7(o�w����R��럎��Č��(�*�vR��H=0~>��[�E���sW��h��5�m��+X5UJ��=#��`�u�+��^|b�Na�C�Y�w���/��PF͒�F�p����~wⳈe��:�������I�sT��D��n���zm(��.st$k1���0�=��sTמ�V��.��o_=��v�C�N}%�НɎ���Z�@}� X0��Q�j�{)��<�v�/��r�7
�]���7���,M�:��_��6��~m��6u�����������e��wa���S���O��w(ч�B�f�մE4k�)�L�!ۣl[w�|z^_%boQl�մ):9����j
r!�M�nc�p��!�Pv�r�2�L�0h����/1X��M��枢�~����>�7��N��n���]`�,wS���qsyi��=�����~��ͷݸVr΋�t�u^�����^^��BpY֬3���|�N��xY
�~�)7��g�/1�hsN�N�9�=�Z>H~w��~�ZT'}�����Ϻ�M�8�<��͋tvп��r%�ڤ*�j�����ɹX�Ӌ�P�F��[���j����:=1X�
+�z��ݮ��zχ�T{.���7}^�������~�������Yr�֦��z9PJ�~��v�-e�:�.
�=�;n�߷[�d*�;Eɭ������b����x�3��o���\���݌�X=�X:�Gv���s_���8�R���Ky]�����
3n���U���{t�YC:��ծ�p6l�1�<W�nEe��
q�g����	9ŏ	�� �I����2�X�]a��k��X�]s�u�؝�+�2pê�O�G����xnS��:n^��_zތsdڜ��י��12;�>����Tx9U��p�o�~����/7�]�*v��N�Z���22�\�5^��<#1��=>�Ur]�r�
2똸|�C0�j���7��W�e\�n:�(L�6�k0T���&�Kn�<���9Ȯ�z�[�8���z�*W	�p�K���-gV�&�@��V��i�{����Gs�v7��fS���d�5-���u�ά۾�\��S%�ԧ*t�5;�P���м%�&���S�� 0���t��\��*��,¯�;c��2oa�b�Q��|��Ӿɰ�VAi�����Á0�oܪ'�,���>�\D�t`] %3��tb��;��4���n��P*-5:l��O�N[���υP7p6�c��BBA�bp�\�,ǐ��f=t���*��K���ƈ7�읟Tט���rz��Ү�_�:��VF?yU��Jw*��f�g�w���KE��{�jo�Y�C���`1�s#+i�5U科cg��p�z�����/�	!�;6�w	���:�1�x+ �̚�*7T1��f'[���Ngv�;���&���e0�q#</����3#�:���.����N*#,�н]w<k�ѵ7\Vt����c�L_vWnW�%YHV_��!n��������ޫ[�ՒYk�-.��Vҥ�J�R���>�ϼQC��,R��a��RУi����v�K��u�I���e�t;�E�l�#�d>�y)���!{��,��q�GS_|���]�*�Kv�T�>��w �`��_���>j���N��Ɩ�$fd.c\Ϗ�S�Ϟ��We���u��[��e˽<2%\�S|kO8�2�x�yq	�ԅk�-e�p;�V_%���bo�Ԏ�*�;�4`��T{2�(��¦re�*]�G1�}���嵑q�^��̥R�Rz)����/`�;&�EE*rT��zm��VK4�]t�*2%�lԗXg�*L��e�8mm0���ڃ	��ܚ�����j5��f����hJr�Ȝ�L�v K)K�NʹɌ��u�����u���]ΝǙ9�|H.s����o_�����'��f5�Y�ݖ!4�J���˻Jt$���gJ2qW��Sl(�G��7�S��_$H�Wk�osF����`l���w�y~8�w��ϒ�V�3��Y�����4�k��/^�����c�T��7)�A�0f��/�71 |�����޽BQ��Y��4��B=����;�k��~�}�޹@�@��HÓ[�3fb����oE���B�L�G%Q�9wt� �XH�_.�7s�k��Թ:�4a��*�oZ���c��oﾴ�1�>��a�@��w�8cE��,��ֹ��#�m��	��(P��|��6^ūa̓�T�K\��-���4�c�U��b���Nӿ߫�������I�67��=~����>d
�=����u�8�������~2�VI6�,�9^{b���W���Zqru����FR�ӢN{Zpª��;g�
�1��u��JX��WB�p����l��+�S�֎�"i�����W5��}�}�U*p�� 2�j����,������U.���\5�9t��Ƅ�X�g8�[�<1�a�mnƀ��W��kc�Bd��"�����V��kn�V�=�?e�U���m�� ��`&��h�Te�4�d��S�I0�$�	h�m6�7L��w.��/Fw0�ЏgU�]L��{*�-sq��$'�ٴ���[mEA��̛�7l��ߣꑶ��[��524b�X�����7��/�;Fɸ�/xg�%I��=�}��1���5�o���|J=T��F�/]�&yPf�8Z�{0�'����^�z�IZ�V�.���U���mK�5�;NA�M�Qk��X��=�iC�嬝���F�J�vM�ֹ��V݊V��Q��]��g/c��g)(��������ÊQ����(��M�E�jք��P0kU�[R9@, <;�e^դ��|W�o8"y��u&�wͷ�sTV(Rl��gnh+Vpse���b�"��e[n���h��En5ȆָѰp459���k�������	4�e��Ec�z3m��3H�a�Y�J2$�To�����#6)��� k~�����"ĺ�ם�c�Nj`�+����T{4!�Z���ˇ�*��H0c+Kڙ����L�j��Me�3W~؆wX���V�3e��[�A��h�4�@+-�����R���Qe���N(�{n�h�Q�!VZW�_��)is�� 00v�M^�o��W'w(Wea2��CV�� �;��5�4O]<J�lZF���5}2��Rىv�%wJ��V�t��&U�X�Z�@T}�������_o@v���IρM��.�o!أ��)�ʊi%�������6��P�C@�7�*š�*B��?�@��%��
�N��b�C�+&�^8R�z0f+(F�]�u�����%�q�6䐧(���҃�����s�K�Ӕ%�� R�,�[&D�(���T5��X�����S�Ly�0tFTYXN??gg��wl<Nҵ??E���V1p�2y������׌n�e<��upg�ɀ�.��w/>7�����[�lQ��ȼBD+j	�z�+�qAt�*��;�m��]tH�w���>����e���m��m�KX����zL�S�����M}�J�7ۓ�ތq ö#�=l{��S'3�G�tE��=C+��;CW��b#��_y=ھg�VK�����:��FG��1Ae9��',ﳡS��lQ��Q�'r~�o%eWb�G�1�-��UN��YP�&й��n��j��Bt���
><z색�S���쯲��7���],��[÷�QMT2��h��oy����R�+�<��|�=x"|g��6�;��R�QU�/0}V�4�R�O�v�:U�iG)�ÅE���"N Ө���闗��L���D��frg���L {S����N%�h�ǲ����YU�v�5�U�����de*�of�BP�<]b��ϰ��@)��v[Ω.[/L���e��7����B��K��tbm��˴Ҏ�Q �mY�9v�29��u��� �\"�e��J��U��{EOu*���	.C��En�b���a��&�]����0�pb��7&+s�p���ЯIy;^����qX}`׀����Jr��Ҧ�	��w�&��v��̺���_�>
�����EF%��w	o�=C9Qӹ�,f�o+1YѵwO�4�z�U!�.(��ʉT�Q�
!���`����w|�۟�$��NƼ_Sg��B��*~���s ��c:�lR�<��Xp�A���蛲��$Te��V6�ϔJpv{7�6b@�a���aAԤBoiG��z�z?�����g�]T��<���ۨH�*�N�>����2��i��.�YB���{���{���I�ϼ��8�Jo����������m�m�e���j�K�WHz�%�.��{j�4��f�k�9C�Laif����Y�q:6�t�y�C��E���Ε��������rPa�!�:��T�Zx�v���L���u:��U��~O���9{�����Q�(�����=�zX�8��"��?Cu�2��Ӕ�.��S�_�L:v`E;��RR�����[�|�Fˮ�E�־�{���Vj����;N�Γ]|_Y�{�.'�z�G$�Y]�wA����f��oR�O�ۗo�D�a�¡:\ƶ&��N��řU��[�V��f�S�ILE$գ-��ٝH�c],^��{هx��2!����^u�����NOX�C�~6�A��=gi5VZ�̝hO}vh��3�J�_1�>T�wP��K�t����gx"�W,5>��sߥ���� ���6��˃ƒwh�(kj�@�]�Q��y���Z�埌�T�����}O��Z����Vz�J��U.6�%m��灭5!�{��m���<Mv�������ڛ����\2s��������ْ^ep�p(葾iT~~AM%�/�ˢ�]��[�"C���kg�٪�nB6s;�~���D�e�`H"���Q�{��!'�<�w�ʹ���Sj�X�f�����]L
^3��(���71�6��b��+����/�A�꺲�:�`�����c�M�]� �a}�kL�e�aI��mkY�gr}��;h�!F�w���YP⣒����Q؋9͸��~�袆���G�\��;W��Y��]�O%�EɃVϦ�ع�q���z��]'ŨRw�鯮~�6��5�ҽ����C���ȣ����!wK�x~WH��������P���(���xRQ�r����u�Wo��+oKǔgt��Q	(˨*rx7�8'1�R��)~:�eԧP<Ьc;��Y�5y�S�7F�ۥj��۠�T�r�u(�\����p
=����j0�7Fu8,d�	B�{��j�h��N]w(*�.��Y�S�xG���_��3�O�|cD�bPo�%4ÈT�@�ӆȮ��}gH�t�`T�ρ�f{׾��a޷�� ��ߔ�L>�n��b���!���YR|���ǵ�|c�`5��q<o۷�y��1�P��v]�����Z��L�<�,ǅfP���'�Cɧ��&�W���Wuz���ڐ7O>l,��N!ݩu��4��:g.ֿ_!L�"�M?�;+��;U�;�>���W^d{��5	+�.�v�U���v���ahU=lZ��L8���W`�2�v���:�Bs��C�������T���&D�,�ւ��9q+���p�Xid)�wê�\7#º�x�!տ}Ն|*��Z��{m�	���l��>�*�+��v4>��j3=k߯1��{A�^�:C�n�%mU<u4�>��>}�6*�g,C=oh�4�R*���X���m�hi�cZ�f�4�(�;��v���
X�NMwe�����*��+�y��|�p?�q^߁aE����5�SM��N�����p�G�c��{���6�nc3w�+w\�����0�P��PZn�R�q��W\/PP�x�7f�KY�)�{�D���2�l&��Y��wqUk��d�����ՂZ�E%�Ź�9،�3�HҮ�Z���B2�1��/���7VՕ5��qu�=����ؓ_Sl�޺vK�>�m#,�֩x�Q$�-'c$g�lDR�NZ��q����{����?m�g����l��+���nz����B�@�
�-���e(>�h��\K\��55�{�@�&��u�k*��h��+��	V��_=�Hկ�	ϱ�Kج[��o�ϵ宜���si�]�P\x���*难�����S���I�u��:cU�-'�Z��۵y[�̯��Љ�%������jwX�7j>�F.��k�
���A/����?
��o?Ve=�p�{(1p��A��V&��cǘ�OTW�j*�ݲ��1җ��4�ܘ����.ӝ��W�4�U9�=�no6V��IG��߀�X���_��'EyL�8߻�;)� ����hV/X-u��5.�=kG���30�)^��%�m���7�sR�Wzc������������5��~͋5I2�6�����ӻ�U�)���4>O�~���#y��fyg�CQּCߨ�e�)�Q�xw�|f_�g�N'X��nAL0�V�Tqȩe�dFޤ��K���(�4$����D��y=ڼ��깫=ٗr��X.6$!�1�5f�&�͉�����<����e�Csgi�Gԇ`&x�V:��`�&�r���MN��|K��X��l�����υt�+^t�-I�C�أ��m��=o�[����>��k��϶�-eub>��_P�}��]�osA_�e�Վ�B�z����H_�
�%�޿ѭA#47,��;^�S=�k���!^`��묽�"��z]
Y��͝t�C������/�W��U'���Y��ǥy=���*ᮈ�5>/»0�l�Zث�fj����ܯ��vv:@,��!u�;��c_���ٳ���mx&����3�p�<)���]1�#r�}r�Q8 �ӡ_��ߧ9���5���v��Sn���J���*�񊳹p�j��עv�د��K�}'��8Я@�a����~�e�Xٿ[�����4b5������\y��w��<:��9	~ƺ��|ʗB0Ck�]��}:�S=}iҖ��*����ͼ��Y��F�NH_A���rB�~�E�XdߦS�23d笾
5���3S��T?#��	�B�߰ٱH�7f��L�:^V/��m�4��������Cg-V6��6�uǝ/���*�{?f���u>8(nK*�ؐ�n}��b�#�\n��6��A�屠���7zʭœ��M�]zk[)�7Y�R���.]G�l�?I(���G��Q���J�<yS����c[T�|���W�/U�v��M���N�=����lIφT�7���
���j�=5j�-�{�����%K�Ʀ��ÈgE���V�������H����&����/7y8�'�5t�K����D̵u����7,��W��E{ˆ��<�m��~ʥ#��6�"�h�3/MΈ��ۼUIw�|������3Ųw���E_�io��e���:o�:�0NA�аm��^�����>轡�������U�к�]y��b��8<;�N�݇T���*O�|�ç�Ɋ~�XQGug19{�:o�_	{wg�n=-��D����R��_��x������-E?u=���얫�j����,f�.h�X����ߜ3���e��=�+�Ei���+�C�u�d�\�O�ǈ3�in�l��j݊�L��)`���	v+.@��Δ}g.}�2$���=��]�y�%�����������w�b�I���������럴N>5**������4n�cG�:�;glɼ"��>��H�j�G�~>�v��hg��4�M��B'I��l���F��"������}M�[���"��O�<m�[����:���2=��\*�wjFVaS��dsyI1�^�.�7��u��I�7;�rE�;_���f&9��FZ+7WXRj.�##�[ǐAҩ��I��i6Mi�⦈л2�`��`��%���\�J���a�j����	���^ig_f}R��7/�l�e�0YhZ˻<X��B�J�w>����Ej�
�'qt�u�GcU?+yh�f9q����_I����48��C�_�ѺG���6����U�z}A p׭�]u�Ƈt�o�*����*S�1��;]7�F�-�j(}�1��U��I7�>����Դ�{��F���:v+Wå�����ݕ'}^�Wp��qV��MXQY%N(i��J�@��ľ���v�W=j��<�Υ��Y��9�o=8�Z)Q��-�j��ק�t��B(F"���8]�B�0=+OnH�3``�����j	��N��R���!z�r�hW��	�(�����7�
�\���v�Q^�g����VhL�;��q1~���B�r���wX�e��P��W�*2�4�f�`����]_�D���Nd6�(�VIuV�P
{���K���:���u�p�uhXfu��.��C�-�~iz릙ۼ�ho޶9�f����.\#w������a_Ec=���n\
��)�*��0��7̄H��TF�i_�[�/e����L;ț^'㸖7Z�T�{��>w�0��PQ��*�0ge���7��S۬�����h\�
���=���)5ct3�f�g=N���� �cUb�2�e���0K�(1�A���0x�)�&Q��X)u<C3��N��r��k"�(MJ�� �d��F��2��k.�:��q��s�7˱��J�F�O��Gf7�%��G�Dn�8�:or��uvjR�k���u�`�c���ȩqj�zoB�;�\�A�5����U�z��co1�u��3.+v��+�K�,ٞ�tC�W����<1���9VL��]�oW�8!�>Q֪�����</�1`��_�4�zۙ^��hI��Ѧ�?����������#s�<���6��&�b!p�M`R5xY��X��Y4�&�X��1r���i]�܌���*k��lW��˳�Y�ģ�X�$���˔'�S��6^��m�U�.?�v�6��C�nŉ�Ξ��O�<��%"+C�6Dr����y>S��NM{Ef��^6w����1ʚU�����U"��Zb��vl�lF�K��9�k�������������J� 5�y����7W��Ct��[�Y����?�r����P �Ggۃ5�?�Κɋ֦��{g�w������������(�z�f]�S1s��eT.��Y�|�
��'T�Ǔ���i���2K�kn[��?��7L��],#��!o��].ї)�ۉ��,=�K��A��Vg+ݱ8|zU#+��B�l��1�Y��)��"N�fΣ���d��k6������
�U�1�9�xKP��y]�=.ktk�^�1o��HP�3��D-[��$%<�겼p�ƺ�Y���wn)	��Nɽ!������"y����-�Nh}Cww�$d��� ���]�³����#o�x\�;ށ1ݎ�𫺬͹ڢ���:�ڣljX9S�a�>Y�7V<I�W�_��oٴV�TK��j���#B/��7�Om!���w|���?nk���D��\��ՑTbj�]��/k�>�u��6�oB��pU��JY�v~�Le06�0��!\S>/r��e��"�JC��k��=�g��Z�B��������Sy]'l,�׭P�5�3�֞kk�3x����繦©.��pc�t�'/��YYK�a�����ђ��Q�t�P�%���}�9��yG�^�ƺ=^��0(���tĿ40���1��+.K�����$��z��M�+e Dp�=��4�Cm�4���>�_`��tQ�5s|���yMQ����bߨ�B�~���Հ:�Z��Ǫ���i��Jg����ΚkkG�{1u�3��T�����l��;�p�eZC�b�'��<�N�W�b6.����<����܃�����eQ�ћ�u�)��z�.LWkͳ�/ڑ�uՎT�<�-��o3\͖�tMt<Z��z��%rɇI2^�S�1ui�٘�1���v�m�N�a8��=�W��sy$�4y�z��St��㝓  ��M��L<-g-{m�Ά"��5Ks�s؄�q���@^��E��׽��iҴ�T&���ּz�.���F�A}�h}�2��v^����z6�#4��;�ͭ��@Q�(فKtjYշ�S�i>�j�'�/f�"�Uᯡr<5mJ�me`��*W�ux�ckz��&��Dڽhlrc��v��P�V��6�����`��^��X:~�]��霑���T�3�lp�iv����;��/�՛}�f��b�f.�]u��k!+W(+]+�5��&b۫锻Pvu�͙Wc��yW��E�RTU��e�Y�0��T6*k��k�3�"�5#�<�v�2#b9�y��[FP�rxw��s��&��ʽ�v�,[{�;\�+�+l]iV��T�V�dÕ�w�p����B��$ΰNL��bљRP��d$`�kpJ�z�ٸfM�Mh��ȭh�1>ɇ9��*�51��b\%��U�&�]�v�-�a�r�r�Vf��1oh��ipΒ<Ū�C��f _;���mwcJ[]Ӵ`���B�>�RC?.��s��z��U�hl�|W�oN���|�h����3�Ď�V��UG:�v ��w@��gr���}�d����n�.?�1\A'�acg.����*�H=��C�J����z볹k|M����"�K �`�]��\��rP:n�}G��L֛����I�](�6l�R��Ƥ;y}Pt���I/8�Y�axE���N�	��j�]�.5!_��.�hK<q�0�`̊����M2�e:�z�j��w���c!Hni�9�Mq�v�B�zV<N�,�	�0�r��Z*ȫ��wS��K�sQ���nq�[��N�{�u�Ck!޽X�N���qW �u�Y%
`�x�{v���Rغ�j�N��s�� �-Yl�z�#m��H�(r䨋%o��lÃN�\tq��=��E�R.��n��ǙJ�k��û��݇VSn�i
崠�K��{Y�D���2��ɨS������\�W:�:�$F�j苰^f�����x���C �당S���˴.v��o�Eb�"I;�8(6<��Q�/,^*Q�$��v���U� G;L"�FP�v�����"�����Yt5�deq�ɱ���]���r�u���R��PXE����[}*��іi����R(z�n�rٓ�_ ���"�8Y:�J��$h7�8���&[� �ݍ�9�wG4�������c_�����V���m��ё�sGSw�$le_*g�sU��Z�J��.�Zw)A�ciN�3B�4׍�������6�c��Hh���=��L�H=�1���mi�9|����'����|C��Fz&��uM�5C"��ڨ���=�JΨ���
��W���y4N+J�:hL勆=�z<m�{�{���DJJkHpb�!K\<m�D�(��_�⢑���VP�������g���e�"�]�N"���)�\,ؼ}�x:8���c��3Ňy,xd�H�X�Y�ep�F�kv���k�ʆ}���;G@��8��s�W�`9a�j�֝�l�h}���Ho~(���`�'.`x]�8GEy���/u��W^�G�ڢ�[71��?�%��<��ܮY��kd<+cς��N�|��[��G�[��v�K���}+��4���ߌd@p��(ϕK�r���a���dNʿ�o'�$��b��	�[�K7��C�4�/[��s�ǳ����J�u���Q��gF�����[�S{�D��"r����h,�w�2��٭	Fg
QU�=���0#ō�B��b"�eA�n}=N�I��Z=b��C�
�U[f�Ѿ��qVH�ǅ��-c�.����G[�k'V�%���OMq�ԗ�Jd�m:��˨	�[:��u�7哟7�Ӯ�SX;�&#.`?
�%��j>ٖ�(�鿦�cݰ��u�Ǫ�¥t��xf��o7�
�T�鈛
H���Lp�R�+w�.9��s�#�q�8���H�a�[s:KY�����g�Uԩ�-iu9��{�1���3r��q�8� (��(������dO ��9�O�lw�
ne��L�����Y��T�ϣ�5b�v�;�k�Hnqg�o>8�t7ޝ�ʯ~�%�a>^w�*,X��������H���Cך�u [�y��}��ۼ���K�����:��x�}�LTH�X���|��dp�~���V��6K��K�����_�����`��L���,R�������Q�=�#՞���/Hw=���iG^����rPq��<�޵����DЉ��(�v��d=�Sd*
�̟1�u#Ǒ�����ϧ᪱O�6{��kᩏ�c�ʕ��S��~}���@��mt:&/;�E�����E�V=�U
z�	�2oM����t�f.���ح�޵|y"ATL4�`��ӊH�u���x�NGr��t����kX�[�iJJ
�OaV�J�Tz4Wm�A� �֑�ӅY;�ޚ�N�e\�tu�������^F������D(��Q���`]�Xp��������$����{5k����Wދ�<	I浽�iƍ�v�$Ga0��u��|*�S���k�;X�X�?>O�	�YK�ś߉ی_*2���=��5qvM���j.:2F�u㋡�o�aN �ݚ�x����>�����jژ�����̱�viEW���X�? V����b}����w�$&��v
	B�}[���G=~�V�S�k;����y8��:�]�n���P�n^U���B�)e#���(4�N�es�!�w�g�6��pM���������X�	�w�.\N~��E���Ѷ,���̘1��s{��\�Íi����&ǔ9pb��[b��r������&B�H;>�����GQ�Ź@t�7�U�pk�Ue�霼����Q	�<�%CF%m-�̻��֚Ҧ��}3�H�]Y��I�_���k�ڄtBR�����z�E��r��dVm���t�)&y�[�gr�yBku��
; ��Q�:e_I��dcjq�,����lF��&�����.�e�[���l��ڮ5k�'���uev��5���r1\��8-�p"�}��nH�|�%�L;�.�w'k6Ll�J���B�fb��c�*�zkqwW[��v>�Ŷ��8V��'�e�����u�8t^�JWѯ���E�~}B��A��<���1�]��;]�!d���ݟv���qk/�BK��`�rK�*���=���^xY�믣���Y�/�hX6ݚn�E�G�y:�1�}��/x��{ŷ�� �'�y�;OBa����w�7�+�����Q��.����
��g�=)����rԂ�7�{y��m^z9�?k����᪢�Y=�������uu�Y���9}�����p�T��e�xs{qƚ���1�F��舩��W�L7�Ԍu��4�W,m��Ί�z�����#�����s�H�	zC���% �nºDX��-7W��+Ⱦ�1�:�"}�r�M�t�p�v�\���t�g�U�=��{k�'+1�����kR�W;��{PQ���F*zb�:�:����2�IJwZY:�6�bB�H�8{	����l_�v�|@x��d���x��7/s���\��Gm3/�f;r�����w�1�z0�C �薘	u�@�bu��W]ɑ�h��l+=z}��Hױ��O˭�����+D�n8_��Z_��Ch?Ս���YQr����[޵2��Vj�ժ�-nϮӎz�C��݆�Q��U��n�w`~�m�"r�s5�˞��y��g�6zF�ݵ:E����?tcz�ר�yj����"��Hz��S6V�3BE��+s���<:��Ұۼ��L����6z�,�|:E�9�h�I`�{89]et�ե���-�>��	j���&��A��LH�s�q0t:����f���~���F�DT��-�j��;"��r��[��/f}h�b�ҧ��7������o��X̲�D�7}�QG!�(cp`�7.�wx·>�3=�5�3�*X�^@ܴ{�n��uT���m����M�2�����<&���9�d�DC䔎l�m3 ����t]>��'Wmk
^VР�b��s���\TPt�5s���w�\�{�v��c�ץV��̚��FT�>�t���9�o�Q��-/�DKi��[�'aG[�\���� �X�*znYꚃI�K�t��߼
�̞�!z�~������n_��u&>�]�B��%E��\ԁ��sfԗ(G�� z/q5�̕S����}�����t6\��{�&��_���e�O2>�d2�Wj�z_f=~:��p�1�9.Y0dM���{u�T��c*�f��9I隆N�>϶��qȨ{���Îx�X��8}mb��}{ޮ�XQ�b��U��lh��U����]`x�Z�m�P
�.�,|of�6�B��+58~=�T���;�K����=skjL�L��C�s��y���������c��߲�zŊ���<{9�ĝ�E��n�cGm����Wz�����ʟ�]�[�����k��ӅD���=Ζf�_���������k�����1���=�7�tr���:�HI��vB��W�c�G�>����9CW}�g{�����~���@�_su� [cSb����&U6x��B*�<��R�AWe��7�WVs/
l�È��]�� �`�t^��Z�$��)�I*���#[�32Yv�u����� �,�o���H�/���f�Y	�����Ϥ�ZUgoW!�᣷����\��Z������%K)�Jr���A����m9�,�F�s�1+�=��|ໜ"����}x~�}�v?��e�p��.��nEo�ܷ3���VW�n�'�?F湄(�2\����M�/&ƕ	k�d�|Z��T�ޫ���+���2���ck˷��Ȇ�(�	������ޡ�b�1m\x�Npw�=������"n��t��X쵦63v�U�:��ʏ�]�̮���f�z��6�uy���:�'y�dx1��5stV<�m�?Ю��J�o���Yy�L�_���xa-�'U��G+�k@�������pbu��	n;0\G�;/�[|<������?�叢S3��Y��{��ǃ�y�������܅�����K�$�*�vӺ�Aŕ�r�\�φX7��zk{&�b�żZ�B�X��oγ}��$�F}!�|߲���3�o�h��v�4{v����S��35c	��츷���Ի�:V��aYS��6�3��������8�^JCQ枤�{#��NK�5�²j֡�3j��H5���J����<V�Ќ��[�µ�;޼՝-R�'j�1d��r�j����긑ӼiWguH�wUe"N��z�]�x�:ۣg
L��!�������j�ev=�4��Y{�0]I�}�j.��h��wħ/}�{�F1q����",��W1N(����CI��8���k���y�V�r>��������5��m��i��%د��z3�������>�B���3�4=�g>[s��Nn�����K��1�ꑎ�Dyz3�K=�0��.���0���e
�3V����}�uR���G?{���M{8��dȺ�L����zZ�XU
.�AW#���t��,`�v����XI!���F�>��q�<i"c�|��Uw+�]��4�DI�3�\U�譺N+�ۖ.�GM���_����������.�y�k�Tn����:���)O�����d5ո���Ew��ݫ���/�{��<�c9����V8� X������a�d�w��Om�{Y]���R�I��/c�d������}�J��(57��=n#�;CYTp&���w��!��e����4��ܬ�pZf��֤��)}��\�r�����=�+w�������&ӛ�wq��5�^�_�u۵Ϻ���>�\�}��|�:�O�ײve�������Q~+D}C�:'�v���:xf����|��н<[��&NK�~��Ϣ����B�*����n�>�r1o?������'�.��{7n4X�}�x����݋�=��(O��G��k���1�x��@Q�'n�_��m1�׽Ǜt�F�y$[o6jn�|�w�x��ݮ�*w���Y���҇0�i����f��4i���!�ל�ٻ5篟�M��P��3^-��=��0�M\�o�{�2,OTbx��P[�({1�;7�j���85�C�5is\Y�Y���g���i�_���Z���g(���{:�8����l�o�N\o��X�J!v�~���f/jke�HwkqyTz�v���D�QW[SK8n���Y�M]�n��9VO8��l�_B��%aL�[����A�v��e-JÚ���^�ǘB������)�C��7�t�����ۺC,�o^�j�X^�g+F7���M�W��@s#"*�}��_!��a#��}������������TyO���37n$�t�J8��o��0y}��rjC:�^�}]Fq��,��L5Z��e�U����J�j��{$���~�C͜��*q��*o��^��	�K����ڧߡ��άj�Q7f�:9��ἋF���,n�+$�8L��1Z����,���=�V�_��[�iz8������˦�doʳ�6gW����Wi%���_A��Ov(�D�C)�t���U<�y�r�_����J4/�٘��?�Ϻ2�稵�/���cx����n��j�$J3F۸
;�����a�@t�{�B8&���_�!�/wU�٣���7������ͭ�Wǎ�w���"�J%�Քs���M�l���[C�'l�Or�f��\��5y俏T��=�to�ښ~��/��v�AY�d���q��i��ʓ��N�'�+�ڥ�R��o���jr��@àE���ʼK6��N?�G�}���f���vOwr�[e�D4-�Q�Ѭe�j��f[��'bT�=;�\�K������ol/o�������j��[�2�罜��iP�d,�)op�N�a��θ^�.�����5����t�
�!���rg�	������i�ܶ�[:s��#]�W7٦��''�R�ҷk���u�1��|^rݡ4aۉA �Otbl��71��M^�ɡ�ͧ�o������m�`�b�������J���W+��̆�9<�\�@?,���x�U�Y�]���)r��]�c��%��dP���c>�}W��iy:Є��QN:���Tƛ+�+�
�*j۔2�D�O��ռ+��Z��	�b-�U1Q�ʺ�҈Ɲ�E���$s޵��%yk"��Aٹ�r�۫������k��h�jnp��k	�+K��ҵ<�����q�d����m�v��S�s��o
2���wyݚ�FR�Cy�7���J�Bgm����Z�i>������v�J��n��w]�]{L�Qk�d�����P��VT���ݲ>��]�c
�<��[���K��4;K[�Aszy��˪ߕ,v��42���v��7�;��p�".ﮆ���r�����5kkL���_e�K��6�j�n���\ˮ��ȳMak�3�=:릎��o�8���]gS�A��y̧��5�k���;M��n����CVSHؽ��΂��x8���r�CA鷪���Bc��5�l��-$I6�L�(��"C4�ASmY$��d4M"$�h�f�p ��»f�ȳZ������q��b�=�s,c4�L�,,Ty��Z:�n�n�r��9)Z��8�m�1�nV�P�&_tͩk%ӗ/�+��
�O��o5z�}�(�T��V�����3� �ư�;���o����X��bo�s�읻�eI�a��&��A7���V���j�:�Ω5�܇z����f�Rsy|�oM�3��<���%���|��;.
��S��MM8�/�����g�x�3�9�
\n�qG�ܹt�R��}���#�"Uo�WU�m�X�0�eoK�7,
�j��i��3��!pP�c��Ƞ��m���:F�a�ܛ�a�@p���VLM1\)�]a���p5�re��j��O�V��Ű1Î�Q�!�[.�%55��A��g�ث���t�х�RmNY����"�����Lg4�����	��޽�3����gp.�c��ݷQ\��ݍQq��M�������*w�%L^�a�|ҡ�֣hY1�Ԭ��CrD4۾y(��UM{����Oe`�[]4=���z�52��[^���a ʷy뒬�ʡ�_)�����eѓM4+��m3Z�̄-Ǣ�/]43'���8�\�1x�dO0���\`{���JL���8w.R�Z��#f���T���-$���mr�R��uƍo0��� ��s2o��]V����.�5Vz�~��\���D�!
���V9,�'^}_W�}�ɒ�H�$б6#�涰�p�۷�� ,���um�3�/xb�3�`�&�U��o�]���]`ҭŦ��j�n�V�fY��æG|)v�s�R������h��V��
[����t����Q�}5A�s�a�L����N��Y����p��hg�NC�W:_�L�s���r� �I���w55��jm@��#[�7�Ã8�>Z�!���ּ�?zС�Gz����;q�c>��M�=�]�l[�7e%��;/k����E_ϼ*+���%��#&!��+��l���w b������Q�ُ8�����9��B���o�v^���vI쪛��25�=���dg=�6�k�5����g���Td��Dd;c�Ψ�6�J���n�[լ��07ô[I�V���b=+����s΢���xh��Ov�O�ai`��ݮ��vr�|��V^�kپ�;AhƖjJ���jr_^M(�����G�a���ֈ~9����گ�dߛ=�2�RL�Ag!�aܣ��O��@N���4.���wUg|y����o�P��΍��]��軰6kx�[1���R�c������hc��ow��쮾kuѕ����gm>��@0�q��/� �!��Tp;�i{x����N��Ԝ��X���}����}76�Ff@��^f����4�V7�
�P��X}N�UxB�{A{��ӎsU��	��GY��뭇	��Ș�`\Һ5^���X�\��s��W�xFde�xs�?t`�ᙘ5J��C9����m�+:�[�ye����^%˱��ľ��E9]��6UƲXA��ex�V���v@�2W���7��s����*�6	��lrl�k�;kg K�k�	�jSu�,L�D��U����*v�WKZ�	P���-��_G���ޯk��/�CO����Q�t@�1�"�z�rs8"�c��q��e�w��]��om$�=N�ohob~�7z�]`����*��'1��Hi�����Ϋ�E�ދy�&G���b)�� ��Ǡ�e���ue���&��|5o��޴����s�3��b�UK?c��k2߼�ׁ�vw,m����{BX�VE6�t��k��۵�������
\)�Ԟu�5������&b�XhC���W����8�F�V��'i1:�R��XZoܴ�������J����y75�x�B������ͼ��&��� .����fD�5hg������eޛ�8V�f�S��Y�-�������/����U�=�W�Ss��N-шd��ާ���'�k���W�|�h/d/o�����ٯ�9�pu�b�<��[!�x�T��>�^���5;�[���P�_^���r���]�W$��M���7K<��M�Kq.x���z=6!T����`�?B�>�z����\I/ڍf���Rr� QG�)��͂�jp"SذR�why��NFK����Q���߁*p�T\�1!w��'_8<��h�����o�w�`u�x`�U��J���V�l���������p"ws�Q�@���oW���؞���
U�C����^/�����_lg�H?<�����~՚7k6�PF��vw���GU�\�_x{ۭ"#=��JJ5t��ϵb9w}W���o���V�g8q���B�ھ���§Y��!�%�Z�d����V�7Ċo�N�uc�mf�0.)�5r�=6�-B�O�U��7z�<0�� oY\��-��s.�@�uaє;O0��hc�]�w�u��ع����Oe���0��Rʠ�:~�޿�r;<�D�|t{�[�f���wI9J4�sI�c�Xʋ��#��$�Kמ�zr���K��m���u|f���[	R^�ciV�졳��o�TUt��'�~O�Ǵz
U��4����S�>�h�h�]��>YqFo2y6��'u#7�=ݙ�mz�]ж�gK��îֻ��!����zT��:G�`G��Ҡ]��s�r|,"�����8C�������Q�띋��`��[�;V�����J��#��k˺���t��W�"���ۻ�����Y`�X~���1����&r'�ԕ2w^���I�V��z��{�oW��K��^#��b־�.6�������C7b��Ӄs�Fd:u��y�����}��ڞ���֠���ze[��:f�{��[��P��:t���^������~��WՖ�H�[yV���Q�w�.g8���扎�v
|c�:ܚ�BKL���n�����6�u�ՆǙ/��*�%���La�'��E�ݚ����f���,1ƴ_�5�m���gH��U&f�zԉ�ץ��,V��v� 5i1�[�M�G��͋�8��L`���[��`ŀ��:6N\j��"�[��K���w��MdaV�}Z�vT�����f��Ƣ$V툑�=��oRCwDG}���ۍw�ý4�gzG����T��vN5���}��5���xJ�0ywS�]N�lז{),�9d���V�3r]�`F�F� ��G����B��y�c�x{�Y������L\�%����ӏ'5>SNb��]�:�;���S�� ͙^z��<�X�J���.��NF����B��V5p϶��%yq���������_K�K*�Z�,��3]^�>�辔~�ϼ̩0m��O�ݯ}��Yͼ��&�h��6�����{�X�d��4��`ul�a����(`8<���@�
����/#K >8E}w�zݫ��_p�]���lSJ68Uv_w
9����W�W/hU���V��;-�_sO���~�~ۜ��L�o׵�~f���<01�q���r�����Mb<��G
��S�C�gG��qHT�ݐc#ovmh9@���bdJ�����/M3�G=Xx������S�C�ιY�ʉ����gt�9�XD�5q���Jh!��ֵ�	h�X��Fc��z��^��Z+�/pr�p��fs�?&��7�]�=��*|��p��/ݻnro�ۇ�c��gW�9��������x�W|��ѷIؖ=��K����Ko���O��ϖM�{�^�B}* ݺ}�g�&���~�s�t�Y����e�F���C�/�l����mě$M������E<�_���9�̼�UΏI�7�m<��;������Ǳ�'e��jE^��������=��9�v���[����٪��\���0��2�Z>�Ma�?T{k/�F�>��P�' �$�L:s7<�ͺ~d��]��n��RR�U,�}�z��΂����r͊�I����y�OK�n/�㨊<�]z�U�ȍ�[��o�s��S��	�"����v����I��W���ZG��^��t�o~�0�$�'aI��qLnE�s܆_V�X�v�b�#�U��h����w[ώ=�
���j�ugv�-��l���k^�]��kV��/��X[�L�[S�Q�0��o ���X�VG�u�����3�W:6�*�Ӝ,5����FAn빼�U�-g�tNz��Vq������6����MZ��;�f��;����U>����9�K��E-��p�]�<�r�_zL��_n5�ϔrV
����L��Ze��_5f&�4���N�hQ�n��l�4�S|ovT�뽪7�"nf�֗��y�Xw~^�/�i��L� �o@t[v372�`���z���g��
ڿ߳"�[���h���[�="{��-�l��T�B��>d-u�@�Vo�0��bY����F����zڜ�˘�A��s2|�2�|y7��>�����Y�=�/S�>Y;�s��W��}���/m+u��c�B�򵔳.ۥ|o�E�º(3Ҽr.=]���"�V���̢$�8����t���w-w�T}��)&�)Uɷ�����1wv���_ܩ:�1{�;��#֦X�9�Y�	�����t�~.�Ω�ncr��qD{{q��2F 8 �3��iJ�;z���i �amdy���H��]	��=�N���|5�]\�ڢ�7^>(u��pVwrZg_M�oKw4���qEC�T�0��M�3�Rw���5��Uyy�qs3r�M]^��+�����Fzz�L�F�8��F|,�5*���b�ȗ�yf#��C�M��c�^�P��Hڎ��"���I��H�e�)�J���/r�y��Qx툟Z�1���8 ol4��
5�0�i���oo�`�(�=����{õ�:�f�v�8�~���a2h���4N�>���ݫ�4���)L��A4�7~��۫4�B)��PV�Q�Nk�i�F��z�}�ëv6+�Np٘�4�8X��y����6|�V����͗�r�!�/�XŦ��Z3���D^����>��b��H���Uo��;5����F�v������ �?�����o�כ��=��l3����&�j>�`^�{��x)_�n���ݷ�Iq
�+�l�v�lJ�_wE^�=�?�Њz}��|��������׋T�5�8��)F$�׶���\��J��̯��8v�?�A�F���u.j�i�\�'̇��7Q:ؤ���it�]=�3GZ���T�e��j�ٕ+�����ϯ�	��S�S���%�4�uu�.�.���(�/$�_d}o4����]�Z�l�1�I_G�9���n���ջS�ŇI�9h��Vo9�9��ݟ�T��������a[�=|�3Y����˰']{����}VV���m��f)�3�%�ގq�q`��`l7v���i����M�@�Á��}o��}�(˲��νWP^�p��\ák��K>��Q�̎�H��=�
ܡ����Wכ;�������kPn+���%%��}�����Wɻ/�v�wMJo��+�Q�je�w���vh܄��-�[����}��Z���E��������j�c���R��J�>�~�x���o1X,���&�ܱВ����F�n������mS�	���e�U�o�y�ڢ|�iW�z�������]&W5$�IQn��p�8�Ν%�h�~_/x7k�jD�<����c�͑я���%��j�o���Am�U��O�ݏL�y�o��!����vt��2���)�N����	s���6Q�K�~�*,tХu�
�{1���h e�đ�iS'�%ҢR.3X%�hnE�6I�8U�e(b��,�&h=�,�*#����p��)e6��P��+��G+t����,��e�mDQ,���{�K�v�� 1�ù�ی��S��!��Q���2r�h
n��zU�}�A��繿_j�U�U�*�B#�匋�m}�w���Kr������z;�̽pF�i^Dy��~��sm�F�\⺤����:�8�B�}r�I����g >�qR%�൳�үI���'�����_]{���&\lI�"%]6�Y��=-����|*y�����(�n|��]�LP;1�v�X5���>�<�V��Ԉ�@�3t����m��w�3���z�9�}avK�߈xq3fUۉw��������{t����mob�Zs�xmg����-���W��lY�zUTwg����-���D:{�w|;�w݋l����m�"�ޱзV�]n��d�ǚ`œ��n�e\xT;�����jg�@3y�u��]���v�Ћ̢Pf�1��m��>��ٲ�̿�(i�9�ϫ,
�%3.�5{ێ�%լ<�,e:5\5�5VN���}-���L�]�F�-ѵA�\T��s�.K��j �KX�B�.L�K��YKU�1ݛ�f��u���[�]�U�7�y>�Hyw+{o��Z�2� ���"LJ��O�I:�"^ػ�2$������^N�/���f:��tn��)<����N]�t}�%p[U��B�҂9�#�ʝ�h�!hB.w��Q%��cH�1'�V�;ȓ/�u�;����O<�]ts�~�/���X���ݖv����徚V�p����C4���1���*/L��2j�J�m�J�.�:�����}���7�	Xm�2~Q>�������'W��_����㺷{e^��t�C'f��*9�[ڰ�f[���v�<fR�i��q���
�hN��'(9�*�~m���I˛��딑MٚƎ7�D=�֓j�\���Ҙ:���{��ڼ��V�OkK�Z�ֽ	έ	�2�<;�kb�Y��)��hK����j��ю�!&��b�����j}�f	�u���j4Ƚ��I��^6=��&+�j���i��y[�1b�}��9h�W-Vb����<��J�Υ���X䀏�@�(S����7�1�ٽYc��XL�F�ˣ)�Zz���aU��ދ��3mnZx���B��I;{�Z!l#�rVu)��=�%��l����zՋw���AtF>���]

��PM�cb.�Hw���r`�Z���h��#�v5"�خ��%�!�!�Vt��hF>K�߭C}\�up.�k�Ы$�YS~���(��\N>����:ȍR}f�t�$_G���K�(�`Q�JʒK}�V5C�g�V��yyI�qlVH�5d?����i����WV�Rܰh��rPή�Z Mb�5uri�چoMsR�H��tL�ld%�u��2�y�P�?�,�p����|�]f�O������'tC�d�]�m'��d<�5]��R������Z�������WZ�z���á*����wZ�[G0�f,����+��)�]'e�d�<�����+k�YZ;!f��>t-��n�*UX/���ĸ�se7;r��.[۳�]Wk���H��� �q�B�-y��J�
 �-����/X�U����BQV�Sf����o�Ԥ5Bh�1X/���X�>e_Q$i�a����{'a�W�mq��8�_Y}�jR���{�b��L敛�V�J�G6�*��/��fӮ�8�8IQڝ�N�r�]�s�~�����]�5m`���,�uZ|Zč���M�����9�p�Yt����:ځy'��D��:ovP�`K��ʨWꪯ߈Q���oi�|�	��%E+��뺂��r��;6E�8=��U�(��ψ���܎����������]��0721��B��kc�4!��,.*������Z�{�9U:^�YV^�[R��
��+V����mV#�W�N��4*�GC�qP��j�T�%��y���^le!�◺��ۍ����+	fϔ]�ȼ���qZ+�U�����fU��&��\ޝ�:r}5�����W�"K���	j��� h����/*u�q���wP~�٨�&'��z���O�ׯ�j�_8������A�χ�����O>:�[�����.�࿫Ӄz����4z����㴾�͗>�s �ko��E|�2_}�Ww[���sޙ��i����FƷ�۵[&�q���n{۽����x�k�~��'U��<��5uե޸��"tر�7P���8��W��v�F�����Nmw,�/�u_G]�>�P(��W���5\d�[�{��Y����=ܣwF��螬�z�I�m��(qέ�����4�'Jg���uc�S�l�Y%v��]+�v����O.q�w]8�]���8v�=�~~L{7����C�g�ދ��9��ѻ��Y�v�JT�ld�v:.�+�І����+��J�]nC�Ne���^+T��n{�b��+bNu랜�|^�ho�{��z��=�;�2�r٬�<N���sqv�+#G���z���ߣ���h.w��
��k�F��PnaK/��=�a��}���;�˓�4y���q�vzM/.P�fwƶ#ۡ��^u�2g�N��f��ܼ)w���1��v}��XiQ3��)��Pk �=vs6%�ܿ��������A'�1���
��M����2����Nw�{����t8�����1܁�߮�R��d�������I�Vpv%��&y��`���i�8�vlm�AX��Ȓ0�7���28g��X�c>�ڲboK;�HW�<�̺\�-��w73��5���Z��z鴲�.�Ȼ�eٚ��#��Xf~=���l����&q���2�/i���$x��Ҿ��	�Wn桙X�yl_��<��
:B��㊅Ϭ�1�0�'i>1d�[�W�1 �lΨ+I��Ū���R��΂���\�ߡ+��Re�U�N�m�L��
\�$���fи�.�u7�x�ϼ�,D���\/_GE�����L��O;ʍ�w.Nl6f*���ͪ��)F���y"k�������V��ջ���ղ���2X��Pâ��v
��j����n߳��w�B���X��Rt�n5���>˭�$@w�{��"�M�y'�({����=�۾�蜞�kZ�t�Oh��Ľo��QͭА�?E,NgoV���1���\f�[񃁝	oP�z_!�z�9Q�|T���e�^6׻^�� Ա�h���o��޹'cip˻G����lF�Zx
������
$Aw�zxd'0m�S=�$iu��}�\y_M����Pz�ju���P�CovK</V/9�S�C���w�7�=ŻE�G����1\�Va�Q����|�G:oUo�J�8�o?��TM�Ƕ�ym��w���(ۭ�ER$��X@wܸ�\W�痳d]mS�,)z���_s*���������ݒ���vp�u��Xҧ�t�g~�+	T����N@��w���)��fU��d侻�#�fgS-%����m��6�F�!���^�� ��޾.�s
*5�Z3kdPїx3���؜��<�ɇ_qr�;j��}T�F3�:� ��9^�?:�7�;�~���x�.0=��-DN˅꺂|�xz!��pϯ)@2���~���|�4�x�]n��||`|�u���=��¨������q7�<U0F=��z����XQ�ޣ~�o�mӦ�W�n���d�I�Z]f\w|�W]�<0.�o.�f�������HQ���;��B����}Q���W�8.���bŞu�w5	ީ�C�����ݾ��,aΝ�Ķ��?zy��gT�j����~J�[e���_X�1&��|��'�{��>�U^Ӊ�����T�^������=���Xݼw���U��;�$6Bn�s���~.�O�!^���W>\g�+��6|������=�v+���������!/@�������v�*�".3����rJ	Z���=��ś���*.^�S��A}o�&�D;q0�%6��ޚ�3�%29n��wI@V�J��|�v�M���{u�q��Y{W'w5��l��_�ץp�q۱�)�Owm�`'K���Y�g�~q�R{�*�.��A'���K�`a�����l\+��{�N03r*��X�X����w:�l�`y��o���Й�����>�QN����/��}����}| ��K�K��{^-���[�N��ٟ�����N������GN�6�<��:�������6�ːZC�n�����۬�G�jÃcY�y�|�s�۽�;������!^%�f�#��^KY�ꅱ~B3��f��g�s3���.�s���S1�32�G����{w�I���垦)���x&�Ҁ?_����:�,��)CO����FW�FK�h:�F3�i�����'V�eϴ�R��T�T߮[g>׮��I��=��'��t��m 7�O�V���k<��g~ϨJ�NӜ�_l�O�ob�S.׾�6b�q�fZ ^��^':�ѩ'5ӂ�B��nS\b;��+��=�j8e��!v��LnK$��cyK��y�Ͳn��8�wCG��9�c�\�q�����
�ڛ��AI�[5%���0��4`�%5�'�1O:�g�[�����kn��1��ü�	�r������9�J�r���B��?�޹v�7��P����+�}�z{%>���I'_�0�@!�7�v�b�����|�3Z�W�������o�Oe�����.�No!�z'��z}�� C}�.������Nv@pQ%��[�8���T����G��~��8�T\z�qT��+�3>�ﯩ/V��.��8��L����~�T?��nv��B7K��t����EF�0<���&�;�(o���qVqm��o`U�f�Ǆp[��圯Q���s��u�TQ��|���2hU��c��}�#���BɚyE#�y�nj��y��}�G<�λ�մ07\a��,���}�i�Y%Wg�.wj��ʜ�.��A��<���$9�)��vO��gu��J���������S$c#���������Q]v���z�yE��ڸ16�z��F1ʴh�o� �ݩMd�Ji�j�α�+ː�u��0Y��X�� �憭����h@D|�l��ji�se�+/(ޙ0���$��+.�31�WI�9*֞-۫�`$��H�)�v����ѽ��7ٯޙ��5޹zU	���p1'7t1>3��J�ތ������;���O��ܸ��8~J�����w�۲$T%��`��K�p��*�+FC�5p�?4��
�~��MP���.�,٦}隗�Z�U�l�:OL��~̿]�6)�l�G��۴���3leG��2<�-5����.����n��X=b�N�Y;^1o<��YVa���}ʳg�7��"�SW�~�R�0���Y��A�Nb���!��X���J���`����ST,ǯ��-F7�b����v��_�
P
Yb��14��,���o�F�,0ǐ��U.����o��ξ�Iΰ}.n�eK�~7�&-Ќ묑����o�1��>���O����;���u.�3�v�ӯ���G=umT�M�ko�n'�>ɗ���_�$���GGG��aW�\��x)����3�߄�g��Š�;�9t�2�٪���,k�Ywi�PT�n�f�<�m�Zs�l{3��4F%t�Ǥ̬��i��+�ݵ���3C�\��f=���s��u6����pX:21:��D+�=�vb��4;A]F�r��'V;!�\Hc>�S{��^�qec��e�X�\���}8�{�y:�� n�����#d��M03���Ev{}Ia$��ʧ�FQ~��~����y��S�&�&���n�Џ:�>�w ��b6a��cHGƮ�^u�Z�ޜ��1_6�+k��j��=�eLL�����VY�5�{3>�����8�>��1���E�Jniq扴FY#0dQ��~�p�=�u��Fu�����2q��>1z_ol�@�nxӡ��%$�[���rwV�{�9��^�@:Ew��g�?Om���=S���ߛkf�E��^j�B��G�=�mM[�t~��2�I^{�SP��!���Gvøv�E��WS��U�u�<��
��ğ�s����ƀ�>�klN{��ϖ��;���M?K�����Ŭ"�c����'�5��]\�-;�اtk.;"��\-��핈j̾�&̑l;
�f\cT�����D�,Ь�݌�9�Y���Z5U:��۩~�+�
��)r���+r&�/x�iq��H� -ݬ�����(���bq�q����r�X�s�K�K�of�(�A������*]���9Η<��~n���!�8�/jWC��i�]9B�>��y\�h�w�0�1ޚ̀�7��>�K���+c]���x���m�O[{z�6MX�}�=y�b�qE�l��9��/Bc&���ύ]�U��=�d^�Ӟڻ";�'Q��W���rٷqs�/H�o+�Nѯ$�K�'�X3}CM�T��ѵj�H�C�7��Nў�g)���!��ׅ�_z?��w_e�	������|n��v��Le���wwJ弔l��=�h1��>u�4�ńW�T_9��S��u5�m��'�
�6�==��|�:���W;�\�u��s��U��O[�}��hO�촕�k���q��:=C|E�k٢m�u��j��_W�C��ٽ��zL���ٰ�U�4o�j��t���Q����c�	S���x�`/�U�#fV��{J��έ�Van���	J�������Sevf��L*�V忮��
^�j�0a#��V�4�G�ɋ��:c\#�2���l���Z�S\�Q��d����%:>#p�����/��ح�iX��r֑��o�r�K��4Z�~ݵ�����Z�����g���<`ث.+���Sٻ��+qk�3�{Q{^U8�����<���|��ՋN�a�2h�fB�Bf=[ެB^����Wg�Eo��?֗���
�g���mYzNhJ��,��(\Y��A�d��z\zr�����z��n�t�1�_w�^�$��wܡ��
|Z�A��:���rۭ��@�x�ܨ)�wt�;�-+ش�a���;�E5KJ���'�qeC���P�T�����ݖB
��ܮ��Ə�_d�>�m��ţ��������WN��"�ƹz�ys�����ZÏ�>�Y�z��_p�.��n"t��Ħ�k���NM��.�M�G�D�^��k�ȏ�tk5/�F�s�x�S����^OI��1���"�g�yסн��'.�w�Y_�=������מ�����h�έ�)��3M*�}^�g=7A�F���ʲ5����r���U]o`�[�Ӯt���V����5��
p��N�'>��g]ں�:��*Y=q��]<�7�4���2*ʛ�	I�e
t��Ŏ(��9Å��/����;�Վ"J<���._���n�kj�㛀mf�j/v�X�fy@�Z;���̄�F.ݭ����/���@��k�v��@�Ѥ���bSw�YU�=w�=7��k�.͸�9.�2+��ص^�z��\]fH�Sᚐ�|D��os�k~�]{�Ϗ��]>�	�dHO�	 I?����$����B��!	I!d ���2Ձ!@/���?��$�5����$	'��ĀII��	 I?����?�����}�}��?���?�������~����\�����8�.�s O�@An��ʋ#d���Ճ�~U���Kġ�jضq��,4�+A�[�������\XVg�q^��a��Y	���7!�mI��4-b�1�I��Ł ��$��Wf@dtQ��(�9��)V3v�^ ndz�ӎ�!�e[9�\�uKCn�$� ��D��]�ݛ�bًh�j��l�n�PRKv��%ˊ����b~�i�� �Q6S̙ER���(m���k%��!쫪�	*Դ�zr�֝����=���'3e˥j��*Pi����W���]aڼ�0�M�	[�tJUL7´?�jͺD6l�T,��bn�1`Ä^��D�)@0��K��?aj�d8m�w2�֌���+j��-ٚ���Y���m��	��"H��Y��ܳ�A<��5X�hƝ�Ye!vBKŮ jV�q�Y�v1
�����GC{2ݍ6j@2�.h�)�Qʻ���-�O�v�R�֮&����q-32m�w�2��X��RƘ�woX��2�u �	�|�eh��)GA1摍��`l�-1b������;��p�LMtl�"�.K��X�2C(*pҫ���T^<��5Xh�V�Ǧ��S�d�28���D7�$���1*)�4,����6��Tm�(c#�voM�@l˼jQG:(Gjӳ���=f�ZM
����P�I͊�n�-f����b�t5B�cV�������V�ܧla���E���)�^�2
Z��ø�yB��Q���-�&�Sv��Z��QCb���K�L�N�j<��[�3�ą�(�4��k2!u��͵c#m���֎� Ȣ�Chu#X^7"zl����J�-���b��C��S�(nj��̫su�
IdtsKຌ%�y��\Ku�;X[���&e/��[�U�P�1�R�#u�v�&��cׯ���x�T���j�q�V��w����A��׳(��@QQu������cT���8�-v�/��J.�A�nJj[�!��۵��m���01�S�Q%2+Hãl��@5�<	⬸�ZZ���O�28^��ܐR���VӅ��q@����՘ z$����������݂b�XU1]��Z׃"a�mP�!�͂^����kn�B6����'���2VRȫ-o�
Z4�{��-�J��g�`�ô��kKo5Y:kSˁ�����`!ct�T
�F������	)�5��`��ۆ�@�`h<wn�b4�#�@tl�t��Ү[z�^Y�Q����0�(��8�{�r<J��Qp���6+	!���C�ol���cTB�*�
`�'n�-Wz���I�b;��B!Y" ��ɕ���u	�!Yٷj�eY٪=-�����ن#I��f�ҍ,.�6��:6�-i�y��
V\zҴu�ԍ#���r���̌ˇ�XŠ�D+:1�oF%Y��xӵ[�(�C��A�6��Nm��gr\y�ҲRPCU�t%�^����,�ܶ��v��e��Y{[X�%P����9�i䗅P�Icv�p	�u+;�[���^�+#W�J`���ZjC�Xe�T���&�m�L��tGB]��;�)���@/�9%i��wTQ�
)�%\�%�pb$�o1T_mv�Y8�	�E��V��:�~?��:0-�ۘ1`f�Đֶ�0�q%T�	�.�[�X����bh�B8��v��T��Uٗ��̼,����'k&���[`*˛�����j�'lX7k!�oAw�9���~���;�=�mĬ�v�!�B�yM���VZ̼"	ıNP�=�e�����' �דh�����m:OU ŕ��8]�+@kU��,ՕB�[;�hm�2n�z�S$�[�0��ݒq�U	xӀ�`q�;DZ��)-������(���(Z׫63��Jn�n� HZ@���e,��̖5�܄��CNES�����0ۣ#R���Zon�y0mǟ�F��Ƥ�ņ�5�MKis	o�,���&N^:EQ�)"�{t��� H��b���Z�z��mmhz^U��P�w���Y?Bij��mQ�vn��F[Bb;��4IVS��)�q��D�4�XG.lV�4@z�(�#×lܑm�D][m���bm�(�On���0�_ؙ3V:��]ЗhQ�Ĉ�cˇV�������K�O?R��xn�qR�Y{�2A�
`n�Ue �A%�˻�҆�1�X{ {Xr�14���	1t%�O�t��w���©%sU��]=w���-����1o�Iz��YT�Ƴ46^Ktf��NX���ѷY��DQݰ��z�z������@`�i�meт���V[Ӻ�-��!XCv6��ę���jȴ'ke�UV�ʘ�#�;Φ������ I�D 	$ d #!$�H ��B�$�H$d$�$��!$�	!$�	0�� HD�$$'����� @��g����ƈ�$����������@$�$�ƿ�$�$�II��� II��5� Hi  ���ه?�~׳f�	 I?��HO�O��}�I �����$�����g�����<�$	&m?������� ����$	?_���b��L��6B�p�� � ���@  nO���Z������kMjJ̭��;�ON��P�    i�γ�k�֎ 3Xӧl:ph����B
	]ele�T
�QU]d@ ���$�fh���    B���R ����K�T�j=v5"E� @K�  ��W����{{�}��[UT��um��f��&�Z���*�k[ �>���o�     @  ����h<��tC��>����9��������5��n9�Ie�����L����^o^��뼝��;]{����t�������d����}w�z�wW�ӻ�n��w�ٷ�{[׵]�=c�t���;n�n����Jn���p�z:޽���3Ï�ʠ������H(=A��� }� PA�������Ҩ>�C�hAB�aAA��>�V�v�ۆ�z��v�����iI���g��/g�j���Ȼs�2�%a���T���4���R���mJs�I	Zt��	�W hj5L�/yl͙P�y��]t����:{n��W;����V�ms�7v�+[����͵*����	ɺ��ӯ]�Qͭ�w^�պ뻫�v^�^�Q������*��k�֫c[n�t����Q���������7�{ڕ]e�ӏ2�m�L)��#]�G{�jԦhW- 7p��B�^5�{�ֶXt7�j�تz<;�u��{Sܽ�mUQ�G�! ������Ψ�w4q���wq��κ�{8�k����w�m�+���6h����j�{�g<�t7�uָǗi�k��;���B�%r���I9R��%xQ�J�}�oc�W���:��OC�z�uX�]d.����**���Z
�P@ض�ky]�w�Z�z��i�vN��_@뽚+�+Km�fm�v]�ԙ�v60��`����q]�ۊ��ݕ�T^�!p�����<Ws����8҅;9N4([z�%�"��.�T�T��lJ�!$�v�t��%�5�^���3:�<�v/Z��i�i�p�f�Ѣ�v��QF�r�v���\�	����e���N� w��%U�ʥJ&kjk`�*����Eh��V�Ч�3����5��8� �)�OF�oS��בCN�,z(7�W��$�^��TT7�U^�U*H��I*���{�Ҕ{�\�B����nzد'y������ެ=t�ov^�r`y i��gzh�mZ;���F��A�Ұ �w�_	��(i���ѫecm@	P�V`6�@ ��h�T� h T�!�%*�h � �b�  �?f�IJ��   "�� J�F���$�A	Ra21z�?7���~ɏ�����F�ԓLl}_,q�l��#������s1��;g�|���$!I3��t�����@ 	!��HBO��!$���!I?�@��$��HBO��$��_��HO�4�n����s*f�5��a��ն�ܼ'ď8=�����&�	Xa%I
P�H`�3&^�y��7����������O^!	�4��'�n��s]s��鸶@����f�
LKr<ޛ���,�5]-��<�0-[�I�;`��m^�$��=3ND���	[�Go�c��Zu�q:�r����յ��@eV6-�O�].b���k6+�7�ؼ�;��y�ǻ��+������x�V{���O�`+����i����ߒ��� ��oQ[V�#k8x*�x�Y4�6�g,��z;�������C/p�JBH��� �#{I�wf���7滽y�k�ޅ1*H<�bN���~��B���{2�4ہYיA��c8�B9l����;s� ��C��0W��?U�a\kW�����!zql�ܻ:�Z��P�yf��N"�wY��1@1��^+OP!V�8�؎��ߘ�V6
�m��-���(jf��M����w-�@U�s.�om{����6ph�E(��"<˱_�]�6ш�i�j��W,�ܻ�n�:������1w�M�%��u_� 6�R7v���?��� �m�A:)������x����6@�h"g���\���y�oRX���a��vk"����O5���|��j��YȈ�/n��B˧�$���ڣ�Xq��d���lP�ɦ^r�u��v�֏7L��<�{5��\��;'�]{è/
�W����m�f�k��{��m��z�6k)��'<���).Y�ne�I��`VAg�W�5����v�m��<���z,Wm�f^]~
�Sl�d$6�Z�7�\���D�v�[f�Z�~#�V
����0��9��!ɀ��t�Mc7D��;��:��D3P�����ڕJ'mg#xiM�y��A��*�6ԣ��Ӯr��cf�Yv6�!����`'o5)d>��u{ԃ҆���{Ef�[u��<��sk�l٪x��xAd��O�y�`���H,@��i�4hs�x�m5�^Y|�ft��q��
Ae�Q%aYP��I��M2z���0ACKkU��e���V%bMҢ�o2^�[]դ^���`�*��sB�pǉ�&�_<��0���uL��uV����u] 6��Lr�x
�y�Ù��q�Z���+�F���	�f��B�y�T�F�,�X�j�5V���=M�0Y�j{-�YkBWwi���Y��M4�1��7V�!���(≕��H(�#���꠬m��m�7)(u^�Wtue�U��aJ��_�~��,k�kLCN&&�!�f�Y�s%g5ךuCZs-�9��B��s2�Q�o7K�<n��n�����T��U��*�Ty��<9�om^mI�i�lyO%��P�T���X-<�O6�+m�+���p�K�u��xSd��ɶ��{�{��Lך�m�B��1�vL��o�f��a�0Hyw�޷��{��<�$�q��ig�{�$�z����r�����|pyT�*�JB�e�a�/��;�C[�a�f�I�v�I<x�įY+ ���w��8s�̽S����[�^��7�v��v]��U�$5��שP�TD��E����+X!iUcYXV�+��XT+���Ң%�Q�R��[T�[T(�ڪ��UFҊ�Yd�TFұU��-j��m�|7�NQ�G��n2�FŖ+C�������]�L��;@�=53�3��l��h��3
Rd.A�[�C
1����"(=[�&+ ��õ�-M%��Uz�Z��ON����	i��5�6�9�s9Ӛ�u��Ad0F�X�k5j ��cH�l1*�TG����j�-�����d��L,+d:És���y��a���h�W�I�� /7c�$�au�-�Nڵ����ić�A�ڊ��<z���R�ܣ?^L�&�c�ռzp�eh#��(��ތ�۴,�ӟ�j�`�����c�i
���y-���k�xxe~��c2$��x�Ǝn,9�+:��3���os��z��Zy�4�I"���������A� �TF@U��d�u�i�WISE��,�a��6�@ :*E ��Yb�QQD �A�
(�U�mE�U
�Ŷ�YZ�&�TE1�5
1��#*J��m/TM%�ul�K�Fc
�i`[@�*J�*�aD�V1�*&Z��
�U�DPĬGQ�B�ĕ1(�8�FT(ƥ
�\eDS,J�k%�5��Q��j��eE-��h��
�[Q�9lE1�1�ʈ�*�ed�QfZR�QC)`���&�"��T�ii-��JɌ�-��,�Ae�QT�F�A�lTq("VQP��L��0������T(�IS-U&%IZ���(�"L&�T"H
�`�B�
��V$ �#%BPAF���d�AD`)!@XB�d�H)""�AAA(#U#�BāXUE��A�+P�*�6�*IX�ŕ�ţUe���[`$����T��De�U[)E�E�%���R�m)#�ʪQ��$PQd�@��B�E#K
�l �
@U�+��Y`�a[#�Z5V�Q(_��5���ʝ�W,-�z=6��<F�h���mf�Y����F������z0�j]l�J�W8��]�����3�`�UH]N+�?d�۱�x<���Y[r�Lܢ/6�j/aM�$�����)���+��WG���2e@���/p�`�7���)�9YW��eC�l"�(D�cie8n��u��{3pQ�I����C��X�Z�tP�����e*˾;N�O�J�X-�Y�+w��,dkyȮ"�bZ��K��Q3 �n��Oڥ�����N�/40S�0[�vʹ9�Vig�
�d��P��'M��[t�^��o"0X�[��="@wKi��~��A�|���]�y���9�����^��e��B� �,z��h܉SЮP�ab�l��f���+$н)�z4JL�˩�#��Y3p��Z@я�%�i;��l F�5lK�u��ZO#d��o!�E`�v��g%�hܛKf��Y���KN���8*�X7X L8���JvJƤ��/��QAe�������,]"f�E�g��#�ᨣB�P�pVP痶����@#R�nٷ�6]Nn��a����X�������0Ky���:�n�9�Ԛ���Z�ܹ�t�)�{�Zٗy��&.�,1�K�Z������Òn��S���+�\j�of�4�m�t��~Aڛ��GD��������Ť��+%<���cr�f0E��[n��#�͒�je����q��a��3��G^��+7ڱc�x[��L����oC�k�v$�:�#������a�}Z��p���AЮ��,�rPk��F/�Ywqs�*�rYy�V(^̤�k@�p�NƬ�]A�k��1�h��Ѹ^���ƯQ�ZB)ww��6E8��h�R���c�v�l�� ��R��V�����.f5Ls"���zlh}��hy�i�а�P˻5�c+#��:�j�CQ͚[�%�����E�]Bh�
m(ؼ&[ǎ#N�^l�+h�U2�6�nS�6BӨ�]y���׾-ya�q�B��-�aFJ�UVV��j1[B�6�u��oϻq�i˚�{.��%�d�YU��A)Uf�-���h���B��-*iKkA���+*�Z"�hQeKm�
ʨ�����<:k8�K��PY�a|�wz��X�Y�B��5����t�:�]�:���;z�<f�k6����{��+ �听���+�3����1-�u���e�
��bcQ�ZX&�+j�\��8�F�E��`�������y♄�5�+ �\0s���f��բV��h�S��鼲5,�*�h����[��0�hB����qgꌙ��h�.�6�x2;��h�tX�;�fܬT�ȶ�l��kU�T�G?"�i�Sq!�����Ɋ��8��A�a�����W�����9`�M0��� �z��d��c�V6��J�,4n�r#7s)X�tC�62���~�!Kb��+Z"��U2�AJ���ImU+Y+k�4t�oʼ��^�W6���M�b�E��5�x�c��X,]�o��n�j��v`ۭ��^^�(�l�M�`���P�ͣF�v�$m��B)�5HM���]7h��2��v��l稾.�.�]b�uCo�.������O��武��Cr�^�h+V^T-T�������a������Q33?��uN�b� }_�jG�A��:�� o`:�U,�m���8m6�
������ۈ����cI����)����C}G}�� �`,��yAR�_����r<Վj1#noU��)-��E�*?�2�RW��ŤYn������"��Y�ӻAe�)cZCCDf\�"�3i~` ^�̉�j���g
�pV��P˓B$f�WO.���K�|�pecM�=�3��Z��*;��BnCZ����4��1۩gD��WIhI@ �3����O7�;��OVV�#Z,����ڬKlX�d°� �#+O<��5�9��o������y�PuaXT1
��w���S�XW8�cw��56����g�W�����Dn����-�&�ky�u����Z7]�;y��l�w�Bu�x²e� �v��f:�l��t7}�c��k}�)
����и"�/�F��l:��-��W��e��6`ɻb��1�׎ݕ�)/ߓ!�H,��N�z��\WZ�/nJ,\$E�v����~�麎7a�NæΕ�ɢ��74F���e��p#o٭�g2�7�m��?U;F.�vf
dN�m�1Jh����ר�&�]�,X�u�7�9�ʪa�x�(�`d���b�V���߿Ah_��8I�Kzի�YҐ×�Պ�q��j}Noj�7�t��X{���O{:�˙)Z�xzY�P��U���
Z�Ӊ.\��T��v3K1���f�Mfdt����*�(���fu�����\��}v��]���J�a7�u�d��)���u��8N�sE��;n�3y��߂g�[��&X�#�n"ƙ��Ĭ�1�܉�g���U�F���wM�F�yms��1�[e���h���I�h�5���R��G_b5�N��S6�έ��͚�L黺�@Kr���$
f4�/,���%�j��F�:���3��:�65f�WwY�sN�[
��^c���K�|��ރM���u��\�ˣ2K�sXz9I�M�Ds��7X��b�)2�W)vG��ЯP=�����2Jjp��4�u��)���}����0�zψ��\�����]�dV���R�#�h�Ժ7xJ��eM�g���������S	�n�f���9qe����yN񷪯��EK83�'qY{�de`Yz3�e>�{�a�����.NJ�H2��pe�x�n�nT����fܸ��)�I�b�0+��x;]��f�v�\f���cm���>�2���s��p}�)���T���EC��d})DlK= B^ND<,,��.�˨1��\��Y�m�j�{�W[ii[7	nI<OL�+�ŕ��ި�#�����߸hDm��+��҅8W\�w��)�݃iYbɝ�+��I�b�LL�}c�Al�$�LU�Mf�=�6���z������h���ެX$!�1�.�e�r')d>�Fa7w�D�6���蜊L1���g>�)�[�9*����;��v͍r�=���*��z�2��KrJ���nm��]��u��mdD�����
��7��ɜ�uY x��\T��b���m8��y��e(7��v�:6_q�Ly�n9�k�*�J�x/<kt=AU���C�mr4�5j.\F�ܘ躹���w�WmP���)�oN�Jvr�D��衽�zSʝ+���.b(AI��t�� x��v�M�Q0��a	�pJ�mhnc������vp�)�4,�4�*՗Ҋ!��l����2��9"�Y�5��5�T�[�(Q5�&a�9�t�#q�Z�N�&�ں� [������JTk4��+���%u}BC��/u���K5����;�f�\�.��|�:f;S��c�;���S}�ņ���Zw#��"<l3�nU�;M��7�%j���A�؀)r��W�9��H
�+)��Y'�&;2�[K%�E�v1e`�gwd
�^����9��{�Y�ڕ1���u�1Z+�����k%Vؑ伐k�#0LN�v�j,Y�Z$x��\$Ҧ5vi�ѭMgM:�aZh$�c�ڽ5��Q��=����6��؈"�m��7t�F�f��y�q��y�r��x�n�ə}#oE<AYK��C3:��彀�6_�qgzT7I������s�d.f�`�'��ĎRM��z�I,]c�Bma3Vߑ�V�ot�x�	���xd	�M�M�K�}rg���:��sh<<;�l��ON>���>�
�o��'>��$�;
��2��~\n��E����.��u+���S���}�G�ZZzHkK�|Mu���/b���Qn�ERx�%-��v(Ѽ9�6;{y��jr���t}���\7���=Sq:=�Z��>B$����k4����lk5�,7Y�9��'[8�X�v�lz�U+�5�E�ƛ�/��]E‍��J�P�y-*d]���ڡ�:��]B��{D��Q���R7`ݗ|��u*�Ꮨ=�	K#c�_L�?32��
g5]����S���LrF�=����s]З�k+A�V~ޚDӇ{)*Q7�h�Un��}Os=�s7\ؼ��M�����D�q��|����^J��W*RGzҽɭf��$N��g^f�����8v+w5�ĭ�q��0��Pd�p��ƭDaʷ��"�QAt����;-��+�Җ��f5��n�Gx⡯1jY%�}7I�|M���N�f�d��B��6�dX��du6y7���%�{M�C7[-3p�Bg �X�e��]�tF�vl��3�g�� �����ռ��a�SJ�ur�޼	
�L�:�
@v#�pٳ�݉�.�n�4g^ �{�\�q�Zm����͐�-��]����.�\촂I��X����;9���hk�1j8�"�^Tz����Daᆋ!��QL�0+9�h.-q�i}coo�*'�eq��"�tᆶ��EXQ�t���

Y�#4B�I4�hg#(�A"(��ړx�g�)�լ�y԰[��}�p�2�t6ج��S��6��.��N��,�+н�vo(�]��6
�n�:է}�=��r��f��`�Y[�u��A[��ƞ�0�j�{u��T�]j��}n�v�.���u	��\����n:i��to� �Vn��ȺH݌K��K�uܻ��)ћ�����ꖡ�FKo��r0�n�/B�:��O\׶����g7�4�}�AGwh�6�^/�w5K ���-R��3��)�;z�u���Oev�l�$v�5:'[}�Ktup�ɳ�7c!ކ$[pTNT��a�S_v��;�#�8Ʊ)cɷ�)I���J��fT�ћ���]��i��[
qK-c;�x�x�f)�y�֕[���]����䨶� c	;a]VI�/c��Y������]��u;w���}ձh$��vj�ECE�����s�+9��b9�S�T:�Q+g]˜׍P��|b�J�
��,Ue'�츼ո�΢Ѽ��da].O._^��NW��=���p�M�Rn`�����WH[�D.��e�X���;tӂ��w�2��c�� �v�B���V��:p���6�	Հ�*pK��Z��,��;�;]L�j�\��*�Y�F��fsej,�g[��Yx�(��)3��S�s�Є'&�\)����'�΀.�6)�슭�nn-R�f�%A۴���C`k]�a��|������g\&�˃���w	Z!�G�v	�B^CIkV� �jZۤ�n����r��oW<�6�wH)j�������4:Uհ��bR��[򼻎�*`Fٻ%LKm�ۙ$ ��m�1!$��"iL��`�� �`   ��m�      m���ZI�~ Ȁ HL�d m�IL��-��9S)� �`6��Rlm� 	�l�$1��                   l$ �`   !�F�� m ��Ȁm9       d�  @%    � r� @���         	&6   �m�6�m��m�     	 @`  4��6� � ە)�mB 6� �    �6�@  �ۑ�����	L�  �� ��s-��!�RO���n[L�����i�� �(!KP��iN@Ā  m�              �@ $� ���$�!�  �$�   ��I  0 �     d�m�      H  ��   � �  �  0 �     d�  @ H    lH r� 0 �     d�  @ H              H  ��d�  �����%�%&�m� �ۖĚS( n  H�b [�N   � ��`'3)�hP�`�d�I�ā��l%��c 6� @ 6�     � $��    H  M�� @   �l�7��A2�{��~��?�:v%b�
����|Z�� ��q�y�$QɷJ�$����b��Z�dR��C��uYm+��މ���L����R�ۭD����,��P�8���y)#oH1f�z�Ueb�^eU��3(�Fn�mv:|R櫱�V�ȻaЧr�u��v�G�g#ڑ�vG����$x����5Z�ǯ)��g%�䄝��4��S���jx�w��3i^��"R�=S*��KN_���=5��r�]�3��"z�f:��N��r놮�r	#N�ٔ*������O��fʿ����]�I���=�S5[�T��w�Ru��T����Ǚ��B��\0�����oZx6��"����r�-�W�Z�<�(:���w^�_��Ħb�7C��cd�
"Ƀa7�V�\q��e����i]���Y�LL�Y�u�+�*��;�~�5m]<k��.���85pL�9����Z�^�F�^�5��0g��L�|�վܘb���i��	}�����A\�4����#[��ee17�5���Z���tp�"�2,��kVw_r��r��R�F��ڲX-����u����mỵ����ܾ#�4�)�)��zN�;�ڕwS�U�(�x�:f<�p�t�N0l�icΥ�:K����h9�[3���n�f�,t5T%�t�kz�`��[�Y���X��BgP��ݽ��>D��y�z��l԰�����[��� >�fP�]s /�n�3\���;V�)B�퐫]�P���f 7��&�R�I��F9�3-7"@��D7-L�(`)�(bC$h        �     � m�6$"d��-�9j�I�9��e˙pЈ�jY.�`�clm��$e���\˔�L��I0�� ����D'
[�9R��$�&�)%���%)M6� $�I2�#ci	J#v��*��s����fAƋ�uJM�p�pTq�;�Ŵ&��b3Y�:�ss�n�����cǯIJwV��ڝdٹ�ݺ��]�&�*�J�[P�p�8��]t���Y�mgH\�Y�����s��5��1�:&�X{��gr�8phȪ�6���,T�T�F~VVX�S΂��8��,�5m�}�j�e��vo��,$�ԝ��Ii�ж|�
��k�t���S�C.�b�{��6. %v���^���%�vÄU��Fd�gAǮ�y�r����!GTyk���̩Z;�Ei���8N�J�[!X�僄�\㩔l�X�bB�T�'Y�s#�H�c�w�;OC��k�z���,�b��Y�#fnGW��B��],Wp\=6��J�� ���Ե��"�@�q�繩�����䥿�O& �2 �6        $��1$�I�M1�3���7#�
2)&%�X	�$4۔  mÁ�$�Ogr�(�4������LH����D�vݸ+r�0���hB� >���[��}�ZĝK�B.�"�[d�zD��S�,�ovm���944�,����c��75;]��G#+��u���8�Cb�t�+]``�i��RhM�Y��&vv��/#���t̷w�9�s����N�lf(V)@3�F�@��^g9��KVʻj�qބ�T�án�4z�#��2R�,�	��A�G�y\L�X��skN�k�Qh��uݭ��*�*�k��JH$*b��X�]&���;�$}PJ`�d1Gu���
��27d�v����n�1q0�=gS�9Xy��K�X�Jf�yF�ꮵ'��_cDh`��/�8r�X�T�g�/����ߋѐ��j3�傡	f%� ��|8R�#��p���D��Am�)�?��*�A^C�b�uBI�HC�i[wg���S�翺A���5ըU��N+9`�i��PS`ݙw�*��yW:V�nu�M��]{��I<�D7�ٽ��r��y�ݙ�L�%�V����Ń�ލ���J�{��S3,[��`�d�6۹(Q��aRɽ��;�h�Պv�k��3��]�� ï����f�_>�WsL�Vd6�+��΢1f�N�QS��ջ]1
�wV���reT|�2쌪�ѕ:����v��L��"��e��^�t��kKZ��ܺŃ �(ف�SSʺTV't�i�g�j���[���[����ğ3�n�yO��8S�M+�� �=w���Mr�yFy���8�k�j���.�JC5��ҵ��"�G*:W��UM�ODc�rU,"��IUw%�r.��i��lv*.vә����S�$a;Ns���l��0:=Y�a��|I]��h�G���8UiA��kU�e��T���A�c/pG%���ŵ��6ѭF�9W�����F��g"���v�wVl��.Cniͨ�/:�*+�q(hLJ��8ֲ��vB�;s�A��]	Ԓ���/=��������;����H�!*����78Df+�mz�2�;N��]6[dS<�-�yW{Q�#�KE�ޗ\��+jVu�Rv��"P�~�U�����ʃ9w=���Ў�����T�LW׃�
�#��ݽ����fћ��=�Y�$N���6U]�rsU��0C�q9����Z�1���Y4"��	 rW0+[��/:�e���Μn���U�.�Y&��k����x3t��Y\������5�iэ����1��9�͙��/�(�ˏM��c)�:V�#�t�Z��r,畷(V�ÂgC%�+�<�Q�qZ�R���aa��F�SA|�����]՜rV6�����*�UUY������_*��%�J��%Ӵ.սC��Q���I��҉��&��d��9��N�N������.|m��8-�Vc ���{v�m�ؖ��7q�s��0S���j��]�o�k�/�����9��Y�0$!	'�`IBIS��$�$6I$���BI�n��R�d���@�Y �$!�@���	"��L1$��	9BB��i�@� 2I8��j�H$�,���������g�a	��I���M�� ��I�P8 y�,�� �	8��,n�wfy�`d@�(J��VN Q���<B@2Nj��Ow�	*�XM$ެ#�p�01���lY1�.��@��8�hL���d&�I�;{���d�ys&$6�\��I�,�;���& w){`f��k�CĚ�Mn�H���$�u��Ww�Qf�q<N$ެ1����=�r��4���u	�oyA_)��I[���Ѽ�+��3k���M��;�q�FL�h�3��h�\�tN3&�(���aj[<���)`mz�,�Cޥ~t<y�����d���z�6���N8ɤәej>Z$�3Z��<,RS��E=a�_i��ci� v�%Vi��am�ʅ3�k�u�w�`s��A��N\�6i4�嘛����b�}��JW)Cyg����w�D�9���� �1姏�h��eM!�)M2��Mssn���|=�C������,���M��j��n�̇9��g=�wg0�r�ؼE�ˆ��dm&[̤�e�,��g���O��\���(Jd^��`Z;vW�U�~�D�@d�\�I|�H�,ڱ5QB$x���m�S�,���/�os8�i�S��u��f���v���iR�y�~&я>�g�6a����>c�d�Gj�f�u���I�O2�M�U<t�Zgw�����3jiP�6�(����[�>��N�%�V ��iP�EjH�*HP�@	
���Y���Ⱦ.���z��/��]{+��5BM�	��"^��,��b裬7����y�0/}���f�n�˽�[}5M������'�ܬ{�6h�.>� ����7hW�*��u>�d+���Ϯ��԰�2�1�����T9WvԀP��е[�G��R�CBt��"�^v_����
���T,�9R*c��`����}�)gY���-
�eL!�b���.�NJo��n�*���"}fq˷��[����5���rn���l̦����U��or��b:�l��t�T����I i��b2��K#%�7������3U�zI�C��t����DUi�:_J"�٥T��6�����9�!�A���j��횞>�RfM��y��Bm��p]�s�T��\m��B�L9�r���b������*��0'�O'[C���	�U�oq��c=�]`Jd�r;������-<J�C*�؍\4j�AI��-��R�[�7u܃Yۥ���C���t�V���xy�h�zF`C����T
%m��`���m�A@�A�Ѽ���kYT,�W�l����R�@J
��mk�꼴OR����f7�Ѵuؿ�������I���P����Ὂ��U�)�a��x.����U�Ƣ;�.�I�A�`^���7	_<�BP�/�q��,^��];���+�L��&�.z�ZN��U`z��)���5J|�p�.����4�݅�	�i`� <�PV�#R�X�뺁���AN�M�E5�P}x�FBD�\7]Y��eP?��D�`�}�C�nil��K�6���j7Q\�^�R����8�6r-�EŲ��ka���r������\
/e�@�2��{n�䒕(\*�:.���댶m�j�-v<'zݚ|mm�;��Q�g����+��!�����L��5y�g)
���[�W:b.���: �I�b�4WkX��ѭ���c��1Qfj��볍�[�h�60�)��/e��}.��bͺtO��I;b���Q��U
���Vi��Z	T �١]�y�h'�e���(0m�{M	�wu�*02�fP��0hP#�����V
 "�x�D���L�>�]N�+��+���`�s�ݠL�0N9o	��ױ
���M$���7*8()�8��11t��Ķ^`��
��Y�By�ImP�eE��m�ˍՈ*ݣYKMX� ����1z��A�su�\�0�:]��uГ�h$��t�c4%�Be[�+	�UL�үۖ).7\�r�$h�0�]J�޷2��#D�%P�7\�f"�(�S7hY�zv*�
chҰ�-P���73�k�"�1^�*�.����԰�N���.Ad-�w.]�D\Y�[���(�!*C:�I�m�d�Wf�+������A�w���B��!�������"S&�3�ŗHPB��z$�3�m��15��]��� Tk2	b�ŋHQ<�6���k^~���I�(�i#�*
���E]c��7�z��[�S,�:^R�X�U����%��wj�Ս�hY0!*$Db�F�`ն1��&���֞������%7�bމ�zq����f���7k)�Z)
��o��ňE�Vm�SA��+	=okwL�/H�wM+�j"1�jD~�y�Hˢ2\��.���(����O����E�a�m�����l"3lm&��݅0[�ƿ'0�,!Q,*Q��d6Y$R�Q����S��B�QzʙYM+�&�͔����<ӗJ�Mʷ���7&]:mHfmfU���F�+6n��#V���X*۴C�V����L��j�45��Z����y���[�&�e,��Qm��w�,�7����i,Ӻ�*����k5lK���bEhKv��t ����V��#*�v�@s�h��s�����,��z�i1[	ۉ;����o4��Y�e�#G%nc[����oX՗#oj�_�h٤�;���e�m֊�Uy�͜�w��=CZ)�1��8��UU�����&x$3��z+)��s7�m�ʸ�mᲨy������ԝ؍T�4i��5�shl4�!�Ow� �h�^l:�X�D�����{n�{i�y�u�f*�5�B�^ʄk��F��N���,����*Xwp�I�Y�D��d,��j�ԣ������X�{07��V@z賸�L�g��/ n���,�4Q�x���Q�oKK�&m��R*x����(���ԯhV����$��f� 4�Ճ�֖�}�.]u&�t��4�����;�n{�J	�EAs(T4Y���K�* ���������x�IKD)\�j�e��bW~E���$euX��ݗ�ų��I�Ǚ���Pώ�ћ�B���U�M/R��ZyÂ\��3Z��C/	`��{)�se��(ײL�=2��
�`eV��
�A��0�%��|Ȫ��_{����������U>�����P;��Ց6�qq�&�.[�G�s�5r��qը�<��hk�ӈ%����M_;ڮ]��d1Xh����є]r]*=.8�
�ZBU*v8[5Bg=[��'"�3֝�6�_�z�����h���sh�łz�6z�ٵ[exŇjN���ֱ7�M�۔�9���3P���U�d�,��Ҋ���.�.e��:��5{f[����H�X���^N;P4fu!�{��5��A,�,��\�8E��C*&�lw�+�@�73��(��SK��:�[���2�n44]��F5�:�וh�0>
�.�+T�{�2m��ˮ���!^4�� �m!�H~I8���Cm̰     �ml���     �m��  4�d$�bD"�2�  �`!��� H              �� !l� Ā�`6�  �)M�	�4o�g+�E�}T��0򠘽i�K�mڙFI�f-��CO�.��H�p�{�NkV�:�dPoa��X�]�R�6��{?�P�mP�[r�	�6�l  �I�2�AJ i0�0$
Q)�3�|�R��ˮ��l����7���znj��Y�0]ӧ�ؙ���iu��P�BϜa�P���@���P�0�A{B�פ��f0\�'Ɯxe`B�ʕI�A]E�d�����Z#��Q��#�
��/�.LrWzw��	ҝ�"s��L��Ñ�����ԭ�ud��z����=u(\�L�
����:��t�R�v��v��Q��8㚠]�US+d0�� {�� ���,�t��j}��h�A�����2�^FD��BJ�f�CI�C l������  $BD� ��rBW\��5G	-�ʅZ��gnd�BhV9j<��ݗ��K.��Q*5&X�D��"�9��.�������� � �	�I�BLa'Y 4� 1�I�H
BN��� �$��$� mH�Bz��I�H "�!�� ��L�� ��$4����E�� �I��@%HM$�a���`Cl�i�y߷���t����E�E��Db���TFTY���b(�ETbR�x�Df�b�"�"",UQE�""�n⊪$UX#Mb��EQ"����* �UU�(*
��EDQFE�F,QQ�iE�U��X��0�Ҋ����,�����
�"�U�UH��*,EV
%3�bDL�n���1� ���<�F*��EEMШ��TDATH��b����Z*�d�Q"�.s�M*"�* ��eb&ڊE�,X��$MR�H�2�DTQEQV0EUE�����b�i�EQPV *1�e��L�b��ыD��Eb�"(���þ�(�PX" �E�"�ڌb�""
*��)�e=h�,M�"(��,TQ���F"��X""F*6�Ŋ�DQ��QUSL�"�cOXQb"���(*�EDH�88���LAA�?!S���v�*��(�#DkY�=5���y����U���
�U4�QE�UADX���*�"���%b����F0Fj�'i`*���TTDUUDDH���(���Q�
�uۈ��
��X�����kJi*$F"�AcZ�Y�XŌ`�iSI_�f"�
��1��Q� ���PQF"�e�Q�+2�X��iES�"�(�(�V� � ��LQM�Pv�b�#"�
�EU�"����L�* �*#P�|�DQQQ��b"�k�`���YAQ�A��c�&aT����E"�ڎ5UT��� ~�+�/έ:�@�=z�M�J�D0�S�a�YX�QF
"�q%UDE�|�"��EU���Q]�Q��E+}��H���i*��PTDݪ��O7qAbj��ً�t�EDZ���e,��DϽ�5b
 ��ʫˋ,+}����Wj�zo0ݪ$D`����b�Ҏ��QA��h���b��(�c�]�����0QADW2��;҉UU]4դ����"#��m�>�������k(�W�
,UPT����G�V,�T`�����ʊ���_)�US��j�m�J��("
_.F1QQ8�f������mU�h�0ED���Q�,��][cj�����"���at���V����5j2�����(1��l�f5�b[b,V/m��ߘsuX�m�� �� ��c��z���l��
�#�{���b��_y�a�f,f�����!����x�����i/�QE�t�TV"N7)U��/�x��U�sJ��3#rʊ�-=֦��U����V&���ڊ#Q`#�	Z(��q�E9e1�����v�Y�@a@}1ZY�^7oJu'cF��4E=���5k֬c�E�VT���Ҍ|�b
�U����;�1�T[=�(��Y�y�{����E�u��}�dģ���X��Z�}����O)Q����;�,r����׺3)E�ֳ�
��G�ք]S�3(�}�<u��GK;�ݮ����,XɄ�@|�1L˓)q��6/�Gw�ݦEQJ��3T��U��**��P��ȳ(��4TE<�kUOis�b�DEU����J嗯�M2�5��W�̬<�4��T���HVЮcmr^ѥ# p��7����Ѽ��R�A�%e��|�9a���A��֢������k�oL�Ȩ�W.�,U�������-TM�e�oۂ��޳�`ĩEj��e�0W�uC���p���)��i�d�C���h����|g��2�2�<�Aɝ!
� f���i�T�U�k�S横�������+�EE����P�ٔ�{J�Jt���X��إoߵ��֎DG��bL���z����q��s�mؖ���n����@���q���L����}=i�
-�.�����/(8S��y\�˝�6�k���J��I�t�yw�J�;�"�[�F{x�����JӖa��ۮ�8e�%YE�^a�kY�<���w�E��b��h�ש�r�k1���C9M��c���i���#k�L��p���J�1���lO���+�J�Ʒ.**��L|@����֡��(x��Z,;jgy��c<d�Y�F%o)X����u���1+nmo���������a1�_|����~B�P-���~=�㢳z�Q�iPQ���H_��;}�Lt�V}o*_���Y�2�&Aϳ2ʪ ����ł(�R߭��z�r� �RVG�}�P6�#$2����Л�d���.rr����w�B�K�%�Uo:Z:��SP�h9�'-5Z�J�"��U�{�9h"��_)X�b���i
��(e��Dm���g��}�w��N&ae�oٴh>f�I2�qy�S�1̗E�o�}��0r�'�=ʑ�殍-(ʞ&0�Ϸ�u�+��Jy��4�mTơ�l��8����8���SN튥H�A��Y�t+%<�S��ݵ@[�.J����q�� "��!��0�����)Lb{����I}�6�'3	�YMZi�߷�y��Lg=~u��4����N�;�0��+7�SHV9��~�IZ�;�i�[IZԨWϮ�����]_m�WWc�1�t=���`����s�L�j�5~�&4�J��Ž�Fe���o�k۶/�hņ�6�}��>�N;�꘼hu��J0��"�ZN�uF0�Y#~�k7�6����S:���H��PF{���{gÍƑ|s�:�66�Z�¿^eE�~�f�f$��8g�lެ����Ӌ�{o�M�ں�-��|��־��mK�Ǻ��!��z"�����*��_T�T1�^G�<�L��sE{f]��6��3iY�e��7�<Bh�D̾:E1���R�{N:�2�u�����E~f8��~�x醒�˙���}�8�J6��~39-�j�a�J�^>�Ks��H�-��6�wL��ٷh��S�5:y���R�q�3%5q�Cl�_��t�<ޱ>�!�iS�'̾P�5���p�ۘш�IĆ�܀c&*O�Ro>����~�]����4@�o�'�u��S��ai�u�}�L�ְ+��v�\əW�u�����|,XcR����2��r{��i�J�R���޼׃MܪX�zCpd�S-��k��Z�"�M��u�{'Hfn�Va|O:N��g�S̤�Q��P4 �lj��q���mOWv��7�2�	�Ky�	z�s���\T�ֵ��.�UZy��0Ì\�Y��e����x�Sf��bDc\��O8��<����̧\�l6�n�2k��*�8�3�SGrT��J́��`�2�S�d�"�
|�@�,ي�y�=�k25�o���g��6���wzL���w#@u/�W�p(�0�4)̀݇F�l|�&�մ������"x��hj>ˬ��+�]�;o]Q�K�O{�`H�$UʏjPD���C��t���VkW���E}{�c�~���w�
Z&���^���{�$/���DE�D�U1$�(W%,VǾ~�|�c�8����}I�1�3�K��)��ͣ�\J�~�f&�2��v�4����g����n��Fn��u�����l<72�gq^ݹ�I�ݝ�t�`E�W���u_`ں.�7AĶ����5�L�f_�
�ŷ�l<f�n& c�J�l���Ǯsߵ�-����F)#r��(ƨW�a7.q-ʁ�3���*���}E{ø���: Ua�{���;��kU4T��s��Z���[��z���ݳ}�h�i�˽\��D@G��A�C5�<��	�<��߽���s��dU��5��N&�Rhת�}W���F�X��
�bm�3��a���J`>�]�i��Gd���=^Z�Kbs��_a�s��U��٥^�Cw�K�T��[�je�@�8�����&����s�Ц��&�%��a߯�3)�vsZ�3�i�4�՜k>��(�uBl(9�q�z��  �XaU��B�R�M��~���W��ī ����I��� >����B&-�R4Dx!22���A��u�a7<>�!#�R0D�=t7Xe>�����h�\2]5�Tۮ}�hi�}�缘ȧɦ���:oM�@U��
�	�����8�V����34���H�9h�}l.�z`:k�>��2a2�32"E�(�	j�v��r鋙Æ��z�|y`�ݚx���Ajt�r�u�.�R�O*|���k��'4r�=�ל&���-���SW.�'�w�켢���}}v�Ix������W��2�0�T4�y��bc�����l����u�Vl��]�l���႑�3ep���MS~�6�����}<QJP��~UUO�@.�����kn>:cmVG^��Xm�k-��h���c�k�t�r�Hh��`;���W�f�9oڣ�͖Q���j�r���ҢZ�|����bfT6�ff��њfZ���hGN�rW��P�DeI&�X5��[�w��H>�DT�u�j���j˶n_Hf�!�������%�&\�����w��%�FhYv�_'��G̚Hq�d���r������g饳��l��>��B>h_7�hк��WuD	gj��|+��R�>IVW�GNo�ru��x�5]�f�hŊT�ɏ�&W��l�5�w{MaH����ϼ��U���ݙ�&�����mB>ԇ]����:5���B��z���-��l�Ɉ�����"T -Y9}Ɏ�K�
z���{��ۙ���S3�}�O~󈋤r˕�W�̕�A�a�։>X3���_�hL�2D�������p�[W̐�����(L/���� �>�F��0;*�ڸ���I\�}�:�w��|��n�5o������e��[3�z͍'p&�r�+UUU������h�k2��k4h9q)�$��ܖ���&rv�0��!��X�0��^F	�Q�ܘ����kL�	�p�,�dd�+놆!<_<����������2���Y�*��I	|���j�$M.5!wQ�����8:��\���pթ�j��
�F ��u��5��2�m�k
�c`����fv��⸏�z���7uMg��{�%�1���d���6�[c��$�C`  �D� Cm�2@�H\a��f֔�&gdi)�ʘ�r�tT�6#me�Aġ�
s�l=w'?�x��)Dp�>c��#�f��h��B	��vg�r`(�P�L�1e�K���_2O��Ԑ=|2	q�Bս,���P�9u�oJL�W�� �PQ%�H��:PB�1m* �-�Lѻ?)��2�
D2�O��T�j���L\ueoӯ�>��I�3N��~�4f�؆y�~����1�4�2z-@�xx#�d�Ѻ�7QB��uj�pwn��X2���2�BkO��> c��֙��%�r)�5������}�����t���f��*���
��V脌�b�A�$��5J�.��y�|���Vr��ύ���@R��Fa2�qBz�Zgd���J�:�WE��Y��O����������~�D��nJ�z֮Zi�b�,/d	�
�Z2!�Ptm1��A�\��0��ht&&0�}l�����6:|��*�}��fF^<�ݡLѢ�8�"��]۪�zS5�ڡr���	2�4�?WMD�0�RV�nV�ʀY����2�熢�RF1ؿ�dM���#�!}d���d�.��m����B+&T�Of�Qtʦ)�?�߲'�wC���@Щf�&�S��3Ƭ/�Z����
\����9�z��|2N(�"\���k+��0Q��8mV�m��E�=H:z�^/�(v� u��㞼� �//o��S��\�����A�E�(с	�I���La�(J����^v�k�;�;4m��n.S汣�zwN�Q�o�o7+�n��7}���k���|[��R@!�C�,�N2�� J�� ~HK��!�'�Ehz�!Ԓ q��+��[Մ�� T%d� @�7��׌�Hڤ���w�| ���d � :�!XH!�d		Ϩ6����A 9�I��'�$������S>�̷~�v��Z�G]憲)���s猳�4V�|-���h�c��Q�@�S��o�M����J��4�z��D�ۯ�2v�f9�቉ycw��w+�<2���Ø����5�mD�zR�0�U���O':nE��;��p�x��2�9b���W@�]m�=�`��|
V.�L��d��+�:��Y@��G���y�݋M�;(k�^�����y�����%b��M���>������hD�5�KB�J������n��$�ȧ�Eg�X��ӱN����^�֕�!�s��fu��3]�B�ck���HO�F	-J����AO���h%ě��&nP�/�:�Y����m
hx#Tk�&+&6L`�e�S�v���&�.Ή��_@о�1�CL�q���ų��n=2�-�Tz�Y��<��4!���
'���	Q2�Y"���Dp�A�ԧ�hS�V�31h@����#�!:���w˛��ο^\��n[E�d�wJ2�מO�q���J�c�fw+&�D��1�$$��D�bty�� �x�Zb�Z%J���:Z�΢�j���f/�zGK4�%�D�e�=�!�$��q64��*����[�;���>u�_\]h1:݊��ά���C弳_�V��ˇ�����3����.���L�*'�ږ@�y�x%��r@Cs;��������,�w��5�����י�zl`�:DiKRa|uC��}��{O^�=d@fX� QwJǢ�,��t�Y�E$�ֹ���w,�5���6�@)O})O=d��ר�}G}J"u����+����I~�V�w&{ָ�ƹ@$-��	���$>��ܚ����!���S�'��� ݲ �}�	'�����ڪ����`�;��R�K|p�ՈJ��5��a
�ʹ�iCkwy�ʢ��H�y4�C�IV��d�=�R�ӹk�bK��\��g�{(��4�B�-oc\�Hg���]5���"����R��]�슺��Wk���y�|���s@�ht.��2�n個����p�5�:-�sQ��&g�&^1�T&��<�"�{��f0Ο���$�����-�+r^� �t��~��P�Ʉn����m���"����2��S���n;x����TK�h�ڥ$��ZAZ �	��ϐ��˙�uD&p�&��+��25��Z5�wT�8f
>�Q����ZULB� ѕS�쬻s�&be+�U�KA�<�0�樱�xY2�%u�2�X�wk�.���I&�k����O�˫S���l�r��/(�ގf����	7 DjYT�(F��_,�oiE+�˧���%c	��ҽ�I��]5�l��5��'�W������ӭ@j�!���Ʉ�Juxw[�Z��[7"�L��U{�J��@�߇1:�fZ�\��Ӕ~  -BN�yy�)L� � �����TE'�7C���J��x�y`���6�EK�8~b�f@�u��w٫�)-kK(�Lzq����`3�O�3��#�3�7��ꉱe�y�n]|�QQ� ��Kbb�ޭL�,AB�:��ڔ�1b@���-Qz��P���:>c�E�-"�U��P�+ܡ�)�y�6_�8\l#�bꮮu�M�ޏ�^��m��/���yf�wD�
8��,������U��ۛ���6�I��&�,�ӭ�����ټҎ:���.�w�:�ۏ9@WD����gl��+%�w��78,�G��r\��Smŋ�d�,�
E"�e>�7���Ć�?N)�;�埢BWԀmVŠ@���7�q����.L$cQ3��M\�x(�OVϗ�wU(BHN�;�Wښ����P�:��u��{�F�p� ۄ������	�ZZ���)3��)I� )vȨ��|�A�>��M�eC ���.'�9���x���I���4�4k����s9�[|���[a���X�u�ј��}���O�Ǘ�l=ߦsރ�	<� �?(v��?x�S��H��>L��S�JJ]}�ߨ����\��,�D�W�V�h�켪�wx*��7�!��۩�9���>u|I��?����U�;�,�#n�P�B<��Y3&R[=��Q�{,
M�"y�CF|H��m��e�$m��&e=�:՛� ̙����.���O1�{
q�ZX����F�
�`7��u�)�����:��!�9�$�2�9wn�Qջ�}���
���
Qk�_WuN�ְ��_qt?ŻJ�.���
g�kf�e�i�7N���Z�-g~(U.\c�-˛�%���z65E��U�a�W�+lGGn�,CM�
BFX`�{䐫&wv���Y	����snڌ��d��UU����T����L�*�����o��U�I�cz�[ݦ��ۻa�M���(jxS1ВDnf���f@��$�e��` $�����*��   �L�6�h]��SP�ח)HA��!�K��g�J�^�;�2t3󽢚�`H�9���e:뵮>xksO�����NL9�?=�"%�����TƘ�P��I��7�5��R��7���螼�x2��h�}l&�K��>�mX��{�B�a�O
�
�m)GBS%�k'ٵK^{5�:����Wt�s��hEe%��{^��vt��*��k�Hd�reJv��z�?%M0�� �y�ȴ���k�B���l-S��˹&f<'֟�#�%~�ې]�P�<��Vf�Y�"��L�Z!阀 �[,B�F(	��,<�MC4l�<�*#E&_�V0LL%r�S\��2]n��\ms�u��Kmwy!7I�2p��r~���M}wHҌ@��r��6\Ln�aLP��f݌���^5�쎺i��T��'n�\��1w]�� �_I�������/��"?B-�0�1_���Qy7P����*�6#5���2���Spa_ �z��EBof5��yB�S:l���k���*��ӡ�F��
�{�["2��]�niG,p�X��*t{��^��|�a�f�e,:�B1�]4�r�W+����vz�B�T�t̷+y�k���2������8�O۩*�]C�A�Vn��*�=��W���^@�L\��gL_������gq̥�t�Q$����ۆ'��8 �n ��䉗W!�d֧�Y��	[�]�b�O ;8,gWB���ۗg$����ن�J���ݒ�n��9�y�'bp�T9%o��T�{B�.r����粠)�m�6w��Q�D"]�쏕1���e�X�D��VӺ�ْ5n� d`Yf�L���>37r�==��W����2%�T2��x�@V��H[F���I�V�'k����V���ٱj�0������)�t<��Å��k
��|ފd֎.��x/+�^Պ����~�1�f����j�.���������b�mL�Ι�_�V)V��-nw̥�"+��sR��A��^�;�4���x��wm
�XeR?�1�	x���ǐO�pܞFX|2��1ۺ\��?)�a�,�:X��Γ{>纨K�āt0����%������Ӆ����.�D^��&��>��ܾ�A}N�����11�:v��YX2�ً�`�to�D"��?M!LD�-���ؤ\�=d���'���S�9�S��2��}�4���V�'�/6��׌&f�(V��������T�G<�i��F�l�\L
v�
w>�s��SX�B鰦I�S��H'Z��'��~_Os��|����]묆�N���f�[�`��D���v����~wҤN4v����n�L5D���/�(��!����A_�2HG/��c��Sgϳ;w4E�; �뷌�b�9�3F�����U���Ƈ��J��68��3�0����N�rl�ɭ�����z�L�i��r��5�cB��vz�x�Q�i��g�^��=^%�a�(��@H�"$D�w��_E�1���^�4U�
��@ΧٔY�+�+:�߼hvi�+����ĩ�߶�&�����P��� F�tj\>��"�����ýl��|�YHȆ>�)j(}3K7LJB�a!���Z�+��UGF���v������w�>�{��]r�{���7�"�Ϭ����ݡ�ҧ�%()��1eio ��v�^�^����)h��|����]/��co��B�+���hK��&���{ߢ�D���Ez���f/�o8�Í����w}�s���l�%j�������x�x�1��5Mg���~��s�_�x���tNZ�I�e���V��6+�����X��Su��2�P:�93�:h_3BhU'��F;�.�%3P!G�p���JD	ipV�6������i~��4��'P�{��I��(6F�Cr�(E�	�!;��u�A3��h~}ʻ�^m^z{������v7!Q��N��V	٩u`��nKt�{�՜͏N�5�}� �<=V���t�K�c�VW&�Cuq�Mu]��M�u�8�Z �,r&��������Z��捝����:>(���^[��)V3�١ŧ�Z*���d�P�e��s�d1�oe��U���m$�d�5����śٰ��5\֔�����)Ն�$�x���sa���gW�G,oo��x������Ob����1��%�E��s-q��d�1hY�wpc��G{��.&��5Q���K���S*�ϓ}�1�]f�f�Y���}x��:��؃71�>Ճ�OsE*4��G�oj�I��)�Yy��\����]�������zc����m~���pBaV�D�t���ls�iZ;��_�N�1�pU�:�՚3�Ѥ��Tǁ���L���݁�4V8.�>;����G5]<Xop��lQ7TU�y�������:n�LO�E��
�����x�#��-��fbE��Z��D�iu��{�>�AF��n���TФqk�V�kfn��`�As}}� ���nľ�͚X����⁤+e�����ڥI��o��qF��滒������b����*����=�>K��T?�^�4�I��k�y�g�aY=���?{�i�Y18��f&�"8���!�9���~LM!�9����,�uĬ�pϰ�R�g��1�ߟ�:�<I���y����������W��^Ö����V�Ds3Z�L�78����<IQc�h}��5�i�a�N��iP�pgS�޷�{z�T�>x��w�u��+�Y�<9����6�!�`��E��T��Y�h៴m�u�T���w��]��s-���v��_���|���g�*`�C��� ��}�㷉�1�ߵ_���'S�L�F����kv����vy��y�H(��!Y�Nk�6�V\�[w��M\��لY��	���ՆٗY��#G�V�\�" ��=�F���f�va����O�DxG�D��AF#��H�&i��k�}��N}uR8��F}x�n�$��Y���:D��<��O����\h�����.��
¦��k~�}��+
�eg��i��! G��^\n�
[�z�*�����2��"*j5�>�Y�",O>�n�;f�W�c�?&�ІS2��oGۚ}u�f٤mZצ���Q��E�z�34R)������I����f��Xgl��XWI�5��rbq�C�._������6��|�����-��/�M:΅�DxT��D	�S |!�<˧�1����I�Hs)Q�������M&ޥיF�/����J$�g��y�����)�Q�����Y1�\g���8�O�P�M>�~����YǉS��y�y�y5�d��S'����WB�`�`
�����{��fҥF�[G|�D���`+�D�^]3V]�˩�Gt�?&�>;g�s<׻�{�%M!PuK�J9a*c8�zͻO���VdNa��1��a?2z̏��� ���Uuql,��z奚ߺ������E�)l����v;C����4~}q���fj�4��0
��_Y�)����u�O�S���bj���oe� ��!��z̨iD*OY��wˣ�k�M��:q�??0��B�6K�@>�9���n�]�_Bl�cD��+�Ϸ��`��_�>��eO�1��1�&_���^���C����g�����bͥH��S�L�k���w�m�~q��g߽����yb��g�q�c����bÏڦ�c�S�AIޣ[s�s��b���P�\�Ο�|�&�C�nfi���P���k��*)P���O�����*������\~LAK�f$ӈS�b����6iM���5��}ϐ��x�ˈ9�g5dĕ1��������""ʏ���]+Q�.> ʬ�§G��pݷ�6ߐ�{Qj{%�r�=%4ƕ�Z�s����e�vun�� ���r-���`Z9��g\��ǳ�_@���nx�;f�GH�<h�ǝ*T,��ă���}������'�oSl���c�3�|�7��'�k)��\¡�+*��Ⱦj�0��
~�M�ٿ��b(�g��`��X>ٌ���~k��i����;��>�W�o���y��i0��͞ݸ�����[%Ad�� i�j'n�Tua=C|��5I�P�a�bxg�i!�QE�1�
"�" �1�3Z������6[;g1�C��<�,�I(3
~$"�|���у��|8���=�E�*,����x���k�8�n�6�5�@i�6��Y���i�E���p��1���+�x���8�S��>p8��v��Ѕb��R�g�c��{a���iXbl����3=��������|�>]�.8�樉�4������%1��O7�I��ͤ��c���O9��4�`��3�{�|�N�q3�*w>��}s�I�J��y��w�������}��Xbqhn����d��@�J�P�x��+i�A;"��5�z{M Vq�f:��d_���0~B��*M��C���n�ީ�4��ֺ�3)�G��~����J���'���;_,4���'{��5|C�I��7����h�$�1'�LC5�����5�k_������\fr�Hc��dֵ��Oɴ��w��w��°4��%O?Rq4��ԕ��B��>���bm3Vz����7`b��"�.6���'�_��q�tΥݚLI�c7�o�_�����&C��o>_35�_3C=
�etԜ��Ye|��?2lq�����ٴؑ�q�i�'r�jd��gp���'<)Re�D��FR��10jT)�Z��G�f�N�s_W��r��C��ֵ(��� G�\$G^Ӡ8����/��?��I�R)���Y1*Myt!��&����SHq��M�1a���6�3��bJ���W�>f1���+�3/~֢��q��o�翜�:�k�3�چ	��z����w���Y�������lx}�D�/� D*0�~ú�J�γ�_~��8â-K��D2�RT*Lq翹�u�N]!���\�F}`w.0+��+��g�o���
�R{^_�?8�|'M�>�s}����0�/�YdǦ���=��gn�f�{��x�Ԭ�~��8���,�6^��a�8����I��!��5�/�~С�m�n��"����YX���o�x�^�~z0؁Z�s��!��Y����Ղ�4Ut�j��x��:��VZn�ݭ
�/�H�0<�=x6h�G��~T1��3ijЩ��aq�G@W!#��&�F�"��?6��)�jdd���a�hT��5��ݲ�Y`]�s1�0  � %�r��!$r�8㪮���A�BI$Bet�3���3*4�;p�}��?�Էfv�M������<6:D��u��X3���~�>�v��S���L4]`\�e�X������I���01��wWI�Syx�"�a�<�\Z���
E���LI���O�p�5��cAO],g���_iSs������un�رv��F#��`0Gл�M�� ��Ր�fx�f!�F��3c|̓�FlϳI���>�������q,��[��Debc�A���O�Lq����b�L�`����˰")�� 8DH�B4�o���U��]|�ҋ'r����7,����)��Xm��8�P����I�.�_>���'�ၦ)+Z�8��V��i��)���*Aa����4��+�g��^ V��o����,�IMr��϶_�]BP���
����6�&&�_<6<� b6��'���Ĩ,P�=7�z͢��\C��gm'���3�l���m�X,�*[�!��G��8����-���g�1�4�w���IY�Q���斴Sg��v;�/�����B8��T�� !j}�i4�P����t�o��`}��5�r>Xma��L���1<|v�]����OSmVW9��6��7�~�b�����W�0�qP�T�Ki
��?�����>�*���w�|N�'SBT+jU�k�:�����wg����~�iĬ]2������:���d�S��٤��V~a���6ͧ�T�o�M��其FsFd4Τ�WIZ����}"�B3�7ܔ���]���" �>٤D>O7@����d+���H��>�.��J�Rq/�o*h�
B߳ӝ�u8ì1���ۡ��bb"�4��0ĝB��_�M$ݲy�s��~�EN���y}׿gO�`���\�w��n�}a�P��M����
��k��p�h#6��"�l{����_�=f8�wFEơ����I��y���R?Z�bg���f �S��Z�ưX���m��L�+��3�Ѵ6����#ۯ0;��(�2T�w6oO�zw�Ï��l��nP�O�I��6�IѬ�Vz�5����g�IuE�5Hy��;L�I����y�B��vL~�h�0�?!ׯ�����0ǉ:����D>����mVt[���>�#�>!#u���v���GP��V?�a]3�)��OkV�Е��*
�����V��{��+�(�}���L4��h���Hc��|�b���?/�B#����0V���C͙�>���w��ge*./��	�Z�%=�N�{�Έ�Ͷ�z ��Z�*j���#s���[Aݓ�u�+[�F���xf���m�W�xʄn�E���1�d���\�C�l��O^k[�X��W�8DA>��d@����	
��߾�;��Hi�ݥL�if�M$4���s�o+���=�4�=M3�E�����M:f�z��?g�Fӛ�8��_~ɮYR�eF��wF ��Q����o��(c�Խ�{E4��۶-��z��R>gy�k���z��Q�_��/���=q�M��4M���ݺO���u���8�*E5�ZM/�1��_�aS�����!�17�̜f�s!׻�t��XB8!<�eYX�i��Mّ]yX�R��M�qM��߷l3(bbw��ӎ�L�m1?=r�DH�8�C��06����fwXm?3��]n��a�K& ���O�r�әI�q���������2��h{�:�3�ƿ0�W,r��~>���s�g�Ⴟ2i�q'�7O�8��&��{�!�QdwJ�fH�:���皕:�}�t�%՝=�9���:��\����� q�;��:I�ۈ�|kl
����G���&��F������n��x������ǟYW�&&8�i�{J��R���� ���I�ӌ4�g�in�
�pq��]���8�ͤr��k$�N=�"�3�Z8Ņ�=a�]=���4�'�q�tf�h�3�+&3o���H��c�>��q�T���\w^��̽Sɨ�]R���C�1�� *�V
>6��Ӊ��y~C����������TG0��h�ɤ��vi�O��ͤmơ��̚��t�S2��c�Gv�@�eiSl3�L}��l�)sfqB�Cbfg��Κ����뮗�[&��5�]?�|��K��i�&��Wd��ٴ/�o�m��S��/В��Y����i��m���i�vE�;�
�u��SHx����7�u��YE���%L�6�t����D��rc�"ݘ� Q����o^��Nk���-��+1;h�Z'�(@W���A%4�f��[^� �`4��=9��ۺR�ݵur��QȄY~��b��N���O'��w3$@u���R�W}gT���H�LVD��Uҧ��wKrp�F$h;=3fB'jB�:�1^a������v�/:�%,�
��ۣ���0��(��-<=w3y����&�3��:���јw�����_;�{Q<��oG���R.鶁�_�t'�߶�;�nW�˹Bƭ�,�n����J<�A�O"9>���$�����ڋ���_����9����N|�V���L�2wjjM���KJ>���+���#�y������ڊ�B�^q�lê�/.�h�Nv�__��I\i194(��4�X�$[�*�CئkLp���o�j��.���:��vS�'���vOY�(ޕ<��x�f��A����3S�ự���6.����;��.ݬ��uL�5[T�I��&��*0�R��TUR
�`"�궭�c>��L/�ŕG�M�
g�TҘ�
���͛
�Chө�o>i��zt�y}b5�3<���ŷ�k�j����F�R8�fd��%0�\Ē�!�3I%S*�O�w��1������wtr.n�j��������R�&u��X��_�߫(B�AM��`�����}V��Kl�S�A?=k�+�G�	�UMfGPMm]�摤 ��'&yLb��)��E�%�(�j�i7����D9��y�N;|:Y���f�U��C1�J���F�*k���PlQ�I
W�h��*m*,Z�҇�e���07��>s����FU]�K�E��J2��(ߝ�(���M�3�c�pW�5��^5V斷1��F[r��{+��8C��m�Uo�߅nZn̯�[p<m!k��q��5hp��c�I�����8�t}�[*{
�4���<�}��%�]>��.q�%w:��ژ*^�{b�{�M(	�N�<2=��RG%��r�O,G�vTě@a�����NPCM��m��z�r�%�鮤��~.����.�N��y)�b�ґ9W(۩�)��U\Yٯv�^wh.��g}]`��֘n֎N�=}ޝ����qB ��������,VP'#Ԫ��e���b�[Fk�lЍH��ylJ3�¥���b"��>\�-y,)�ԢZuxPc����?I�k*�E������ayj3����U�����j���B���S9�m��tRۺ��T��5D�5�閲Tw�SkV���H�H	2D	�!{mM��;�S��݇���[D��H�
}�ڛ#L����i.�W��ߒ������G]�.)���B�!�&68���w쪽�<����ۏ�^de7�E9X��&�_7��B�޵�B�9RVc�#&���3t�B��W�oSX���'q��󨝞�����O���X'���5�Ȝ<�o�Q^*)_h��t����I��R�$��Gu���]�Mz��x�eH�k^��}1&{}�{&����H)�Q�%S�wk�|��#����Dp�/�	�e(�}E���[�6��|$K/]�.J�}2���^���F�К��n�7Y�UR��+�p@�b����X��1>䑻\ʘ�jm0%]K�H.�I�9��� E���z�Q�;a�O��iz���V�YK��iT���83Ջ+ի�}�+#��Bڍn��^M�3�X�9��j�[wG���}q�"�oh��gڦh�US;ٓ��k��y�g{���I��2�>� p�Ϛ��y�?�t��|L�P�].���f��A01$*��ձ�v-n����uR��~�AO��2L��$����|~΍W��v�h��9V܌�փ�ta���.��:�Fk49Ɵ5���n�#WtP���rՔr�����i���ݪ7���m��6�4�$�  -��!���d�$�l�[#�r{�Z���D��{�e#)����)ݽs-v
0��:	�F�Âp�I���?��)�'bJ
;����(�N7�������d?z�B�v�D;��v�d�����,U����6Yo_���/Q	�G:�hU^���+�=t�~3�R"�A,��T�dy���Q��FO�9U�Wi/� �/���s���A�����&��t�� ���D�g������,�pqQ�d�z��,vx|p�+��2���c�&> F��Y��o�ϚJ���B�)�X	Q7���C{D)��"$@�Hj��@����}~�X4a����`/$#�칫����^��xH=�5f�̘:��46��9.��v���Z��<4���{G�P՚v6��R�f*t ܝ�7q;�m��.z�*����b,����)`�c��#R��7�J�b��Q|�W�s��L+��t	{=l�u�|�����SW�s��R!#
��@�L��C;F�︌�ŎLOs�&jmFS�`�y�+�QP7�Y���:==ty+MB���_�F{.����aC%�3T?g�wq19�3ɼ�P%z��$UV�r�V �`4���;pjxl��K���H�R��v]�;�.ov�DRT�%ur\�hQ��zq�]}o�*)X�bs�xL%�~<�OMR�P:��)�w� �fjLf�$��򐰔x(A��������$uG��(d�ttÕ�m����Q�g�䦝���N�����u/��ҭ���#vrGx';��:���y�gC,Cq6��\K
[pD�8֐�*�CP2h������8L'rD��y�{@���yx޾Ⰶ�M���D��ה����Dg>�D�պ���F.���H��y��u�M�	����&%f�|9�'��$�c�H�O� �j��Yi�kǾ��7n�~��	��E�-�U.��Ή{�M��)�z�g��4JS���w��A�0�Uv�u��d=)����M���U׊���+��t_J��ު��k�j��a�)z�<��":��.K���*���՞E����sRF�>�Y�%�*�t������v������:9���#��j�*I	h�L"����*���uG�NCC��G�0`C�y^��oӾpW�_�7�5��ڽ��'�6.���)���O:����5�A�u\c&f�֤��H��S_6�r�5n8�ҕv��zK^٪&�������ۜ2���_�(>P`�ZD�I�]�q�t��]���Ya�o�g�MVl%qG�)GI$����������A�����jNqR��A-Z��
>���F�Y��׎a_��Tpn�PԲ����ol���c�[���׍��0�`�c���qS+m�:>���uRuL�|%@�����ɽ�v���so��EI5AE#�϶2�-V�Mj*��<�%ںL�.`��c����}��'kBT���렘��l��F��4���;n]l"������33�ȫ�J�-p�-;�^^̯�{�̊�}u�W�r�[c��-�J����9\��iY�g��?�c�m�����E��<��N�K�(	dޝ��Y�<�[��]t�:���=)
�l���J�89�i9JU��ɚsV���t��8�J���mӮ�
�g"D4Ùu${lՔ�]����Y�2i�<W���dH>]�ͦ%t���b�,���8昰	?W(�8���*4�9��O�g5�y�\p�W�OR�1��>����7�Np��s.���?�Dp�׫�F�o���p}��H�6008ϵB�R;�{�z9 £���
T������d�_���jI�Uwj� �8
��M�^]L��Ǧp�|h��������������1�kB&3�R���@�_�pK0��;4�U�_�D?]Wړ���J�sQҸZ&h�
�9�ؔ�H�l�H���
ӭj{��}�:��cj%�x��&2�ˀL��qh��)!v:�ύ���?v�۩�Ϩ&��ǳ�fNʥ4�V���֏)g�����!!x�˒�6&$	93�����LP~���/�p�V��+v�ݡ��~;�p�nΛfh�6LS�Q��T���^���?h$P�l���E}5�|��@��3=��Nu���	D���v+����i�3�_<��AȒm��I#�Q�u,+�L!�F6�r3ME���P}�&{�2� ��$u	�*�Dq��]�6���Fu\z��r��2Są��؟z�J�b�NGfWB�X�����&�ߒ~���|x�Q��a�b���p��qB�w^u�&�晑Yw`;���$7]���{	���M��"�a0�.c.O?f�EŠJzU�l$5����t0q'Yܧ����4-��i�jJEe�!��f=�4���a����m���j� �E�p�;��8'|eR�c�Ǯ�E��f�I�#L�����v.W�u�@����.T�
f���ꡧ�b��l��[���(�q��vM��H!|F;��J�Cz�}�[����S*�N�E�b�'~tz�p�:��>��cY���h�V����E��)J�J^y1bh	�.�:o�:I�X�3b�kq*��	��-N�tUH(<���_�TKt�n'�:��(v�<�j��/뫚v�Da=���!�g*ǃ�ws�9�w�"%��ۏ7x|V��[K�qU�-�iw~��?��T�.g8]B6�z�d�Rӽ}'ڣ"N#R �֤1�J	lf~�A��1��}�ө^?�N�={Y�Ws97/���	�#؉|载�w�3�R�V��+v/}��|ua�ݳ�Em�Oq�SB���荊B넍|��,��^>P��v����t�F��=B0��VEջ�K�8��+���\�PW�M��v�����VA���B9�UA:�SA:��D+���W�,�4��x�Ӄ����yHn�y{�����BF��ܠ}�a͙�"~���X �������^M:cp
k��fih��C3پ���������rwq?>5����S������횙�x�r����c�1;����^MH��UСOD����L��0�.���/�Uy��0-n�H�s�^��k���V8��A�z�uf*�WGBP*cF��W���N+8��@�����V�=�f��e��Ru0�9����ͫ�̽B��.��b�����r����q�Q�I�RJ�D[
*l�|I<N_�y��M3�`�j�e��6J8�E�f�FɊ�i��L
�蝘֙nʺ��S'q1��F�Ҿ�y��i�Qm���*w{�[�E��wS8�^{�+��$9fuB5�,��E/�9G�;X�^
�y������5L�l��Ӄl���z�K��%Vg�;f9�f���k�5Տ*����G[u�r��[������+�i��Y/k{1��YaYsp�_��z�P�*�k�+q�{ۿ�BI���V���_T:*hXj�2^��7���b�dS��ٔk����oK��[��9�� v����y� �e\�������b<�f����vb�殲P~:�
�N�n��]mw�W�����p�0�e�j��zQk�r��zE������n�ﾈ��6&	�������̳���yt�յ�DW�W�D�V�~
�����d��|�V����ŗ����γ�%JR�d���yY^~���rj�>63�p�w�^�5��\��7T�^��W��>_Z�S��hǴ$�B3��UΝ����<���ij^Z�o���w�^y~}�P<�.�l����{�u��PO���X�+����$��S�{=�'�J�h�mɧ���rN���Z�֑M����*q����|�K�O�+�xnŜ�r"��5qG�����nN:Sܺ�A��9ڜCzsj�FK�k�;[�Y����Ͻ�i	�=�VнC ���{lYLeM�~3�)t��X(>V�i�L��xa5L��t�>ӫ�\�,xv�AW���m�@���%�9B��o
���@Q s��hk��6�j�����x{U7�	,4������v/���cI���^w@^�N�q!�ݢᬐ�淚��j�	��I!��J�O��GC�z��i,8�6�Pi@�P)8�Z��d�'�
Ȼ3�<������ccl  l�ڄ�I$��e�Ā   l�h`��   �   N[m���   ci�f\�    m��`1��  d�  @ H   n  H  ��24�2Cm���y�U@69l -�   �$w�y��+��ڥ"�Nz����:�2=�w���=T|�)�3�YZ8���[�w�\�j�d���=��6����o)8Mȡ̹� ���%5�����n_�-92�x�ڲ79wlh$û���gx�Z˨(�*�b��K&Ǯ�%�)mԀ	ډH�Ҙ	w	IU��@��ٺn�<���Y��<�%-����e�J�G�>5���9�0�Qի+F��e�]R��}%N�k%Ia�}�{�{{��I��+��*{y�|"�s���#�]�����D��h�pd���N�l����BBN�m�m��
W�u���_j98�u"��W���n�v��i�g���qN��c�ku]s�qj�9�� ` 6� ��1�l  > �$�۩��__�0>��8�^��.�M�UV��j��{�At�-=o)p{���c�n�l�NR:$���|۟�fI��K�����ϕ߯&�S�sĝ,9�5��ͯ�%D׽���'��k>r�!җ�s�!���y�0ꏽ3	v+��J"�y	��B���P#QS�
(�3+&S�w���:ӚL3�"�mKxw������BjP��].�N�ٛ����S��x�>�^��;n@E8�`�#�阜Hc4)m���0u5:�Nʅ��x����Ez�.�����+{" �|�LxJl�󎅠�.�.kU�M�r���3x��v���mu�I4L�"� Ь��Q�1�Q43e��3q�(�c(��L3Â�BIWx؄�p�~���l`��՘�e[���%06l����!��t��	%tz]��c]�>\�$���w��E�:�wC՝>�C���[�A�#��j�i���J���d c����s���Y쨜�Ւ|j+��'d�!���L�wwC�$|3
�W${����lS���j5Z��滜��v���h�W�U����g�'���t!BC$~*L�W\+�x?���u��[���RT�a�,���4G�P�X��x+�X�J�.�f[�T^g�ce��R�,�&��̭���d$j��/����6�p�(��RT�C�A�ޛ{&�n��у���f7x�v�ĥwa:e�9�,�jx���*���楃��� B|x %����T]R>Z���~���2�`��t�(��_�G�����o�d�u�ܐ�b��������F���{�bZ{��S����?�Z��̻�^x���������>�U�q`Z\�nLP�11\�uD�i��#"���%R��9繋\��h��mEE�3���F��Q��G����DN�&%�ݳ~x��U�*�q�{]�_�0h��,"���O�{�%�+�`L�ݬ�e���^7�4��ZΫL�`���{l&X�t��&&R秉�Z�/������(G0����h=o�ӝ[��>\ݝ�vf]٠��З* #\��xw<���>��h�ͤ4vU�����h��Z$w���+�˝�v
W�5�|ik�^{�Pai�<ρF`��5'(�a���ގv��*0l����������9>|��6ST����d��ٴ�/�O-4�����(H�b�Äx,���I�	x��Qc4���"ef�c�x����À��nK���#ؼ�M��mN�ʨ���S(<��yﱞ����j��!��W��Oy�B; Oo�ܭ'rLZa-VS�+�f^�<�0��,ξ��vb;�f��`lq[�7T��Ӿ��S[݋o�]Ĉ���8�܀Ӹ����`;N+��w���t�lXs���Ȥ%df�%�;�k�r�O��|�4տ���>�Q�)&N�ve�-�����#@�n3�R����M��"w�KǗ)䥘��@ ���d��� {v��9�)Y�%��gﳷV�nh*���/5~��%���7y��i�s&��CG�����p�yt��D�7q�2iS�<��'�e<����4! �=3빃�4�U�(
c}�U��t�������=�$�6/O�<I���mn��� �(9���v�U�:�5�L��X}M�>A8ruZ��Ϫ�ۇ�c���|�`ʆ^}����~��릙����OmQ�U��,*�QWX&P(�
$�>�B�K�wE,���ɻ���s�q��ѹ�b��F�G�Z�<v�9�@(-�w�POgJ��|��v��ꐳ'ªj�V�s8D�9�a�Rj�����<��6{n���Њcĕ��T�8y���{�{��_Y�c���yy�k�e�,�`��J=&+��Xca�B�uL�U/���EB�5��6A��{�2�'�r�8��a�XL��	���c��zrr�	��jyLP�o)�s}Fb��sH�r����>Z�vQɱ��-�&>�,��y�;If�h���n[�Ѵ������[W�7z�\x+��zVJ��r�34���6�����*�Q⪱�Kˊ�v�&;�/�o����/:x�ߴ��0/n�`2��$�sc�=�<癠�/�`õ��+�D!~�^���6H@�FZ�V�x�ȮFg�$���y}�.��a�l��ԁ|�l�^�:+?���CW���G�Q;`�(�tq����V���0؟z�%��KC��WwS�� �9��P��"O��r�]�&W]�GI�E�O�8g���a�O�-��ߺ�益a�Y�Q)(�A��<��M���'�7�COisk/���aJ���.����]�VB�;��B�B4�X ��p(亍���*�v�v !�E)����C�^����q��d͓'D~�2_�g������ǹH�����}Q�k�s��_�/��"d��nf����y:�L��T2o��#J��Ѯ����%u�=FWV�͑3�5^^K�y�P�&�W`�.CB���/"��*�-u��;$���\��d��.i�yT��3o�z�꘧��6����M_{׬�7��Q�bO�q��T,�@Z�
L��O��Ť/;�F�m�<$c��tK�&��F;P��(x/_mL�N�2�>�2ި��}�_������)�G�y]A��^42�tzN,��IZNOf��6��_/�Y`�'r!wϳT�s���&ܩy���=}�'K|�	�sVnǌfImD�����V�v8������7�<����Q�f���2�/��  A(i5c$ !	�H	$en�2w.�@;.@���J+{A�K#3��_#:V�~���}T`��s깽ו���Q�m���Ū��}yꢊ�S뱙�?4�[�E�:�˺���(�ϏG����.�M�"���>�Ge��HƆ��b��d��l��B~��[�sd��PTr�'Mxo����A���7w[��1�w&��W�'ua�W���Pz�f5,�M������w�;M/RF1�����g�s`�1��"T���R�U�L�?X��N�~�������m���}w�ۛ�U��R�}�-�Z�;��2�O5J�tpq�:{���]�T{M�١� �`W7H���/Ĕ>X �9-�-i��BI. k�D8eS�1�����o��ԑ�)�	��XWzLI�&c�k�<:�ɼB{�)���&q���t��r���}D��^�B3T��o9��sS�*#�)����iR�R��_����۔&o���"0����y�*2��"[M�S��]WtG��|֙�!��s�E��J��X�>�Q�k�C��Иܸ��-] S��uۘ��$G�������4�X1��h�J�m��5v������	�v����0���_C�n�za;a�h��+�Ӄ�Yf(^�L|uY�eeՂ�L�/��?Zם�n�a����P͔�C�J}7s1�5��u�Vn�K��2�#�߬\�
��զ��1e2
�G#%�}�ة�\�X=��U��;+tU�������_nϝ��� <M�H"�L�S;N7+�D��r��<袖=������Yu��[��
>>t/����T:d١�� z{�r��6�L�?��~��̓�c��l#����R��a��1�4 �ɦNi�HU'x+��5�XWh\D��b����ϳܾ�#��Y��Y^��2��  q��EY \��<�*(��F%������)�:|���������41��٣�RT�a��y�Ɏ�Y�/K\0�y5k��^���G���'{Jr�ۻ���ݳ�f�-&�`ɟ���\Z��g�~�N�����y`���	и�g��͚��z���|�qS5�����a��1Ý��zSB+��ʬ�I!�I����zN���[���#�p��Ϳ��ܼ��ο�L< w]='�3ë�$;�@����͆�n��4&��ϻЮ٤|7���&&sgF���1��c��W�� E*`�%]�hW���}��ɚ^�'��H�Z���)��ޛ�$��:פ�ǣsv���Qm��T���AP:�*����W��{�oL��s���bײ��R����,�3/{��JwkM�ag'f�f�u*���m^[9���a�5fh�#o[�}!U�"y�+M��M"sWc�n
5��T��
~�bl*��7�Բb� ��h8l�墨�k��l'lh�hH�c��2���rt�Q��z�>��I�{!ǉy�ו�9e�͛/�Р_�G�%L$䭂Ѽ�3�	&4r뛎�&*����izs�k�y��(
0�N�]E�������ꍘ�y� >�B
,�����5�o�}{�q����B���0�\p��3{��:���?�+�/�#2c0j��U�����}
�bk;���z��J$r��~ĥ[�K���HN�MGVW��O��������"�t����b+��C�#.�li ��i��tT̏Qr`���]U~Q`+*���ZF�nгS]��X ����1t���_��/7Y.�c�E�{L����d���`�;z��c�֬���sc�x1>re˵Ӱ�il�*��&E)���BX<���r�mo�3�Z>�:���k�"-���'�;e�$��TP��5�/v�pT��\��)im�X���{=l{��)�X�^Mi:�<=C���M�V���	9nG��6Ҁi��+���wS(3b2�;�<�h����;is�]}፪�Ag�����H�{�M{m�֡a�s��i�+ɐ�ۢn:;���]V<��{���Y�ѳ ��#������7w�P�S��J-�Q��p��;����{T�Gۜ�V(�̣2���m ��7c��h"��WT��ʟO��+j�05K�CMR1���Z�RZ��#����������,^��a�N�� ��X����k�S2���H�4��i�����3I�!3癩V㖨�7'�)%DV�Iw�97GZ0o�za�k���v�I�[u�s�e���`1�Z`�+d���kT�� ��]ka�B��@����G���2ޞ�fTK�6�X�"��1޺�I��"����j�$��^ul���翼͌���w��¬�)�:a�}O<L�r��P����*ֺ�sq�-����랗�@/�:��j��kh�
|iU�J5ؿ��G�WrO�ź�[0��r}�smv9Y�RPZ�!��h
�<��?����.�g0׳~Z��{�w�[���k��%�Q�v�I�~���� ���C��8�l����'�JY�~�mҤ1����C�������g,�}xQ�������O���C�����Sc�M��GV:  X��P��(�]�f-�����L\��O��,*ɘ�$��eP�n�Pb���L]��u[2ى�����y��
�T����׸5ծ��I��K���oei���F�qF��M�]Mm�Ckc7H �3�S��ڦvksP6_k|4��n��$���Ȃ(�1�l   $�`�ƫ��ra��I)I#�qM�Ú;X+���P/����j�΍wt͒	"�6��R�UХSSQ=�����x�8b�m��3Q��퐫�3��ﯲ�Gr����z��h�GWa�-nZ9tL)�?_�}<���u�Ř���G'�.O]��B�權�x�י�S��7MT,0l�/�L�������C�X�����-��v���>�GC��+���e�]cW��ũx��������@fs�k�P�H�W�4!>0�`&/�{�����������̭n4o�Uʿi�<���~*���{p�=��]w�)���O��V�N��&�~��c�"��\���^��A	�Q���/⁮�߄l�QSѣ%=٤����k�����O��������O�Ֆ�7�$MXYG4��,.�x��ܽ2�+�q�X:��5��jk���	���*ɌJB:��QI%�a	~�C��ߖ?(|f�)ίlm�ƨ�m��� @��6+��^Ķ+=��:z��G�6���<D�އ����7G<7Y�+vM?OrC=Y�N��x'�v(���
�>/[�-�B;w�̱���m(�?Wn
U���i�T�-�L���T9P�p�͔/#yA3�s�����Qp�vQYN3�U�)�v)Afwu�y�9iFQ�q�h�@��0Q�SwR��
!i��A�l귞\�%�&G��:�o%�zצ9J����X���ؼ@_���ӳ���(�V!�d�b���=�m�zɯ	i�j�R{E�Ƹ���Gx|��T��}-��Lk�4��tu�j�]^�-$O`��n�\�!pr�  �~�������P���Us�a�zҸ����.�z��c��w�������U��T���:���� �<ς�3Ft6��I{�p��`�����Q?n��0�f�ԗ-�k���|��Y�\W����i�W[�	砙��Ȟ)v��w�$E@Ki�'z��z�Q�ti}7EW	�~�ߎ�zw��y�ECTQ����<�J;�_�z��$tx���6滜� c =�j@Pڰ�9:�3�Ay�ü�M��AX][���K�*iI���Ωq6U�I�#�w�o"}V=�5��h����p a�X���5*̆w�`�Mj����n��w���m_�l��e%x�l �� }6v����|��������,���qo6����#������$��q�A4[�ϻ��u�r0�)�9�3ϻ�6�
��YU�ԙ��̉3�֭u���Bb]�ن��n[S���w���v������V�3y�.l���j6�@�M�7�{3���miL�MV���V��b��7w�� �QP����Ki����
�]�_?���CL�&��uh7�׍�vޫ����&aS6�?`�v�^"��Ղ�m��Ӧ��K0mu\䜃q�}ۛ��Jln�J�p�)כW{W	c$hYs@K#͔���U���tջ|Sֻ�e��6>����^�U��2��9/�ρ�C~��|p�o]bū*�`ћ�p�rY�C�Ōf)ׯs���r��+%f%-�z��_~w[��׈<��|NV����ޗʢ1{J!z'���4w�I�L粧{���xܻ�t"�)�~����P�5������U�<lh�}�!�cEa���_|��\��K�DF��ٌO�5��#$��U�-��{�?+�}Kz����?xxxSK����Ζ��ߌ�a�� ��﹌�жt�w��>M�o��k'��oN��[���d�,s�v���
�oM˶;���~�oHJ|]\�>���*G�q9�y���@�Q�;ٲҹM��ϲ���u��,%���R5�
7���*��3�U�`[��E��S�4oy�����a��p-5K����{Vg�`��3E�Y[���=j�;D	�s���ğ���ϫV��
ȍ�EQ8��ŀD�ګ�t��u�y7\yi�H�ٯ��H��lb�"�;?-�,��}��s��P��XeNg����xʼ�O�bC4jk"���y-�����T�Á�u�WD^�kC*�ۀ�v^Po6p�k�t���O�Y9�MG�*S�5��E���y�ܫ�#:��	u��]ú���,��4�[�6H�Z(Pݡ��d��K;��3(��PN�ʽL뻓*�3�:\�r�Hv(�S:YZ3^v�r	���ͩ���<�%��f�37���X�CbQZj!��go]��'3/9m��*Ln�j�ɛǖ̬� ˗Eg)Mjދ.�����K�B��6�Gޔ��P�V8��#�ʞ�ds(L-��i"B1su�Kw��\��.�uI�V�+5X�\�A��Ù�Y,�ta��u˃J�wg*l�x�r\�� ���ᬊÛY�k$���X..=�b3%]���2N
�u�j�K�Y�����7T.���P�4n���$�Փ-[p��:W4���J(�ºSm$��g@Y�Ň�����8�h�;��� w�iy�}̯�n�)k6����6��W,6v��"��wzH��34�LER�obh�Nm[����K�cQ���J_�隸�ۺe��^��h/�p��/�������v/![;ZQ	ݮYꛂƉ��2�<���(PZ�ȹ�/He}Uj��f�T1}��"-��&d�O#r����]W�q>�9����MM�B�x�e�(�� D������U6��O����vK��8���!��ȞA.�yӟ[�qw��G����1qn6�A�.���+S�f�\>J�nq�r�҇8*�W".�>VY2�mV��&N��w��|�qи�h���#���ZK3��uL�.$���h�7ӥ��艞�v���ågd��W2��ƽߚ�i�x�;x�"2E��A�,��ʙ��X��2��/�9B ����8�J~�]�QZ�h�j}7�<Y�$��_-3n<:���A�@���n����VQCE}�4J8��{��csX�� �xR�j��(8`�4;ϟ��0�2N��*`�f�՜��p�%��=���V�P�zl������;�e3r(��F�v9��j޺�%l|W�2H��S��x��\3u���¹I�SҒ���q���7J���w�w8wb�W�q�I�����S{eo7���YW$�Ʊ}5�]~3J���/oyZQ����*=y	�!;�n�M`�G���u����2ڹ���&x�����a;����8Q�3>������_<���vM+
��1����d���l�p�,�hnz������`�wWR�f�N�����Ԅ�B螘iM�4ĭ3��j>�Ϭm[QWeʞ����xlbZY3��idc����0-M�l�t ��W.�L��ߵ]�6n
A���Mߎ�)�<Z�۫�-�����dq}��|(u�n,�CQ���7�;i����d����m6���l�'�)GQB����b��.�
Ԙ��-d�����^ۺP�<x4%�|��+���Z��KWea�3:!%*��d�)U���1G|/ģR�����(Q��3��z�g]D)��h�L̶6=�~ζ�$:�p�I2����C�m�œ�9�w�l�����&\�Z��aQ/�3�3{jZcic��k	�ޓ��=�~�)ص�[d�����l+>��߂��Z�k����N�z�R���L_���$��\,�W@�{��hS�ƺ���7X��n�f>���2U�r�ݹS5�������&��%�;θz�h�����vd��b9+�P���2c����r��h�"Id�6� 1�%�	�
a�M�mlx��/5�J ��k��PJrBa%ݽ���v��S�C���d;&ei�	JH�QQ�jnjV4�š*t�?ufAu��o���XZ�1�Jݨ:PNb�13y77Y+"Ƥ����6~ta��M�/�4h��M���j�]x��ʐ�=1��*�9����(����aOE��P����`��i��	o�b��iP�9�4eLޔ��b��{ާϠ�+�*/LZe���K��:l䉌r����%�E4�jxh��7|��kU�ny*M�Z^[�(��^��1)27�@�W�k����3	�"�[V����e��%��`�J ���|r�c�|ϴ��8*���ٖ^��s�*��jG��_��;�.uNt�r��XSW�9�s�g;3�r���i�7��+!��	�1�1S��}��[���y�¸R&ǚ���K��{+FS�U]�0[W�?n��Dui�����y�WӺ2�;�K�!���mP���mL��b���p`�|�,�u��)�� GWs�ViPh��cvժ�z=�ڦcP�N���u�)\�!�^����ߔ�$�=�գG8)��x<4���*�?_��5�
x�|5X�᭜�lc
��QPK��r�W,�,��ݺ���n8�t�^@�d�N�
ݏb|`�kf.O�=\�4�Jw��L�mw�k��J��=��:v��3e��I������J��]V݋\(/qj4ψ0���zy �oZ��y��}��� �{n���b-@2��U;"�-M�w�h�훰a��'�D�+�R��\η+#Y4�1�RLE���*��1LŔ5�ȿ��tz������t}�>u�L�`���~"��wz-�v��4)�(����.��s���YIJ�~�-�w�څ?U��<+{����_��}7F�$AM,��mpn��w5庝��o.3��H�e$w�K@fj���4=�$�YCA- c��W�%@�D3d��G��*�����oiCx�����RQk��P��L�o����LV��{��f_�[L,��k��c5���u�*��Q�+�کV+���ªߎ�פ+��/�6@ga5���%�{x��8*��7��x*
�`�˰?f��h�H�@[>�,HԄ��Y�Q���HL=��y0�YBp?��l��*�y��1��L��K�e�M��	��r��B��P�ߑ;���hW�E�����&���6n��e�A��z�uݵ)�U�x�\�+"��3��M�^��;E8�J��4n��v���(�Te�S��f��su�mc5��rI����L�Rr�z���R�عH}���C>[ ���`�Je6+u��Q!�[(EV�R�xI,3��z�k�궷�l�B��j�̇e��*��N�"3C|�b��qH4s:�,M�"�T�U���_���q*-f��q��@:}��(�)(��´��dY�'��s��U�� !����0�~74�=�;F�l?��3���,�v4� w�䭓���Dh�=^q0��xu��{�݅���[�m��E5  ���������(�[1ܩU_yA�=�ƃyh�'K� 7�N�uߒn��4gl�|s��8O��/��D_)�$�e<�AiUH���kD�{*xi��ws�6& ,�=�����~���������Q�����ዬ�W�U��-�Wc3K��?T�;�����'Rm)>�3��5����]*:ɲ�ܜ":Fy��������Q�?5�p�G(����P�
�pp�<���&7�	bs�8eP�OO��bLm�j�bfb� "����>S� 	��i��ı˜R�>.g��S|5}`�غ��~^���^����ÓmG眍G��������a�=;�NW�zh� As�� �*��k��l�Pڝ��m���ЌL���k��bu ��uP��rxoM�+�W2�(��4�>�s��(-�Y�c *y0�S��`{���Pϒ.`��'�,�z�L9#�	��At_';��x�˱�@3D�k�.���}�`�]<0d&���z4��B��ea��_eM����6�P� ��v�ee%�)P�A6�E�E�}P(�3����vY뭏P+LW>��R��oNA�ˍ�����ʼ�A��c�Fi;ЦM��6.T�{�60��-3��h�%��BP�&�+t�'�d��9U����,�����m���:�f�咧͓~������ܼ�{@�`�x��/��~���~��3���D/�u�Uc-?��3��ƃ��+u�o&����ϽV��(�,1�Z��f�2�|7=g�P�@��9�5U�0/�=^F$F�VX�u�o�{cձ�1么*�w�7�P��$�ya5�E��i"mP�9x(v��̠8����K���ӹ/��I93/��k"��o�V<L+> ý� ��Ɖ��pFn���uX�.iNqj�ċ����	ϲ��Ù��|&9G����L�QD���L��]*�û�"���e>%�]�c�Xv�
��X��íѼ<6�c��lsD��0����K�kv﬋��[�$�h��S���U: ͜w$�6*�7ט5�Gt��.�@�Pb�Ê��h�wd��b����2@ #�	!L"L�����n��Bl���l��2݊�vRWg	2���"]���製{2��b����б��˦㮣�sE�x�*ի���94����!��oyz�ذ���&T�mEI3��R��A��L���K�<ltp�#���^1�h�K3C�ô� ���)�4������{�Ǥ�2��Z*�Cg�^�X������s��|�~OY�����uv%�2泣ǋΩ��٠/������-]�c=V�W�Q͛���I��?�T�����6�}����y��Һ���N�G_� ����͈y�Y�ly߰���1*�V���Z7/Esza���W���oz�)TC\�J֔�6�_��� �5�����h��V�5px1�90�䷲
���<�C�r�i��+�_V3uv�'G�Y��k�#��2$@bi:�F��8����k����s������"�L�0&�f�T$���4ʒ;7
��L�k�Wj1��Z�p"�	3O%�=�ױB���@ik8��#�̵����*+/4����g�{eIrl�Q�D����$@a	����f@�=PHԆ̃Z)�(�_�b�݆�+�z�ý{�Қ��W��uK�F�Wi��;5n`)�ѝ�:ƻ�1�ͻ�bĺ|�Ǥ�{Td�w:�θnZ���lS:]�-�#P__����\.nQrj3��qnq�S�&'8� Ŋ��^�?|=�W���Ѹ�4!�l�W�7΄�xL�@K��@��w��cН?0���_k��@C���|]� 8�,y>�������~�h�r�%I�M/���:������ļ�<8u{����{�e'�����}��%�F�Mq�sNҲiٵL�wnk�:��0��)i����S�/}]�_uu�=>��עs���y����n3ʻ՗�9�O�~9��ƺ�}��>\��"�Y˿r�J�G�v��uK;�ܛS����W�k�~��hG�V~�w��P/����(BI
_��U��/�U���
g�ՃK��j�J�<+W&������X��Wl����,��d=���t&w�Y�}K�#g�5q�&<㬯��=՞��啞����7��G�l���EC*h�I�/��=̣*g��bl�gC�
�U�a=X�ɓ9�j�yT8Pd`�p��T��
��v�o����y��ƫ�q	����T\xq���D�����b�W�t�4lmV�Գ:���!�>׺��h�C÷�ep�klRrT觴ڮ;�)l�q�+��h��ie�1�lwR�Xq�����xR�.[����]^���*5LJQd�D�_	m�z�AP���~,�ﳰ�FM�Y8��qƲQ�"��@���gm�*&,M`���CU������]��m=.�_/��my0��A��>���}�8��f�S�еWU�̊wF=Sm�^o�[�����F��W`5�[�,\e�2۟J��Z� ��s�Oa1w�m~���w�>hg�ۅ]����^~U��a�,>KX�y�6D��7֔�vi���k�;h�5���Q��tF���8��9�ǧ�cj�YGD���]f9=��ϣ�}+<�⼫&��h�-�o:�Ka�	��k��8����2�\y�~52�Ly��	�Q��P���ӝ���Dg����6~��6�����O���o����d+^C<���������~�P��,���>\�i��ʹ"S��b�&�W��L�o��qwM ���}�U1)�];S�E%	.=��Y�����P��1��uʃ�I�펾���+VWeNĊ�--�1ܨ�ޒ��/9���)��۸�Oh~&J����<�f1����M���"]����t�C%ٕ}3/Z�yO�^p�֮��n��{_v���|dh
s���dV����Y�uRy2�s1�p���{�]tzw]�����YW�툕�?w���L���M�A��F��@���6�k���G�Dx���ȇK����
����/_��O�U�\x�9�y�͹<��:I޿}�s��/�h��!/��+����%g����a爪ޫ�X�J��OFf���fWj�d�+���F�������xbB,�Ӯw.%�I�$L�dy����N �q���YQ��B���)r�{�|���w�$;����_{�G.5�S�~�1�K��8s�@����vZ�O��.WʴN��hA@�ާۖ!s��M����t+�B���ۂ�Ə�����ǎ���v�or�5|9'�r�B����8�1��{3�\����0���}��F�d�i{c��.ٕ�czm�:�E߾.ks��|	�^\z`�d�:a39�K��Vtv5&i5hi��"�,���
÷3sE�䭨�eu�v���b�*��U0��ehv��}��X�^p����<ref��Y���!�ڷ���&Ә-&�c�nF��@\˜l;zOu�#�k�����0�.�����F�+٬n�[Ֆw��.S��4\�CMÃ!|�H��c-3TxL�tᱎ� %��Y՛92��[�������e�Ep��c��4��L ���x�6&6�=ޢ}�f��e2�×�J!�tY��
��x���i>l����'\c�X�~�6@,���zIv�,Q�̬-�4�_-[���W'�KtD�*�X�u����{��1�P��7i�16H^�sG5mȆսw�rJ�L�g}.�`��t6�]�W8����7?.��3k9֌�-�<��lu��ګ1�sB�\[�w�vr�ɡ��wN��:��ɝv����c��ZY��ݴ�qaJ��u.�b�1[�}��<O�6�l�'�33�ߒ�z��a��9��I�9*^��͋ă�S��m�U�7gs�XY����ȺlV�蹔���m畷g��=u�IN/0��������Q�<KVw�aB�"X�*<DX	�ݽ<Zr�o(�r8ȯ��Ќ.랧�rM�bm�v���2��
�чgI�#��:���x�L.��+y'֗W2��b��x�J�y-?���vB;H]}S�ٺ�&�:�߻:6�NhT\O0��MUe[灧f��<��K���rp��R5Wڿ_q�7)�_���m��>�������٬/���;n�#z�s�N��G�I�Àܭ��%�34Y�;�ٗxΕ��q�KCo��;�Ʃ���=2ۺ�\y����8CB����ݥ�ɾӰs�et��c�� \�ݶ гj���#]s|���wj��K�����h���NTM� 9�    H6Є!�la2   m�X@  ��6�[L m� � �0���
 D4�� �HjH`   6�m�r�7-�              H�� ��!IF�  	  d�r^��5+L��h �*$�og]�@��ooM�3�le��t9V��wpew���C+�O�5qr���nNdS�,ȗ� m�KI� �)$�$�D�BeB���8n5a{���9��D�L�Qd�Yrk�l��ϩ�S��a�Qz�.gV�*� i h�	��	kt�K�k��Nֆ�����9�91
Y��Y���7D��6�u#�W7d���qB��[,
]�;Xf���z����bЛ��P�G�7�L���suɻ/
�pJu�.��sw��0�ɂM,vO��"�{7{��N9]�^�c��om^VS�\�?�� x��r��_Z����Ϯ������W<W�er�Κ)�mF���LR0I m�HCm�   "�RIz�l�{�ݕU�Th�T���粐�vH햲�R����Ѳ1�2�x��	$-@ �H����n��_���z���F4J�յ���s6�\;��#B���j�.o8�N�WGs��?���v��=���o;hCݏz��>�����co�̎��h���٩;��G��5����8ϻxӫ���~G��{=�c����Z�/�p�VSH�h���j���I������7�:�%��yC����{6��)m.�o��7��ť�d�kߊ��R����?�4O�̿SV�3�i/��b���=�ַ�ڭ��u��5������w��u���4�yP䤆J�~Wv��bk׻�n �e�157�ؗ5���Q U'&��8��^������.��n[��~��{�n�=��f�����!�lzI�K���D�꿦�V���!E���K�ѭ~282.@����۱���W�-�8�n6�2d�� p�{2�q�mΎ��������g��)d��غ���Z��s���%u�)j�gnKy�=��ZH��%���-�LY�`�]L+��U��S�ޝ7C�E6���lz�^�t�ݽ�ghq7]�N�|��fB�#Ѽ,��gL����YӸ������˩_QU����`s���huE��8.�@�^�^�ݽ�zFT�zj|sqM7<M�U��>fw��޼D�����`�z~��#�bW
�c�M����ŇS���|�ކ��^ϰ���o�FS����AwSs9����Y0���zj����A�쪹v�b=ћ�N���{���{1n'2��3���[Y�j���*��v�LoJ��ު���q�nU׾nb��6�t�;�i$�DUS�t�@��5����+�k���h0ly�ѻ�%���7)}��\�G\Ӂ����=��;��V��`�"��pr�������pgt�̨�֯&f��Յ,ˁ���rS:�}5�o ME��Q����f{ufuVq�S���rb��fq�=�~��O����(K�J�e�O�߫kWtx"s�~�9�fi�WZ+̂��s�h�������ul+�ٌ;x�3)H*�_@��&�����b�Ti�ݝ����G.Vį�l����tE�Ql,����3�97���Vy9V���N��g�K�P���}�{��S�.�]|�~��f����ֲϳ=h�m]+}����k.���׫7��.��:,�� G�ܫo�Ԫ�{����n����{G$���0�zoe|�����\�/�A.��૦z*^VJ����+���[��I���bs}�Lα<����р\Li��,�^���2��^��2����\��;7�%9,C̒1�7�.N��>;J���v����U�n�����"���n����5�4�D���̙;.x���
�׆D����K�5Q�5qg�69[���%}Ow�)N���F��`W�ψN=sN��(r�.Jg�I�6�p�}����˼(g�������t�odc�2d��3�iR��4$��<=�tea������.c����=x�#��6]	st?�)54_`���]�)��8���k3��]VaM�T�ȷrx�h�ٳ��R�+�U�^�*�{]=�����[�B�5uj�`;�#y��������i��2�r�u$'e!�� �f���,��cr�o�ٹCU�	�[9Kk��\����=&�@�^8�	�Y�(��衦�����8n�oϣ�q\ipϺ��LrM��W�ՌT����K�~�6�վ|���<�Uz[��oٺ����-��쫓����}�4Y��uL�}}y7:�͒�r��7c�)J�O������Y�C�Jf;�,=~���k��3�i��*�ʧ6;��j�\�H��	�w+Y�硐X�c��q�u���Īn��K�'�fxz��G���Zq{�W�w=�Q���Ϫ+�u���+����҃ݔ����st<�>�P��D�.���ė�tW]�K��$�uL�=y�G6Y����:�ك���.�|����p������}s�,���݋�h󼻉ڬ���=��Εl��2�n�w�dE\�5PHZ�N�z-�B��6`�9����h]����LE�ll+���(����$ йv��Հ4{c�x��j�I�k/Y��������1�iUޝ�V�\;oV��716�y'W�O
½���P�qӛw/�����t}�4wV�#�j<;�Ҏ�t�+ji��gfC�r�<)=���l�,�i	���Rю�2�qΝ��6�B`� �*"P�p� � @�$R�g\�eu�Ζ�� M��M�3��;�����ڱ殲�������$ݮדq�ԮU_iV�;��دnq��v,��1���v켟vd.�k�Vz}�_�!��| m9�$o���e�����9C�5�q%�����MF39��,<��>�Q��݈���{�����+u�E=�V��9�g&+���)|��1�������Z捴3�����W�I�k�U�_J��/c�u���s����w�y�矪է� ����p���o-�^��ň���硋ٖ���Z��Q6����������W�*�F����EQe�Q��(�z3)�s���SF������Ǻ��>i�P{1��&�Ss�W�^e��8\�, �:��y>/}�n�S�=g�:���??���I�5�ƆiB�
���1���oA��I�i��n�����O����_{�%5.�_|�2:��Q�bbkk�:斪gb�t�ih�ň��\���XU�} 6�r�r������{���dG�̂->��non���Պ��l�/o0��Ζ��sl�r��8n�����2�2��zM�<���XD�Zԧ�Y�o]�X誔��/E�ҏA����V⧥H>�ݻޏP�x��'��O����/�0���>>��v�.&X���v��?m 8����)�
v��f� �Uݸ���w9M��{f�^�|2&;���W�%��.����/v��{6�����|�̀�Ո��-��$���:w�]��=��g�xy��{����>�-���υ�օ�/���<�x�^
ؿL��>�zNh�ٲ��דv�B�I3��S~� e2!t?y�Y�&����.T�����ܲ˺ֈƣg�Ҕd"B��It�ML��\��x_���D}藓�v�@���QA�鹪���;��$�QMY|���{D�#Tkո�y�.t㬓��r��d��y>�41�a�������q�w�8!�4�������u�7F����t�=2�9���"c��9���fn�쪦b\�����S=�^����5�^,�F����O<���:�h9�n���fYȉr�K��ܻ�{t��`�O�����b���LX��u�IɗYYe�pn���h�A�r�<)A�m&T��7�]�GOA�Z7J�[���qo���X��K�j�F]O���qV�V�Q�wY�ֱV�;���������]�g�=y�+�@ӑ3*߻�L_Oԕ�{��K�S�מ*�����3�ϝ6��̨�-.����,��*�VL����9�xd��'�K���P���qꎺ>�w����ꏧ�Z++;+���i�Q3U:�W�H�7����r==�r��i*~<�	�u��D����G<>�����H[�5�j����}>���o���>���B���J���:߳�c�Ǳ���_o�[�p�*͏&�
��,�/�K��~B3�V⫰�,ݸ^X�9fj1�%�=�=�`wz]/��zn���Om�sV�O�j������Ѫ-�X앰"}�<#��U��+�<nM]��G��r,?C��fkr���q=��iwy�G��B���b���X�'L5i;�}��+4����V�#�}Y���zo)[��K�Jw۝Y�Y��g6�:jKw$Ԫ�r���!8����':2�.S�������ogB3M�c�G�>�P���ڼ��
t��0ww+n��	����+�zU��ᗬ��tL���jb�E��Q�GǪ&���=����v'v�v��6�����ݏ�~ϋ����~�v���DV�� ɻ��RBr�6���S�%'.a�ٙ�g*��մ�գ�K}8�FP�g5tg�5��էx���X��s�v�N�qX˗�u�K�r�W�&�}]ޙ+�O����߷ϝ�x�Y�]��������>�03�V�4$�/R����Y�ڶ�~�n������s3r�]ߕ��q��<�OU�϶��{:�ue�����S��ܿ��_I癋<�R����S�+~ΧW��ꊲ|�/K��2���=�S���n-Z�]W��Gtv�yo��W�w�Vf�{w��3����N�y�P_1��/|�hr^&{:�{y'����׉�<���s�vÊ���U
%��VT)G�g�0�q���6g�>}]y��q�^ͧ��C�OkS�ܴ��'u�O��Y&�y���] ��;��浇�f��|�^�Kڱ���ux;�kyLʼ]F'��9��uh�2�Q��%�vV�h��a��Uc+� ���ctR�1�oZS)�)�m�IM��c$  RL�ųrgS�T&��]�Bʪj���-�YouҸ8�'~W��t�b�*K�@���l�)8�ݪ����U�D�{�}\z�ǇTá�Z:��>�Z#u�Gv�)dR-��6�
���>wp>����^�w�Y.U���m�<��.*F�{](^�$]�L-H�f�V�h\j�YM������0m�?|����.o[�������Q��m��G9�kx+3ю�k�y��/)�J��f�E6xw$�M����fx%��஽�al;܊�P�#�Ã��G��5{k��O�M'�8�~Xn����S��xP�c������"t>q�y��pv*��)ѯ�o&/
]_n�勣so�;���xnMzn*��Q�vϑmCI'>��v���ͬ����s�Oi�΅�M1ճ�7��h����{v��ΜϹ�қeSQ�gOP�������i[��{Ǖc���P��ֽX�|_���>���fp9�F�������;�ݑ�3�>��,z;�P3/n���K߾#�$���|��[2��*�F�fn�&��ӵ�dS�=��l3w{$����A��b�v��e���"Ъ�3�x��IVX�`=3{mL8ڽ�8��:u�3��[a�1�ev讀�@�K^a�yϠ�	g)�;������{�o��zߵ�^��_���s�J�Ù����Y�Wwl�L���ɱ��!�}N�q�b>���n{7�S>�<�b�=���..p�3�c��r���n�@���6�/1���B�׾��齜�L���n.����R����y����wȤG�����<���A�{jEY.���إp]�=]���f�}P&1X^sfD�����F�l���K�o���}{�`!�޴�_W�S�\f6D�Ծ٤��M�)TI��>���D+�f�f2_X�����&|�����l{m��&ۯw���|����癟w���~|̍��j�� #�����46�.Os�Z7���\`C�0s���^�d�s�w_dڱ{ t�Ww��!^{<���㳆���� ���0�<��8�\���=R�|��:�yw�0O�Ϗ��+#��p�X�\����fM|�7$T�;vv�����,`�N�M��^�Gq�{��Va���Qx�����.��TOZ���va2���m�ǵܬߎ��@�ܱ��ml �H*��r��s�5�*��� �Kr������'����L�s{�W�.b��YuAs��n��
e��N�䂚BH�lo\9�R�l*ĩ�r��wD�_�⫕1��d��Y=o��*�'�%y�F�����G��{<�������
�y]ׁ
'��x��\XG���겠�nv^ni��T�g;�7��Mt�i����)��˰,c����H7b�V�Ëޞ��*���M�s�'=5�y�)��=�ˮ�<��r�.		��`$�q�W3{!	y�v{5d�g��;�';�{�z�P��]և�2��s� ���� {����i��q��a�m���z>�{´�F��?�����Np�I��|�BO{�λ�`�w��{���=���z���@�$���Z�3�!�'��}�9�y[zwz���3Y���s{��I=g��.0&���<�;�{� ��ao�	=���+'P$�:�{I �w������ļ<�$�|a��&��v�&s����K��4�{����1	XBI�q�x/�0�ܹ"A[��+��ӑ�f�ŝ
�; *k*��Z�x�=/�>��0`��i���G��%���dGSw�g{38ʹz�wԵ���U����>�W��_*9}�ד�MPU˦ws��L틂�G�<:��������L�$�x�6���� �Ҥ���vy�S���vo�o�I�I&h���{��*����Y�Z�]� ��߀���e�OӤl�S,v~ �xڄ�d q��'� H�!�,������Y����r<7�@���D�/D��[wYK/X��u��f�rf��,�ذ9\K�EBk�0��-�X��񩕵��)��/x�S�8�����x��w_�Ǖ/ �U��>�]^Ν.����zuIX�Jfqc�M�j��z�}�l��>��ھ핓�I�|�e��!�#�;���J�Ւ��_: ��0����	4ufԈF/+3,� ���U}�.Y1�y���M��׻�Z\Y[��,�v�~&�)���#��$�0�;C"�]q�u��v��:D���� -�`.�tK���-MbWid1�WX�=Q���-�����OF��*�ժ��l��\��N>K�yK��Ap�ʆ�����R�`5k��b��_Qf������P.�qYe��f3���U�L'���ɭ̦��j�l�|h�p���ɗ���Dvѫ�oV���t���r���q�>��kD��P�n�ZuЇ�)���nI'���qV��,e*�^�@�!Q]T�.AFNbM}k�� ���GP'���]c:��w&rƱ�k
!d�H��Y��2j2ɨ^�йک5BZ�G5۱��-ò�n���H嵽���N=�9�dJ�U��s�9�ӛ��(يܻR�9��NN�]}ݡ�3�2�;�u&���\�R�M���{_�6%ռ�WGak��p���}��TǓ��.�̆��ޟN�Aks�c���3vĽ��rW~�����l�s�;��sW{�ɩR�(����Q��cӺ	����k.��)nw�-���v���e�Z�U�o�ڍw��ýC�5/�ɱ����ݵC�Sbw|r���۝�hN)II2�ɪ�MZ6����V	�Ѯ�������nv�:�g��M�����򑺫�ۣ����\U��k���|a�]tbd1V�i.�s����~��z����|��ݫbfpW�םƝ:���x��~Q��Q�Q�8�}�������(�f��n���͑ㆩ?{��N}�>�Z?rGy/���|�?.�}29q��X�Rp��
�V�����d]L9��Dװ"r�{*x�ft�տ5k�B��޹T:U�k2-��_mrE���e|8�T�c�����el��]_�H�T��P�9aK��TD���/�������),�����.���Km.�=9��Ãb`�nq�WkK����ܤ���0���ґOq�]��;�x�r�7����h��7��=��+�������rw�)�}��UG|��|�a��Gc�i�K^m�Lx��)v�dW��%�z�k��Ļ����E��-��eQA1훘��_Q��`Vy��+yx{�T{d�Ha�̉��C}&�~�Y��������b�'�mס�2���i�Q9�X��}n��@���I���8z���{����o�G�t�{\�oԶl�̬���������~�\��<h��g�Ԏ�֣��1�e�y7�p�l�����9p�l*��^5���������S���^۫7�J.�xn�_���J�=���^��t;ܽ׊���꟫3���Q�6#P��.��^�wQ��@>�p[�U�=}��u��7rr3�/B=������t��S�^���R}�ב�U�uyP������u���627'������Ê��^@����]˒�-O�)$ff�Z�#ް�b�b��T��t*��zl�w/l�ᬚ�s̜��4N|�����qf��+����0���pp���V'n��µm��ȂM� �nH@`  �I� ��f��], �2��hCͭK(�럧4f���nG{���m�d[F�I"h�D\)Z����l!^�~w��/Ҳa[�����f�_�/$i����mgr�d=�G;�}��/wˀͻ�{��-�W׌��;���L�$ eL�q��BO��⥟MG��z�A��\T�{�Iˊ���fJG��wjK$�{�ѶkQ�����O��w��Ѹk��`��컩\��`�"���u��3�d	t�nyz���ޢ��q[��G�T�G
��}�Ej=Wa�9���S��� �u��u?L1c�-�1'����?U�.0�z�EA熞AB��%�U�O+5��U�ƽ��%v�9�x��q���(�KQ�V�{��5fvc��}��>���w"Ɖ�d�GN���	�A<z�yy�~�D�2�ɝ��1++h���l]�tU&q'��pz2w�r܎J���]�wfG��1��rӕx��.�ǝ ��o����<�_FF�q����/g��E�z�m�}�����ǆ�}]�I��>�@���*�eӇy��h�Ȏ#3��94TRy+�S�_u�v�u��ZX� �Wt�Z������D|a{pq�v�&V���-e�׌�N�+;%hc�J�V�����R;Ъ[�y���:���&��}�>���/v+���8��oWI0���'>S<�ͼɶ"K팪ɌX'�����楥{�W
�������W>����
���R���R��?4�+��n��5_W�#�;��*��z/9u�1|��}�h�wws�}��t��c�q5����l�wmk'蝑+\�^���\�������3�}g�pD{�]I�w��w��7����+�0�x��E�K�v*ݺ3}	u)�ުT��{w�UN���IV�??*���'4]�]�8��޼^�S��K�F7$��+��׮���[�[�],��It�ݭ�7�-�p��31�����_��^vJ���.L��ӫǮ3�Q�]֬��0أ=��<���C7�!���ٵ�>�>4�ޫ�d�%J�`�]X�f���w��J���\Cy�uj�����;}���V&�mK�����:=[]�t��A'ȩi��\��}�葱�����wF���2��ٷ�q��'jӺ V�Mל��y�;s&��)s�k�KC�%�gP�j�g}���p������*��]Hy�Mf<v�aS�؛Y:%~���G;�?�.�b���Lԯf8��Tdm;�y[3?�V�7�NF�{�鬺׳m��_��OF�-�L��@�Z�L����}Y�|x�ڹm�i-�`��Fsf�͙�u�&�Ě��|���'X��9��������/I���Dʐd��st\	�[�佣p�ӕ}���t��C�ؒ����kۙ�����OT��ϻ�ٷ�#�e�X�c�d)�U\�l�o���)���MJ�;-��&N��.^͟D�Q��?u������=�=��ܬ��E�wb�w�-H�q�����S�?R�އן)��8����ΩO�(M���9�W�͔0z=�i��5��WH����y�}�	�����s���2�/c��+�÷5��r�ƭ^�%�P��雗��;M��#�V�aݽ9���άZ��N�ܽB���o�Ui�A�{��&�uv�������l�9���s�-��f�}��Q����W���G$B�Q�ھ�\�iH�r̦,s�E�>D�T��8݃W�+�[@i�:����^wrw2r3��H���T�e5rs�=�B�UqA�P$M�S��yo���Qn�?[�9���]��~�����^9Q��O�][�=w�[
&�����3�H�3��KRSؼc��'�y��^e�����P�AS��򁏸y
�N�Dn\yK�X�ջ�Mb��fL�~^V��㞟l��X�#���=g�34��`�66���C�"Qy��qUVzo����V���������|�� }ts�8����[3��߁�4<��4���G'�k&�WW��L�Iq�iHG�x��}f7�p��=Ct.˙����p�
�b�S��|V�w�ҕ�۾����M���o�f�ޝ�.���t���z�<#���OG��ӌ��k�c �߅�\�������fyQ���շp�ˣJ��^G��h�a�s�ւg��+>B�޹w&m�*��K���(f���q^�G�P:n���d�8�^ծP'ݻ���wݴ����t���ާ�����j�w��VPY9��v%�Ze�❈�lj�W��T�<�4�SH���y{�$ؘЄ0 !�B�� RR@�`2c�ڣV_�FjB�Ll秖K(X���I���5�<�h��[Ik�޶��O��@��1~z=�/b���^�G���W�	���;���§����`Q�����ele��&��v�Lf��W^tQ�y��*/}�?H�v8=�1��w��U�?�L��J͜�7��������^�T�f�^GX���t��U�{)֋�{���}��⟣�G�u��k=�˘E=�`��p[���c��pb�R�8)�w~���nf_���C�q��닁�N�~^�ng����܂�U�M���Z�Ȫ��]h�=�Wo[=��e��]1�ަ�������
�ǩT��wuO1dl��q?GƆGi��p�w��U����/c��3�4�jb�<�ٯ�����5��*ng��j�g�.=�[ݤY>�V7s-y�B�jL�&P�Tssw�}���{'Oб�
XZ��F���^?yUIY�dk{ﮭ�vk�7PrVj�Â��+�=����hҋ~'LwW;�s6�P����5$�,���Z*��آ�,���t��kM�4.l�Ya]q��0���kf�f�s�O����9G�8�֓��){VS�.�I7���wo��>��j�����%�*��OB������Q��Z����ܓ���+�컔r��+z.�������ؗ�ٍ���h-_�>M�a��W���to��v�blO��7���š�c`v�RU^�2G�ڱ�-ym�:V�ڼ��N��8tT��&3o�:{�g���P�!D���~�K�8��3����G�W�0����Vn��ϾuU���~ź�Ϸ�n���f��Y��*է���h�����ܻ=3Ŷ� �RV��=�,�'b�/�s_y��ҞK��%���&�sv�������[wc�)��	�(���+׬��,w���gЅ睛�W|(�������}��>�em�/ۓZ0���ҕ�>���Wvĥ�<+]w�1�����ٟ����iz^��7g���%��Zmҷ��w��϶yF�η5��}�:04��_z<ں�᣶wW>[��]u�(%q����J=���a�Bx͞�ܛ�[V��Tt��6��vUv���$�T�o�&Soo�%%���硼��5�&9���X�8$�V`�Q3�
��k��
�\'�t�ը)�bټ��y���+��k=�$���@,�w>𫚟E�?����j������YQO(yE\3�{��"~���-G[�b���/A��Tg�!����q�w�_��Nǆj=��WѰ���Z�G�>r����aM����W��ېz���BQ�/�pM�g�σW���9m�.;���<ݎf��صЪ���f�^�Z�g���zOM�_of�B��7Nw@"���뻛Q̔���l-��x�t3v��M�m'
��z.��V�f���g-��
�rP^��y����5.��e�׍��Ra@ן�"km�d118�r�c !�+�����X۷�Z��j7[�Q�7ٺ��3�}+'����sS^�b:#]N�]�ƭ�����^��+����"�n7<�����m�i��9�_�~]X���Nm�7�m�`����+���t������6��`͹����2#��wu���S�6`��Y�*Cj(�v��L&� \�۷?�UN��s{�k���-R�ښ%��>�nn�7�JUDs�s1:��1��|���YDµ���^8�s���ťd�>�>V}����.�!�>}~x}�݌�K��{�Q�9`W+��)��8& �)L����xHv_1l��4��^<��7��sbU�����XR�o��x!�́��	���gcb.೤6R��+�˧�7n�^T�~d��W-ȃ�c0;�V�\���ۺ�����&�v�4)�������m��!�<6�ghP�v3vy���:{����K>�o�CS��{�nF]o���'Q����<R��U�\FᎬV�c���x<�ߪNKzu�M�J�'[j��:E�]�ŭ���:6D���lp��y@zM7�t_xס=��צM�U{Csݚ�:W��z�J�m�׆���͇s o��Nb��x*w�,��n�}���2Tv�S�ENF�Q��Kq5d�y�GH;����ä_B5y�{�ES��A���˭����WNZ6�x��X�Ѓ�h�T]��F��]�b�n�m����cW���f]9ED������X��5l�$�-]�+yU[�Eq�M޸������*��٢�ge
!�	\$��Y[��Ժ�YVx�i�����Sv��5_P�*��h0ii�po6���ui#nRSUq����8j��34�P�bɷ4L��%A�8"]X����ߙ��V���l�sN�,u
=}9E���_����FE|4���b��U����#U!V3s���l��2�ދqD��!b�T��Ջ{6#�|:��ŭY.ib�v���Md�ٞ��sdX�Q�ˮT��j��y��N�ux7]�&�^��p�v�l���<p�X�f�U)]ݚ���.=�#D�5s��f��G@�yB�-�P�y,&� ��V�����g��HUr� ݹ�ST�>��L�F���{�xRŋ�[Tn����&�3I��|�\��WT�:J��?�t2�ܫ]�#�@&!����3��Dƭ4�%�v��__J���n�}�׸��w�@s{8��^�F�L}�"�2��ZR����y�$	y��g=j��H�����U<��Z/�lbY��7ҫ��p��j�{��ٻ�D� �FW�B��9p0jc:s(��}�\m�n���;�!�Z��6��W*���}�Ҷ�C�'/���qC��f콌g'�^ɳF��]�t�Ws�1���v����D(�"սsEO�M���������4�m�1��u��bYRU��4���%�o�h�}l���*����.7�0��k$��Zk4�<�!�1�ǗU��O�Z��av��n�vG��z4>�w�'��ۋuZ�M��r�«}eQ����U���j�fD% +�>�3�Z�:�Z��3�kz��d��!]��u<�$�}Kqn��N�(�7&t����ƧSr������ɔ��ASb�c.Q��}YrU�+/9�Ұ�%�-G6vTv�)�޶6� l m�%$�� m�e�2�  C 1�     6�M�� ��  &[n '�S2@    6Ɔ��� �b ��   � �  �  0 �%�P
D� p����Ӑ�    ��'8m��+��k?b���1o�9�L�M�q��{f�8us�3+^;>{�S�Z��I\TM_�ݣ�I�ZW,ڃu�&Uh�D������e�N)�!!� 	!K�&T�D�"T��?���r�HLr$a���xV�i�ۗ�#���5�;:W\N^��)�:!y��wm���f`Po7=[g����q�٫�7U��i���Nɜv��:�7��uK�1�S�҈=a�fTTR��R4�:{�h�P��c�]g���&��ii���j�G{�j����n����4�^�E�vL�v�Y�"]Ϣ��ٗ������V0��{�z2�3K��Ag��:�èVV�ѓ�������Z�T�mB]�!��c��n  $�����jsΒ��ɖ�0��ު�J�
���f�	�cp�\��a�WN*��<{.���g����k|��
 ,�B4�0/�힞ƈ�ۓ�nX�۶5��_U���)0�c[X���4����P4D�v%��zP.p��R+ْ�]ot�o��N0���5�)z�:�-�Uo��Z����jz�T�b�x*W��vK"�����Kb�]
��`�k�~�Kt����އQ�wa���-�\W��owȗ�g��8؜�AÏ�<�:=/���&ow*�����Q�I����������B�<]N5�H��%����V�|�Տ*��~w��S�yz�L�{w�Ξ�7IEW��+�%y��\�����vw�L�"��'_���H<i/_~g�Ce
�̉�݄5�n}kD�$95�w�d+�J�:�#�[�=��[T2U�.{�?gG]�C�̪���]V
�������{��9<�B�ɏ\$����I�!#�3�c˽�l���ͣ�鹵�4��u8"����y�Nɪ���KR��FyYSIԨά'k&C�v��.y�8pg���VlTi�i�@�;�G�9���c�Aٙ�0�Y@7���SO�m�L�z���'�Ě�W��QR��SI���M{�m9�楺۠����m����{����r���J�^�=�ظ��1}�Q��f�Үa'�!�� �z�Q�3)8Zz�+.�������+���e�7�W@�3Oe�y^��9;�q��{46�Xl�Kz�0�W�l�CR��Z�}�.�~�"vs}S���������1{|����c�U��f�s���-w1��G�
l*P���n 3׏ב��ۢ���(>�~��sF���v�j5�9��T��bl����qz)��W҇�29��1�~�Z;��|1�@�Қ�l6m�铙�Eh�����3�;��z�|{k� _�'�����i�D���]��	��=�<�� ��l
�jpEA�:���2�M��o�h}���&���_T1n�RtRɘ�ƟV�WS�Po �dybN��
M��hP��:��<l�A�{u���p�[]SS�X�+B�n.p1��IjJ��%�|p���J�"ҮpV^�u��%]}��ڛ�a��@�;��d������驧���ԍ�=������E�M�î�Ս��~}��Yɓ�%6�/NN]�����L���W��K�i�xH�v�ܧ+���+}�Jo�˶��
�dO���m�~||ea����*{GN��/��8�11��[�Q0:�ۻT�uF�&o�}9=�(圯�q4���;Mj��)/KD+]R����C9��9�y�W���κ1�z�:�,�׾;��F{�.3:��qd��RQ���0坞���yǚ�G[=7ky{�A��&.u�_�v��Nɾ-'���@Y~��yֺ�dˊ�Օ��δ��2(6-,�e���oԪ/,��;v���i��҃�����!��plp�Xn�J�N����?���ɛw����^Q&&�guS��4�{�G�4ˍUr���2xB/�'2~��n�^�	]�[���X����A��]���[�ν��&��X�e!���R�ś����wϲՙ�8)nD6�X��S�ƣB����+W:ǳ���t*F�`��y���4M��{��xQ��xh�XW�8qATO�3I )�80އ���v��X��O���}S��L��j����	��{�:�wy�9Uu�eS�6�H�.�G�Ȣo���A�(fuM��M:<�-��������6��Ëɾ����=i��8T�F>�I�צU�7�t7��|4y��qe�J���;NԌ�6��x�Q��)'2�_t5Q��_(�3�-��*J������{0߱��ɤ7WB�}��]n��-�PFvz�Sv�@��l�*�P� �d]Mo}�]Y~nʯ�x�k�ёQr��kݐ�D�!^Lu�j��㦺�ْ�"a��S`����{i��=w뜕pK�zt�rCxL`���;��U�Ɨn�oI����u�f�4)���v�X�"�О��'ې�ኇm�u�����-�ǐ�C=夿'Z�.��PFe�ڳ�QS�F�MM��f�wf��0S��udx褗MJ˹�υ��.������e�0չ�s�Vr��d�ڦn�������P�]�km�����@`���`� I1��}��]��uF���J�S=�X+Y{Ww�j�;�՝�:�4��n;�.���,�M��R^�����s��'u�e_΅ïu?vj���-��;5j���L�^��2<���4�՛u;7z������/;�y��p�㕢��խ�t�a�b\=���r��]BW���E��u���_׻y93�U\��o'����h��]���G�5�X"�p����g:��9�S��{�Q�YA��@��F�h�,χ��Nnף0���~�^r��淖��9[�����=N���R<f5',�O�v�l���-���t�}�]���%�����R���{�O{I>�l���<�?V�JM=X�sgSy��&��.��ߗ[&v�Ì�O6���:t��uL���S){O]��-,ma0���"����W�ڣ�0<�{�=��Iy����{R�YZo���ѷӏkC����<�7�x�P��=�U��{�,k�/k|if��YƦ/�AS�d�bt�SgV��,��)���_��)*������V�ła+����P��5\X�����ڨ���qS�ƪV�twemY�Y����҈tZ���PV��Xz	pq��U8�Y;����o{���x��	P�[z0G�k���9u�����w�o��(W��	;p&�6��ى��XR�2Xt�Thl��G�;�r��حj�od����zw�2�-�Ivؠ��d�@bҺ}\�{`阺��{�hc�sӗ���+ϋ��G�f�z��5^�s��6��ؾ�u7�Ee�+_��ܥ�یY7Ԙ�����'�x��D���לS��9SԽ��ﯻ��R���J��2zg6��m�+7����M "[�J����ҵ�T�@^`كL�^���ƫW��;f�nE��*��^�W8u��9AOk�S̺47�~�����8m+����w
v���a���~*5)O���0y���hS�~���,]�����S�W�۬w��ڨy��x�� ��:��kK`�]^��?m�r�&}�u$��*�丙��WWe-�7�e��[�5��q��97y��1N�і^L��Ղ���qE<��JJ�P+{��Z�:�r�Fh��YX���b���,�N�ի;U�o��E�9w�g���]*+.���\ž�-�i����~��QE�EC����LQ�j��j�]!�1�w3ی�2���w��k����̥A���u�}]ʾ��ݮ���\2YLӊL������

=U�{Ճ	�>�U�;�dk�m���G����c&��Q�㦷a��ޗ���m4b��hV�`W^�e��ˮ��\V7���>߯,l{�2�z��ZGce������:��n>��B����;G���M���|�1Ƣ1��bҙ���]^-�4ǲbR�͓�R���\ځvc!���Q��r���������8������\�	��=+y츼|�zh����݉��wwFK[yRX{��w��,�Օ�TY�*��in,�׾Vk<��/�N�����v.f�K��ޏ�pb�ѺZ�ˢ8s�]Ba���vT�gO<��x햾�p��t�EwB��#U(��˲q	O��-H:��)��k1����qA4?ׇi#N�1��E���ǅ�/��6�ݾ�ն^?��[P��2���|��J��ӫ��oi���1g��myF�XI4Y����3o��~�oǪ4�~�Wϙ	�.t�r��Ak���*�"}���qW�����ᤴɀc����*�͉Or��<�e��Khmc9��juwf��`�S{��K�O�#�l8b���5�+�{n`���D�[���[~�"j[��֧ ���f�];��� ���_���\��ͷ�h�ʄV��ۼ�~�ڮ�s���ۑKLnO��[�B�o�z�g����>%
��1����.�v�`��qܫ�4�gW���-i��*���5�j�G�y���jw�m��~D?4r͟PB�ܱGI/�[�8`Et����uOo&$H!ۙ�MeV�����I�W���n)�=Ia�Ŵr�O}*�|@�`����3;��~P��Ê�a�pq���@�kj��g1}AH@�Y�H��7M�W����TL�\8J/��v�*vP]3����u��(���.v=��.��d^����V����m�Z�jǪ���d��cH	��D��m�C   %)H��u %�����e@ᣖ3.���&�����d
:����ې��M��ٺ��CH�0�*h�}��;���L�w]�G����WS�R��ځE�h���#��y*��J�m�Q�:cwbd���tL�C)����(y�/�F���	+zX �S=���U�Ӟ�=�~lS&*���?g��9w���K����	�='ލz��v����}��G3�l����[:'_�v&��4h�ױkr�ƶ=��9�|�U+"zS���*�R��}ұ�c�9�{�y]
&7����+�׵[g��r�no�vCfp�� Fk�4�[�^2��F���T���g$�y��^���))P��b���[ڗ����4M��7�ܩ���O�.�M���+�~ O�����.���c�$��&*�r�NACQ=�׏�z׺g�����;�Vtu�`�ßK���ͦ�c��轓7��߶��H,��fj0��*=݁o�l(�ӻ����ks9����������/˙�f�İRV��9�n
�7�e�v�/��a���jsM�]{J�[�Z)awB`���\�oK�sq=ݧ�~�έ�!����셨�[|©�8��!n����(����Ű�$���u[4�ޗ�T�3|{��U뭱}>��l,E�y�/r�j�Вn9��E�X�N}����؄�����x=�9�뛽�m3�Vӝ��T�]g��Υ=�7*9_��t��=��\t������v��ş�m�^��6�/��C��l�޷7��1!O
��>yt���_j������<������G��~TUv���E�^-��R�V�v����f���
��V5�5��ݣ������-�g��;����f{�w*�.t,㒥#N���V��7l���O��ڼ{¿�)�z9+��5�#x�Y�<�g���{�n���ݩ[7R�M7�|��j~�\�'6��K��v)~
sV��n��/�>�_tu��<��9�z�����:W�vԩ���.�����g���ߜ�����p
������c�6���n��U��%�H=տz��:��e\�N�j�����=H�%�%&���\��ve�]���ٯPdnJdDzW#|/r�T�O[��\@f�8>̎�{��Հr�52�W6�E�f��5�%s�;�1�.8e�uz *[���v��`OivP����T�Ttb13���Ժ�@��	Ǵ��/y^��Ʀ.��;�v�AD���&Ay��Ӌ5��W�#<�\���W�\�\-憍r�tZ�zu;G���e�8�E��<�L��֥qWL�w/������X6�dW7H�)���Y�S�Sܖ��Q�L�.B�U��lf�u�|"V�U��Qи�[���.���Œ1��KP&����p*�e_�ʎVlv���˩]����!�y��l�XyU�뀄�
Jk'v�X�K:J��(�2ٔ�+�Ee�Yc�/��Pk��䜈�.N��hV ���m��G���{e�OD�=ͩ�Q)y�QڙUW�����6�GGF�����{c�Gx<[��#��2�l�k�Y֜��#}���PbA޼�V=rHP�V��2��mL���\�{�p��I}��h��ELG.bF�B�RY���9w�}�M5��ahk�5��r�B�m�Mܨ������rѕQ�AT�ohiΒ��R�YC���z�:<ƣ���CAb򐵫��>���۰A�u���K���c$��dTݚ�l��˃�qb݂ۻW�/%B�d��W/n,[8ӑ�!7��=��`����B�Z{�F�Ȥ�ò��s\p���4�=i��ݬ���Oy�8�7c.ܐ�b�w$������)	�Uq.�ξ6�j�-:u*G�.�\.-�z2�A��<��kܮ��,3mq�l�i�p���:n4���*xΫ��ne��{�5�zF*�<#w]��P$Z���v�g��qb4=dK�F,-7�*oD�2-�{3og!i'��#�#�=����(���v�+wk�r��)�w��������-u��AݬZ��O39�nb ����r���b���9�G�p�6}Q��u�r�==��Xȕ��]�8�g��NEN�Mr��9���vt���A���a�>]y�����m5�&Eԥ�+�vi�hΰM�Q����媊��c�z���EdTNUצ�������=�z]�Q�]�O��2�����;<�dV�c2�X�.q���u����OZ��9M₥wu�Zʡ��m����9��1N��'ZE%�ɚ��C��xn�;.+�;�g
X�6
E
���gR���  ��?�|��x�"�/�|U+��	u»e�[�*�>�7�I�5<�Aj��Xh=�ᕻ�Z

�&D���Q�=�4şz��grG�<]�R��/�}m�m��9��Ξ�$'�ztq{�="F�*7�u���xe{���M����y�uv��Ng'��>=�.;c�6��a:X�M�����7�1�FT�Z�\롇��i�Rx�����ˢU���o��xUr��.�RÉTy����������|��U�*�|�|k8Y6z�*����\� �M�W�m�*�z�=Dwr�w��:7�pm/���f���KJ��B����<&�d�b���yUu͇yE���~��ǉ�ޅԢ�����|��ߢoއә]k��U${=��ԣ48=<]�ٴ�Q�|$z�iG��LO.3���0�j�Ӿ��׫զ�n\���?"��]�*�ĸ�$�&����A�/��H���f�߈�O	��_n�c *ߒ��u�;�E'3�~w9��AH�).�w�j+�,7��,e�=���)���N�>�����1�N�u/x�NEnj	N��72��l���N7q�ThC��g��+Tt�Qh�+#L����k���w�YY)��g�uh�	��,N7��M�Cj*~�ճ�v�ڎ����S�l�ʉ�g��U�0ú������]n���T� �n��*��R�r]���"�oP�"jX�Y����#�7kK���@�on�MM�;zp$$i옾�����伹��ߙ�Ł{3�U׫;�L��r���Ks�d��.��/���}��y�~Ӗ	U�u��.J��t^k�����Ǟn��/�oe�4���'���6s����/<w�ỦE�W�%�@�y�7�<���gL�\~;��B]]<ٓ(H�~��:�\f�-�^�Ň%G�6�v2��M�ݏ9��#��v���`��_C�{7���:���Qt�m4z�+���ߓ�w����N�Ρ���z�3Ԋ�Jek<q"���܆گ)���x�Tm�I|����*]>P�1��"Tc����{݆��Lr�껹O����3f��Ɨ���B�VK�Ev���}5o.���v0�Atu�q*���	@�ZMi�:}7¢T�8��޺��G��E���b�
>\��ɚyS���u�]dܷ	�V9^l�����ToҶ��7��u�k:	K.i�ZOv2�7��'ٖ�×ZG�O)�}�ZS�t�M�̶�m� �c6�� �~!$�  Q��n�����S� ���޳z�m��c�c��[Ų9���M����Ļ4>�nj��n�ĺ6�S	�)9�6��.��h��_/y�����]�`�b<�}½�;�H��-��#��9ڌ(�z��h��`uOO����c�A��J���3P���>U9����]gj���#Ÿ�Q=�x�5�P��3�U���\�̼��w�vP�=�n
ܖ�l��
()�֮�)�,�}���g��d�0�Q�̨�+��!�x�v����z6���Ȍ#)7�c��E�S[c$��{mg)7y7��q�%�7Q��}�ݼ�7�g���H�ιhS�&q�o��/f��8���X oUq/S���g�������/˭({1��Z}<6){�F�h=s>q�/Lӎ���R��o�,��n��o���+�~�gܫy�����=�L�b��M���<xT]�v7��9��gF>Ŷ$Ɣ�L⊘��r�T��E�* dR豈��m�*7C�ǈ#g��J�.1�;mU���~�q��ǫ��jT����mGzohi��p%?=�((��z�� �2�����v�K�B�ǻ�(���u�� ˳=��hi��Խ��U!�GJ�QʔD����.�|!C;qT՝���^)�����i�(:�4����p����1�L���fUޅ�&of��á#��8"�;�p�K�7:o������VR���虉�u}����%;ip1�U$e�Ɲ)Έ��ĺ�VB���튣޹���6y���ÑƉ��3
���L��+$ޖ��}��ϗyzLy���䲰̜z��e�zN8\zdp��;=3��,������E_OJ��S\���\����KƦ_���"�]-MW[�K`��#jMM�����e��U��}N���Y�`L;38*���x3�c��M���>�D�����}A�x�+����~Q��#��s7S�C�O����J�_=�t�:���援�=��2R�X9���&֤�F��J��Y~Lׁ�2S�>[�w��63ʺj���h�^�^�@v��,���>��f�s�ʘ�
ƣ�3v+h�W�nV��,g8����wn��%�OSC�;˘���sۜ����7TRy=�Nx"/˧<b�6ww'�9��g.uV��F?^�m�`�������k�E��Q�WOEl&; -3���y'.x�9Q�k>��Y���\�]�D�m�q���˒�U>x�\v_!j���������]�G)�W����+�&p^�Ѩ+
�p�̮
R��z��zN�Wr��o��������p�L]��r���y�{]����OM
��Gؕ���>���_Gx���o�zG�
�mm�S9tׯ�Fh�m:���kJ{z�
Cb�J@��e����Շ�Q��hWNќ�ZϟI�H,�~�˨>��c��}'��E�!av�UE�ϯ��[���#���I�ƻ-�x��T�����V�?G%SQ�>e{Ʈa{W޻��N�_�i
A)J$OMy��{3�,�G���T(-�M�́��>�M� ���qVC����=k�Ut�-SI�+it�n2�G��Ǽ�������Y�X2�ސsaX�i+�=�fX�ô�O���'��V� �k��1�8$�Ȩٞ��Co{�퉩+�{3"3CC,b!����Rf��ǎN��7���KL�5�R�G]�{V�3t�76#t:4���.:�:�ɵ�/�57�_Z�"�em���/鎱>oٛ�p]gS����fY:����eq��ۦ��v�~M�v�?X���~�S2�����Jj��O�Ea���`j����K����x6��h��ՎqWBm��֍�8�q��p�Mjbv�oe��-�œ$q9b���&K�ٮ˂M�"c� f��l�߾���ـ}C�'��xT��R��1l
YӀO�u#o#��`����7Ǩ�>̢k�n�W��S~��֓ȥ�<�r�ƍ�^}+��ߏ?,�q��L����;|oeF[T]J6�
��JqѝlP����k�N�S��N\�rB���(�t���9'����b�o��4���}2�o��ڲeQ��-���^��֭�9�d;��׾��2�1�����ń�Ǉ�y7���B�͕��:-�����Sy���̣^�l1Hv�|nzsrx�9'�I��N��ڟl�=K<�z5_��;��ϧض
��gG�y����2�E�d~w:���W��~Fmχ]�팽ͩS3>���?t��T��#Oy�U�:lr.�����x���k|goz����o�V��u8=�Gx��s9��&�SL��3|�&���޹ƅ�ޮ���O���ϗG��T#����	v��V����>�O���#�s��Hz����m�_���{k�b�ʤ�+� �݊c����:��1�#{4S�uXH��(�[y��k��u�y4Ń9�2D��W3uT�WU��ږV�Ҩ�j��V�RO`n�l �� ��ܰ` m6 �o�����lNS�M.4��kwdʄ�)�5ui�a���r5��2�+�w{0�6	̬�ٜ�[c��Z}��˧��\������=6�(���3�UL�T��{=!��՟s�?��s�]�렧�©��ˊ����-�5]{��ɇ��,�v�}�鲫f�.���QKIgT�'Z	ixu��ISw;o'�}w}���kơ�>�d��%�\��2�<�z�FPul�>� �Y�l�.�e�ǡ��WJ���rD���i�T���}�L��M���K�M)�/�K��i�@���vG�(ܠ)|eA�t���.K���ث����c.Jb��
��b�l�!�7���L��w�,�L�5�>�����`�}�����[�k�S�אַ������"�BG���y����v }���ƽz"�S]��e��yŻy�YVufƅ^'orc5��I�'R���壘1b����9�S��jrsN��4�BV��*�p�Y��i���\��\�|�h�k���������0+�6uό���x;��U��׻��z�;�G��Vd���V	�[��r<]�u�zti�6��ϸ>�u���5{ݘ�v�Afլ^�&X��ט:���y����Q�;w��&�UJ⯜���tBERs{��@��-��\W�jì8�ɽ(+��v]��۳��-�s'
���s*�*�d ŵs�>��^8��s@��)!5��������Nb�{TTi|]]f�k�x�i���4/�����:��T�Abvp\�B���Ov(�8�gb��;�b�Z8�BISԗ�A����f{��|=����,�|W���ݑ����Ԫ��Zg�Tkiz��r����Խ3B�f����踴I]O9�9�����
.�E9�3e���.��!P�p�Qrz&]*�c�{{D�T�Iď�$�Ѩ��zk畃�T�
,==^�9,���K���Q���O
{�ҾU�L�Q�v���wu���3�F�wq݊�vBrDB�������Q�UޫSj�A�=�����q�՗��TV��5E�86N�jr�~�j$n����;�_��5`�JB��;�K�u���h	��R�:ĽD�3nnQ^��WCE�����|X�s>,�]`���j�W!�n3��x�
Kܖ�ή��u�%�M��:uA~�B!�|;�i������F��t�1�A��9�\�+�M�B���U&�Q�vb@���U�{W��o����̮�L�9M�.���]*C�z�gv�-�y�/\�{�F�j>ƻ �:��"cy������1�!�;��ʀ�GT:u:]���C��Q2�N�yN�|韸N�}�v�W�D̘��O���n�bZ���+r�){���'_l�]sy��gH��w�o�,*W:�mvN�t5�x����Ě��S�|;r�xF!�����E��Q�02\���u{x����,o���Zhh��mb�[��^�ǹ�
yZ��ץr��ܡ�{�uG��W�ˬG�O{����".Gםx�/��Ӕ	&�=k�����~�X6;t��� 5?:���#������
̛�'�^�aQI]LK�mN�x����O#]Trrşm1��C��/��V��V͌#8܉�dy�M��7�m.���;'Vl�a6o�VZZXު��;���d	�6��Ks*�o3���\ܱ+У��9���@�]��.D�z\\a��w��+K�b�l�$}�ׇlધ�xL�����#!�#�V��vL�I���Ƭ�S����^�¾�%x���ڻ��0��/�E�Գ���"��z�n[��N]�â��T���sd���PG���)s��alUg'���r�e����7��m�oG4mD��aӘdI��:���o6L�+)#0��ξOb��ưᶷ�N�Hn��$�Ǖ���$;ʹqp�A�o���j���k"�1�28�Ϛg����T�z�%�n��[��u��Ws���#��p�^�p�zfƊ��Y<����{��{X��ek����S�^��B���m/}[ڂ>��2���JMx�K�{g�!�VOY5f�0�ֹ��p2���0�- Jj����^����У�� ���D���5z�9�gLh3�.��E�<�Uy^�#���x�����{b ��gںF��S���C���3F�a=�/qV]gW��O�*�qLKh��(Q�~�D��E8�c:��T�R�Q��?W�y����ch�U�mT{8*F��x��Q�P���t�-�N���X���Vq�2�+�8�
�tis��^.NpW89l�Ъ��~��@?9��O�����w{z��g�Y5�X������N��1������ W�����q��v�^��mR뮕b��nbR�W����/��6;�Ө��M��3m���j�N�(S	ɻL`S+�V����+�~��TD��
�A��v;!�*K�79Z�ԣ�V.u��&2��I���:���A�W/uY�'�x�:�92��Z�f�	ʵ��Ib�{S���*���]e����F�.G@E�O.ah_�.�������u�r���aiʁU�B�i��Ĳ���Mu�(�Mͬ�&���D�˵��
�)��a:�*b!r���f�ޙZ�2�gi���.W���:��	��,�ۿh~���V����A�긆��8/�����6�{1t��H��W�^s�ZxΧ]�w3r%vE"b2uk�4�"������}ݥ�K*��y���-.P���U��}T��Վ�Jf��dr�����Ӵ������flX�!/Q}F��kEҴ'[�s�r�2��?�j�bh�,�z�dy1V���d��r>�7x8\D�8�������)�4N[����2����}�E�ɐYP���	ä���PQ}YXr1�J�����U4f=�a�r��e����y��+zd���kǏ9`Zl�i�Ss�̇Q/J����&ӳ�s4�'��<r��g`� �L^��&�(��9�Y�[���e��U��*�֤?}3��ךC[���V����i��K�5�r��s6EA��^I>좝Sړ��j��6æ��D�0CvIQ�%���r\����zB��SH-g͸���^�x^�Z�k�cU�oQ�gm�쭓9
�q7DS]���=���
��U�U��LVk�UFԘ��[u��)�f.�)���!�2�I��L˱}z��$m%�;��б�x����+�0!>�vi�pA:umΜ;*���q�&��j����W2����^�?�!D~	���=i@��^�9B�X&��r^t۬6)ن�\XҔ&-�����4�\g�L�ܑ1*ڽlt�"ݣ�-u�)rs��:oo�C �� 6&7��cl�m̀    	6�  $�`  	&�m�1�bm� �� Rp�BD�ې    �H�l    d�  @ H  ��  H  ܦ���@%(	�nl�  �l�"̮&�p�Ʋl�L�z����t>�7�u�ù۱m�0(m<�J�˕Z��7MB��vf�Ӷ�T��텏g,X��;����5��L  JdS��3�LKr@���)�C5��l���Үו@�rT����.��{]�p�Ê\,Y�J����[�:1�&�.�KO�"�$F�I�y��۸7uJ}c\��-�;%���.����x�������w[\Y�]E=�Sq*V�.f�).N�죦�j�}")'�WT��D�/����W�ͅ��X�u����Pn�37v�+��Uސ7�0(۹nil(�mS��YN�ISR�n饋-%]R~�x{����m5jN�����J�l�e��I7����)�D�.���Ɛ   �� �  @� ��H��#I������i�	��lUYM�<S��z�M�tf����]@�R�=�;Vכ���"K����/��������UH��t?N�u�N�:����J}����X��tc�W79�֮�s1���{�1>��H�	�Wjn��H�D�{K���(>~�`��v�����,�w�>-U���?>�"�T-��P��Z<3aD�.r�m\�F^7�}�੗G.|th�HN�u�2�wzc�,*�p�u(�N�^s,��Of�s�p� F�rƭ���������-t���-!�f࿨M�+S�SV�i��g��GTqEֈ��ZP��s٫iy�!o��9�W����s9F�QM�a����B���C���B%�$>��:��KYWb*�L��b��Z�9�q3{A�}䗋d�_zMB�3�7ǧ��.�ݏp�k���^��m5$��E(�Oo�7sJ>�;�����'a�˥
��sm����Z�h��������>	�5�us�:15c��};t����E}�_,L���OP
9�uH�������	��7��v"TMyJ哐@랍�拾 �#d���{Ѭ���:����0���ι�[��3���"��lgs��ܽ;�ݐF{�����}:�_�vǲ�};�
��Lvʾ\���Nr��F�
/ڀ~;��xuv7�����,Ko�y��#���mu��|뇴�p���o�hi�2DÜب=�rl8�O_�Cm6b�Jwn%F>�x~Zg�Qv��xjF���&���揵�/��s�:|,{3^`���/ʫ&�o����>���L\�>�i�(`���0�RW}�a���-ϳ��}s�RsP�J$u;�=2}�1a�*<���i���]aTc�k��/}�����P��{ʳo6R�]f�5*VZ��\�m/#��?K��{>u�}���m��,Q��s0�yT�
$xh��,kKY&�z{qE	Jv�g�кϷ̜b7�7���9f�� ��Ѡ��I'z<���^69��Y�]Lv��E�P��{�����y|EΈ��,�5�\�e�s�3�
>&���ґ�J]B�{�>��Sڠw͹ܳ�P�3�U�E*��;<�}�O�yt�;|:`�W�9ntj��N�Vϱn̯<�����qx�mF�i.df.a��Vh�P��:�КNW[k�B8�gF����|n��U(�:�y"�'u�١�
p3#��+�eK��p@��ʅR�ݑ��n���t
Ӄ�!��qG4%�9N��-���,���	G��:;+\���q�ri�CE���������e!�a��tSV�3!gt�V��U�İ�':v�b�N�\�z�2�`�<�ޓ֢�ȝp�����3�lʤ^s̹GF�\�P�j���=^W��g�呧&Q��j������k�̑
jgG��}�e��۰�A�]��f�ɠ�z�#v���/e��.���Giۥ\r�w�YN����Rpk@Ed(��1��*���f����6�M��K��� �ƏY�o�t�W��ՠ���rG�\dÚOH��7v�r䆅���������y9��|d�8�0+w�bj���4�,Æ��4��חq�\��&����L��B��3CD{ӈ�Ӈc �M�_}�(P�K;y}w�I�6&��e���O=6c�sn�u��g�z���n�g�P����nNR<�����������2��t�_B�����������{�;AN�}��;Lc�r�N��YL�\ �G[d�3{T�u�Q'%����l����K�Ǽ�:�j{7o��kĺ��=����H��ŕ�nۮX�Ω��֞Ç�{Kݕ5��	��>"��[T{�O�����qV�fm@P��TnOz�EFc�8�}و�l��q�K����營�ߦ6f2Oc��|���f��轄�ӑr<��H�T&iK>5x��{�O�^���.P�?��G��0�O@H���'yG@֒�R31��IΟT�r],�>���6�H�,�r�+m{fg�x!�����	�˝�������e�-���g|��>~�/�����ǽޘ~���Pf=���r�Qu������1/x�롥6g�צ���B�BS��(tV�g�֪�HH���,##}P"t��Xn���c�4�ct��"C�i��1ܐ�5�Fǔo�L�Z>߹���0��od���ya����<`���#Y<���O�O�e�tK	�1��~�r�&}7���7���dX��=�5\���b����ޓ�̈́���{���h�������s��J"+����<�Dk�{&1X�zU�rnS�p�{βOi�.�9�Y�*r3�Aj�9H�������]�w<��/��˕V��]��su�E�87V�Q1<b�����y/Y�VnL�n�҃ue�T�wtm�L��m��P�M
�  IL�)��!�9قk5�J dF��f�0��r�����A�]���]��dks��0�� B2�B�P������c�M�W���5����"@�sG���	9<�G����#yv�O�~��~���*�]��Ϯ	��/��ğ,4�9�����g�<P�p|��p��J��sG�'؝��V#���q7��5�W�T��Y6 	ݩ/�뽥���, ����V,/ӧX�v[<�:E{&tu���T�/�f5���q%�=�sÜ�ޠ^;L�N꩓N��1�pg	��^ʇ۲���ii���$G���"��Y�.��Ω�+��1ZH��<j���*<t(�]3��tJ�Ar�@�!T7r&�Ĥj�/2c��zr����{_���[2Ql%��oc�G2W��S�6:���0��U.��:���^Z���kpLr�OM\������l�#�C�kN�J��e��s=H�����r�����*��DޮG@��/{�@yy�^Uy�w�H��$�/f�I��k�m��=����Wv#��}�i�'_�ӊ|���?��=y���>;]vԞ�wyp�^y]�#Z��R��X��jů�'�q �5ʩ�`�Q9*����`���p�ϱrT �3`�fYC#7{-�7��ޝ�\����K��(�����eۭ}d\�����Ye����ڋ�f�H:�X�;��?ϡ�
fǽ��4���i�1��)�`��:�]=�����M%Tk3�V�)Ԉ������ʗ�����%�v��4�GV���%�;��3�wZwaIt��"W��@=�>��H�>�t\ɝ�����!���fm �Ď��j�%q�=F)��HY�{A{3�$�q�49A��ۼ�Ƙ<�]�����z�&�����u�w��<�>��0�w�{'��y�c�}���cjk��inٮ��2�U����w56t*d��� pov������w�е�CH'�}���J)��'-{��g*����n�~{1�O5��h�N��B;��dWn{����� 8��mKT(�a��g����͎������9�~�g�k=}��6��}=�� 09�����G�N�Fx��Ѷ��7�V��cDb���t�z�wd�;���=���v6��[��;��M׆�}Q!T'�7��O�Lt:���>��욟n;����r��7>��ИB{Jy@��5��GA�X��r�M�O_�7Ւf���I�u �n��#���x�T�
cq��9G��6Us�#�}nm��:�5�W�g�L��pJSL�j���VU>�s.�ŎV�q���G�`�r᳚�Z"�X0�G��<���A�|�:≕���Y-M�}j�}2~�<˛�:+>6���vVS����}��c�7r��'f�i��(��z+x~{�����x5�_( JN϶%=��Ou?�8��[O��W"�RI��OYq�g�F��r`a�uTc�����#hFm%�RK��pۊ	�6K>"�|�F�0���G���L*�ϥ�Ī3ϧ��TQ��O�����_g�`�χ�����������Vi��y�����^\���8秒怭~��οz��Q���C|���lI8���V�g���4/Ł4U��#��&���Vm-�AOy�xo���02�����(��~3b6av�؛ܓ�-Ț~����fW��H��Ĭ�9/�nh(L���5���5HBb��~c����Ȼ����,g��[�쮥�Vx��<Ch�:�����TH����:�DY�5^1Џ����G�X��:ߠ�)V-;��]�F�5�
�$y�W#.��}�]y������4,��s;]�-P�\���3J��j¼�e�ζ>Ӱvԍ*��jRm�W ��˫�ޡ[�qSs9O{��#L���v�=�̞���G[�v.
���9b��uT�u�j2.ڹ#���ԑ^n73�o�x�<��8* �=�+;=h
�m!8�U�_]�&8X��M�6��T͏P�Q (��'��Z�˕Ӝå��9����^޽�U���j������ɪ���b6o2�}��=�Q�3%6��xC�:��>�{�9FT���#��s~�=��k����*����i��Q����ZQ̟J�����t������>EƼ���K/ol�II��-v���	o�<��{Tܪ���t�]��!���}�@��8����1Cj�������2�����f.��%t��g�}��~�+��� ���>����;܁̗ިz�?Eǘ������-� <��\�P7�	||��_A8(`�H-^5��LW��FA
uޟN�2f/M���\4ކ6�W\�r�z��S�w����ع���S��5�\�?Pg[�l!��d���]u+���J��8�,�6%��s],9�ӌ��5(O�f��{�n��|�=�M�����}/���b�sR�]��| �I 6�  &��Jl @ BD��,����R��5���9���2����d�#�c�=i$-�����n��Lé����N��T1U�' �9 k�;� ?w>"�:&��n;ƕ/i�U���qg����+�`��ytḛ&\�9��Ё~�����ykQ �|ʮ�H��l�������E�9����;{L��(���O���8`�+����*����@{w�i�/�ϲ̎�����騞q�:�li��y�m@|�F�'%���N�=�4�<IJaә��@H��+SP�y�.d�]}NEw��ݶ$K��v"o�\�b���˾��M�����4{�@��F=�ͥu��o����;rp�B�s=�&�s��<�^�d�ճ��T��>����Ȏt)��Q�}29���)@T)Ǳ`j�}ƕz�_+�s���lQ�>�ŻU��<��P����Y��,X�:��>���sU3�.H��B\I�� *��sr�k����X�M��vx˅lFCƗM/�i�qr��杙�ݓj��\���%Zl�F,����ؕl���*�W�>��SëJ��7����w�/�Y3&����+��y�<���,�����وwo�Is����r\!
�C�*<�� �zs.�Z0s94�:^�b�s�[z1jpwv�Y���U���z9�s��X�!Kmiܩ�8k5�1�6.���罫�`^%����� �E�@wR���G�,��U	�����d�^sܗ����9�sD?C�fͣenj;�p�Q����2��+@���7���,�]���~�S~��F�K�Iz5�٘�u��`���y���t�<V��yDc��֭��b��Vc.�����������9K�i���Hp��?L�/��Z��~�8rFGN���^�v���>�oV�}(d���P���(��jG�;Ǹ������Ɂw(�J�>��W��k�(YU1�e?*�i!̃��N�VA�����-\٨�����&x�2�F8���X�#IlMvo����J*��z\�n��ѪH���M7���#�����1F�����oh._D0�����w6���l� ��*�8u�C����z+���>� y�#|F��#� ��E��JE�Z/��O�M�Mj5�4ҍ]�=������^��L4$�tN� -������>1q��Q��&������>���;�A�k}�(�L�|6��Fo���
����uEƤ�ө�;8:�s�t�|:�]�V����d���]<��_앗!���E�// |��XQ	�.�#�orJ�V=�N�lMehn�Z�]6�X�ܮ�f�y�h��+gci_WB������s�dQm-��ktֻH�2�V�q �o�4;F�v��_{2_iL<�ʳxU�9���2�K8>����N�:s��[c1�ͪnl��O��8۝|Z�ƌ��'������/�V���Pw�g�%1��i����7o]#�R�Ǩ@�v�G�%�O����D�VU�!a�n�xؼ�Ei�n�f�s��G�	X,��%Yei̺9���r��e�Ѹ��%��YIRiA�� NX��K�3��ډ��b	�r���a�.R��+��V����l[��p�*�Dsu�u� �z7;��(�Ǟ�K�"v/a�L��� �^�z%]�IB�����i�S��ǜ��X��N^���5D�k����Uð�Y���p�\nce�����G-���2���TPP�ۦ�Q(@Z�u�VA�ҹ��0�K��w��C�0ֻ|�ȳ@u�JHM���.�õa`��^4�X�{�P(b��mq�Ҷ�pHX�����i�'N��zn�|+��ۅ���H�gp�v�Q�0`��h^h�%�ǭ��O��,���MZVU)����%��,gl�=&��ZW`żx��Ы�M[�c1��c|�3d�tH��ӵ8:����s?� ����à�����zn*d\�V�4�C�4,Ξ��(�KC�&U`'�ھ��������t,�Dqk7I �k+3U�66u��8�̛Xk��w����u��Uv��5��뮂��{�-=������S@o2�[�,T���tST}���R�w��xk����&�;p��<��=m�;�] ��rr=���M���lB>��s����wf����)7o��M�'U������S�,ą�Ι1#[�����ko���M��b�`ʴ^ˢ)�m�����;��J��Ɋ]p�,L6z����F�P���J��eM�vZ��xr�����N���C.�iz����]Z2:,#�[���M�9�_&x]�*��z��<O�2s7���Q��=�-��;�vo�D�L`�z�`u��H�PVTaОVvLɱ��T1nH)IW����
�u���i��CYLe��.�U����� =�G���dF��燻7�ty�\�b���J�gR��D���v36fQ��� 	{��l�BqM�No���{�&&fl����`�םլ�1�x=�����
稿tn��R�vU���mm>Զ����HZ��P�N�fP�Y���{���FE��D��wM3��@e/\\f=��b��f�g�]U���U`ezm�,�W�a���	�cn,������2'�z3_�
�oD�OX.�¬���ٻ�komK˧��%��#��L}���y�5��V�w>�"=1CNR����Q�d.ä����⮃[�a��W	R/��_�����M�>�ôK�7&9Z�8�u�L�����Z�)����7�����e�^ږ�齨��/�lY�� f2��ѪIQ�iɵ�&�	\�Pߴ�ޏ]���1�#e�6��;���esV�2]>ȏ`��\�y>�-���;�|��>�����oq�5=wǳ$��R�R�$���s��v�2w�-�|��+.�)�>=�F��k����qUW���=�Y1ذJ%	և�Ua>s4+�RW��7 L�%��Q��n�R�|}�0�.��a��8\c�N:���D#u���^���U>���乆jJT�wR�b��F�T۳Z��C��x��]@��l�&,��[�]O%�nh��~B�%�{�S�Vu͚������>DhTG��|,�������h����`���u:DƉ�\�U�����}��(��U>#>�Rǒ�t��~�����K	C��6���e�t$De�s�0u�f8ۛ�M���h�7mUJ���i9���uC��O�²sL�ߧ:��4�J�/%CG�,H��`����W>�W��](d.��Y�u���҂��0c5c��Q/��>���6���i��#޾�l��g�W��[;�\L�hn�{��_E%y}=���H�{r�b�b��ʵ7�3���,�X�m�\;ھ?qh�;{��HW��G��{I�+�6=�j��z㩓�p}f:;�>�唉+��𪳷�1"<������4����ڇ4>6�U�\|���r5;�}9�m�Ux�$��[PcGuG;�/��/�P�������Ax�������r-�x���u�ƒyZ)�	���j9����=��w��]=&�]������F&�u8dIɭ묠�**aWr_���2�uL��_u����2Z��ɜ3GT3�l�k5B\�� �d�é���;!��C�8� 6�  4�4C8m�$  S)4�u��wxκ�	�ʄS��W�-�5T_K�.��#�3,nY4å�����Km��P䥤W�H>�<�����!7�ק�0�g�{�z� t��g|s�U=c3+fEo�/��2�f�zw�fm�V1_T�T��'	
�B�_A��w���N���xgg5uj�R������B���%K�����}�c�3�Nk�Yʝ`{�˘gݽ��f�H��tL<7h�=ә_wS,���]�՚w�5Q�ï].��9�r�4w�\���Y�8��w��
� Ș:��tO
�J���>5��ө�xd�[<���#�V���`�O�%�����TsK�Zٞ�q>�T'{6���c'�A��K�粞	�$��C��P;6J"�����^ư�Z�E�_3�j���@�ʙ��
�ۚ�g���{��n�ه�(�ۘ>�Y��
��K�
2�[�j߷�����-T�m̉����y�;Wv��;��N����X�с]G�"��qG��Q*v�%�W���z��U8;<�yP����Ƿ˃���q��<���P�0On�~��s���d�pa����e.��N]�6o�v�0�`��݋U�ۜ��A�'R�v���w�L�[�Ja�z$�&�a��N�ď,�V�/�X�r�29��raZ��3+�8����b:�i��/F8�9�����'+�ĶWd�����_����� �5���'�/�iڜ�O<�:,�@��5���dΑ=E��q�o,��V�����{R�������C�6��)b�� �u��bK�wnX[�0{�@Ӫ�݇�B��`γU���+-;;�Ķ'}�<�{~�@Aւ����E�ɬU�~�K�?L�{���u���ޢ��8��N���O����C���z�;�ޱ�U�6W��*" (�7��� ���6�X=�,ǿ�;�z`G�M�7if�
щ�[:K�죜��/g۵c��J�M8~Q��10��M�6��\�"&���i/X��}U�tz~Aq�F
�����FO���W��ɞ]��zGg�������{�4��ϻ��և�����@�<��LK�ۚ^� �S�௾ۿ���Q�u�wJh���+]I�����g,=YC�Z� ��m��ux׈����z�s�x���p�ߢ|ҹ��F!��-�=���6�A媺�OQ��D�U.㡑8X�䡴|�N�f���0)U�΀`.�7�������$�"��Z/�)�t�ڃY@�t�� �\O:ZAꡐ3����u@p�Tμ���׏��Pq�tIƜ��V4�_A�s��D��i|��+��\ri(�9��W�}3������y��&��w�,jjq:/׽_c��+�����B�q:���%�6x�x��:5��&	t��#�h��v���������c7/����9��u�������\\˒7�8�>u��{]�-/�7��Pՙ*��b��i�k�K^Z��:���H�$JA|E:�� ��w��ڍ���j�p�,���M6j���
��q�na˺��]��vוjO��}�XUEn#*�W~�V3�s�>�A�3��E{~���{�r���Ux���g֣��;�CNT���W�P  �����賽�Q���[������&t�Ey�^W���Ǵ�q�	�&:9��PR�>�EiA�m���ۮ.��鹃T��:�{1>yꭁ�I3I���J�(vyyA��r2v[����h�^��Fx*��j��z���i�1�44�Dh����j&���9	����2�Ys�G2l���C��V��h��Ywbp}��Ē��VOU���G�;�jV���n�>*��.%\�V���ck��}#���ݒE�x�H$��RB��K���˘#E����p�}��*V�}��/�G���iR���t��x��}�4-�m'�?uC� �p�^�ݸ/�h���1J,]�=}ZOF�%��T�f�=
W{��Z��H�� ��#��J	�B�Fj��7�A���5ިǊ������٪ө�����L�o��]�t����2R8O���{l�OI�G6>*����`��y�qd��䧋��R/d�x�5���F^ǣ�3�o$=�$c ���Z^���Ѷ�4��������]yz;M���f�����u4.�Ϋ�˺dB���A��(v�/Uc�޻ndSǍ<Es{'Ew��3a�􁱲�NA�2��m��x���ܙ�o��{�\_g�Y��J�����u,^S�::`�鴆�za�zge�߭@�&]F����GTkn*i�\mX�U"n,^��V��Д�K�@������/��}<��h���ʆu(�p��cX�Od�Q�h�{>���y~���\���%��k'#��}�Wh�SX��P�������<W	L����S#���u�:%9f��3�p��C�hf�ߎm �w=�v�p�fS���8�`-�~rb�|3�X$�"JV� P��A�  �"m��
V�OR�[�*�{
Z@㷁�Y���j�qQp��4.̩r��Ox-xU�����s4m?�s�� 3�#�:#;��P��l,:�|�Y;�f;k�R���T[��/*`���3���^�@��x����eT,�����f�m�UH�q\_�=7Z��~�g�w�Rӷ6�����.��xn/�4�rM�9T��\wd������G&m�G��Z�̟�0MhQo�tK>��Hz�ήC2*tE̥���N�Q�r�L�v�r����8^\�n`�eЧd4J�����Խ���}c�R3���c�u\�N��]��Kk��7�7��כ�5�6��ռk��^z��!j�J���O�;G�\Ȯ��|���>ŵ�3��y����/��5 � �6�D�^zu^Z���yůf�y����N]><�#3��}~�k=`���=��cIg�0{N�UK���y�#g�Ur�>H$JG��W��q�������W&d�>]�����t
���g-`����F�J���&���ћ�[��|��
���^O��1���=������ƬD7R�"I��O�pL#i�AC/��-����)�-���^�C1�D�`v8k�E�Mf�ν�D�t�󧹃
$�|�{5�f�<�0�,wit��K�{@w�˲X'�-���+ ��X�m����̕��w��9��m��k��1\>�Θ��s1QH��(��`{��:��Q�Q�/�Ss�����&>�H�z�r��,LW�ss�7�L����:9=�@e{g��x�7W���Qr+�[F���T��5�ʩ�򸿒���Y7���@w�h�qj���w�w�n'c5�&3<�b��]�H�ޞ[��4imJɮډ+�|k�Wm�{aP���kso&��B$Y�舑�9�"̘y�1���B�O�Bpʰ��ږPL��|�j�i n�H�~��;�#���s7�<����ԿT(��ږa��튫J�A��I�l�b �G��Y�y�U��:���TU�(��6�kn#����{(`���Η>fl^�c�Wљ���<���$�Q[�BI"�g�6/�����m]}��b�6v�]��xNV��V��һ��]���2��t�qGz� �;��@����Z W���m�����r�P����듌;�GF�'w>��x��}�"_���7sʤ�*ջ�'?+��o��.lºf�1��:��;�
�>!,��s�p�ˏ/�t�����Fh�w�ׯ�/��y+XZ��rT(�[��S5JYU�K��#v'-̚lc�i�^m��/��ޗw�=�PB��U���{ۯn�8�?Tӽg���s�~��z{2�Ѓ�9��fT�����t+~����c`��C�;�D:��C+º#u�[�Y����}q](���r⌅�ģ�H��h��kLwb��{F}c��>Ͱ�vȣBc�m�*EOP5iG�ˉ(�##�1�ʴ��x�*9��gfx�jB���}*��~�Y��G��b~�	���P�ٟ��h�cS�Ko�H�L��7�8}反�Voՙ��� Ys���['t��(<=6t��L�Y�df�:������g�g������\��_o�#�Æ�8�������YaZɑ;;9\f�j�_����S�ԡ��z6������j��B�}l�91>-�Qn���^�f���3٥�U3B��x��ĴOZ#�U�E}���e(t�De��(}�O�Z/��sLvWz�il)�`m���P��PQ�/*�<��`����e�A�Y0��b͎����Ya�ƫF{��뵏}�9�OL�֜�=�g,|*`o!*��3����ݪJ��k.�B�l��`��X�x�\W&e�k��Q�]�D�;;o&Ci�\a�A��xfgs�s��B���]<!� g��ީ��oE`�B�oʣ�T�p���5ڨ�@ďQ�s�vn��������Q��bG5}R/�sW����)zT�`��H�$�*N�Hs�nZ��G�S�l�B����j�
�0pm�b��Fv���D��ܵ��O�t<G��:��@�Θ��˰8��꺎G�_&g{7	hWNx�Ǿ��k�:+�P<�\��,T���A���Q�G���[~����N�y��Y�f��z}��ҙ�~=��B�E���Z,l�����P���c��lq�A�oo������A��o����Ư�d���T8��#3u_��]y�X�6���Sv��=?N?.�����8��u�6b��%%ݚ��Y��t�W�۸�h����� a�N[��u�>�ޘ���>�ԴTa��X�}����#j\zSH���	.�ʯ�NkL��Q�B��sB��u��L+�0v]<��$����3�ZA���՛v���L)w���]Y&�ö�s���������w 9���I����6Uv�Z]�G.�h�ґa�v6���l
�y�޵�;t��l����}�H.�rӼ����~<��to��t�����Y',���իJ58��,뼫�8�,4+��¥Lu�o��*V�&���,Pa���&�W�u4e���>�'3`����{O�����Tk`[�	M()�Np�b�h+����*�q;$X�Z�{.�Ij+7iH�q�ɽ8�.�.b]IZKŎȭ{�+,�y3�����!	'�IBO��vI ����`I$ ?ْ$		$���HI� ]P@ E�0!@?� ��&��;�HB�_���$�����<=�~���������xxxx{����������������_ş�`i����꠷s�����݊�]�ܫv��Öޝd
�LS6�j�Z�)�����IYɗ%�8��Y��f\eP7I9a��\���kQt(��
mgxλ��#�Wwm��v>�u��(�s�*`����؝K����d�N��mb��)	ڛhd�5�_��ȚPv��̛V��<�B���jFn�� f+����H�r���RcxV�b���ͱ�&b��f�E�L@��(� ��7 ��ɲ�oR���%����b�1�%3^�^⦡�\e�]5�[��p������a����I�N\��efa��i��m���Ml���I�i(�L-4B���n�Um����Cd�݀�օMEbת����-��n� �ݴ�S��%8l��R��z]��?��:*���μ�?��k^lӋo�`�e�Oq$�@�Ƙ���e:T�X�0��kkJý�k�u1i:O��u��w˖k4$t�P:��'6�H���F��WmU�۩�z��5��7"�YL��:t�S�c�.����H�r2R2�b��
ig@͂D4�ܭ[,��H�;h��MW&7x��o3Kƍ�����ƁX+�z�����	��g9����ev�<m;/�Ԭ��i�d�WF�e�)��B��@��{.^�: ګ#\wh�\C����t��*�V��Z�c��E�r��elk���X�t��"��axr�bA
�l#Xj���x��ʔ�ͼ����O�i�������i�\I(к�V�N�lͣ-"��P���(s������}m�+8����;�uַh�b�E���#WK��*��R�KQ;��j�4��ͣSR���=�5J&�+�;jHi�FiZ�����K^�����VSP*�U����&KaLܴ�^RU"4ͲlY�y@���f��֐֍�Tw1�.6�k�����A'a<�<V���ؠ�b�U�D�Yt�ah��[+��Wu�7(hX�VG3X��6q��;��f��9$;��\�����%�X����*�31�+f5�y��!:�0*����L7,i��a�b�J��2�VZ���5F�1�S�d%f���4���R1V�t������� k{gNLr�����n��M�wbz5`gr�\���E�M��lL�ф�ѕ��|�{��Q�]�]�b[x9�ղT�v�'�%@���S�TM�v�m�"[gN�n��nZ�zU�!6�Ŕr�Yt���
���K����7��vʋas A̺M�q��C]��d�Y%��h��v��4aT�65�S����ȧo!I/0t�&f��<Kpfӕ�-�x�I�6�*��I�iN�C�Ÿ�r�Y�]��&,�
v�k��f v�&���T�YY�3����
�B�G7e�0�m�P1[n ��f#o,���;_�T &���գlbn�Y8��Μ��W�k7
�[z�D�tl�w0h2��0ؙpk_�)�L��f`�Ԉ��ׇr�p��i��{f�b���,�/�6��u3]h�tL5��JT�w��m�mۤ�#GN�E��.�ԥՕgi���6�= b����ۧI���՗ �f��]��%�V8k��F��sn�ŶEN���6�X�� xU��hպo��jRP����GK�2��*��-٘� �Wot�;��?m�q����ګJ�z2�3�5��l4���	*hi7{[x�C��jn�
�ꌥ�C����ʩZÛWp�SwP��ST�YP�n5n����F^L��ؼ�6��mVݤ�.�;Ĩ[��Y�Tv�X�TLZ�8��g�m���7���k��u�vi��6�ہ���Mh����f���|�`��Qݘ^Ԕ�dF�e�f�JZdK���D�/5���u��wP��\.�L�ɍ����+5I3e�EF�U�A��
SL����fX���#6�[��E���U��#�6��w�2l�X+	��Zuj�x��I�Aa8Ś�lm��њ�i�ځ<�42 �i�&���O@{+�4ڃm�(,�m���r'�SܹZ�L����FY�W��y�^Z�.�:Z��Atխ�Xn�#7Aڳ�U��,�,D�-6n� �o�����ՠ��X�,L#�7�
��d��	�ջ����5�Zԥ�H"73)˼�;����	�mF�)::�׷�p�����ܙFU�˽�^�˺�`'0n�W���4�ǣ���Sbڼа����X��%�W��\��Ūk��E̒\��ЩvoA�8�^V	��PU��%ӽ�g���E�K�@^Ͱ-~�IfY�z��6l�b��`�h�Yd���,<n�	[���ذ� �m([4T[�/47��G�y�b)¿E���B������Q+^hL�;�=���H�O��֓�h��k(�ݑ� �R��sp�0Z�=���A-[��D�@Cm�Pdwm�5�� Z�V0�*8ubl�r�F�l��X�Ncw"{C2[���,�����r�D=�P�bƫ]�I8H���wu�^�n{2�dV�z���,�
Qղ�ƶ�@���ww)�۬� ��Tґ"V��B)��Y�4�:�	���x�)�����E�"��v��*m��z2S�/��y�k6o8�H�2B@ 	$A�� ��$?�$�R��@�  � BB0�$@	  �!	 ���Đ�!$�ݟ������!$��~������@HBM�o����$�IBO���HBN�a�B��\��5�٣@HBO��! B�  '��_���$!I?���!$��3�xk��������HBL�����Ϥ�!	'�-d�!	'?�����
�2��L#�.� ���9 ��>�<�      @           ��   
      ��@��� @�(@  	@	     P          (  /` )P�    *�<=�i�{Լ͝�Ҙ�����i�y�{I���7�[kW�5J[�ux����w���ݬ�^=H
���k�w)Uch��h0���;c��t��i��z�����}���yW�9�;�U��=i��U {�"�\�X.�ҵ/�l��o�c��� T��    )
�}f���{ޖ�
�X=�s���V������UǄ{��m��u��=���hvŲ�n���w��U����n۞�/_�{ٮ��z�e��u�d��ʐw���˽q��s��R������Z��J� G��Sk��{
^���^����޻�z��  z�	   ()y�[�x==�����qު���mmǩ����=S�޹�S�ػ��&����*�����f�]��ov�s�=�q��{��K�w{6��wt֖��{�R�Y��[q�@W��R���t����%������n[���py P�@    B��ڵ�=��5\vꕧUS�w��5��@��OZ��{��뭫[������޵*x� *�*��ʽ5{�:�s���gT�N;uMm�	Vy�绽�U]랽Koz��i��zԽ节wz�G��J�W�^󺗬��׫Q�  z�$     �[�����)N�t^��wzگ=�6T��޽V�z�*�{����j����度�{�T
sשU�]ޭ��wzӖ��۫¯=����*@���S�nU)�{{�+[��긇u�x�B��R����5�g�y^�Ϊ���U�>  �O��R��0 ��1JUF@  T����Ja�    ��UI1SJ   T��j��UH   	H@�MQ�M=@a2x��>}�������������=|�~z�׿^ �(��u��J�(��(�?Ҡ� �A@��DD�aA@�
"��"������-!�P�BEB���äJ��mAJ�4 U�A5T�jٿ���0ӉJ�lji,��m�$��J���	IM!\����ATH�QM1,��GKM!H��Z���IEP{�AEHPP=IN�5���PW1�	l�o��hJ h�
�T�s&���B�D�HBP4�@�̩UC�1	'69�4�4V�b�J"
����:*(�'-���)H�!BD�2�1STD�h�Q[f���1"�%Q1�m�*i��&���琔CRܰ-%%S�MDT�Z��Zj9b���*������ib()���QQ�%��@��f�B$�qpMh�d"v���QpG{JD�����ruJcN6�*I�� р~[��8$��H��b6��8d���Z��&��Q=ZB�h�SBPDr5H4P�Q4�)A�J��业l!��✁�(B�Y�*�hJ��h4RQ�@ـ��TQDH�B���<�V!�;���2�EG6Z
uJ��K�)������b(Z�(�e��Y*&�DIIJЭA2�u"qi�I��Ҟ�IDQ �4�T�%>B�hy��<���L3*�5M�"�mQ̛N&GAE0[b`��J��$UTΪ���D9
�:M5MR��!H�
�P��[ |���*(i�."�I������"�A�' �T�3UHiW�	�P Q��-*P���9R!H�y�


��(N�!KHR�ް��R���ZQ�����������{��/O��`�ۧ-S��8pAz�ҵk1���7bdۡZ���'�޿kHߥ��wb9���DQ��v+���A��yl��SM�h4&��[�#ݪj��#�È!�b_WP�=U�`��{�1Ը����>�=�W}{��yh-�.���yq:��q��iO���h���=t]�RoV*�Н�|����^m�G�cY�(伄��5շ3��.�Q{��GV)��T���� ���w�&��tu=cP���GW9N���>F�j}lU]��f�s� N�%���$ $����jK���)4{�*�R��۪��m�(��U{�M|��1T�����~�ʛ�!�F���Wy�9.T��EEy�<�.r�QTG�i}H�!4'p�BR=]������	�%-응�N���~��|��׾̢z���@�DR����(y*z��^��F�4��/!qTm�"��M,UKA����:��#c�2%�T*�����KDm��,�ըֈ�b1�����F�-��D�("V� ��((��"�:�b#IIAN�ZNB
9j-iF�t%С�E��]��˸OQڧv����@�J:DY���T��F�iV�4fJj$)�:{�ܲV�J)�[KRX��(�P�
*�d4N�h6�Qlm�P��ڨƌ���Mg��58шm����:CM/!8E!HR�Ҕ�6	e� �j����"(Rf"�婨��D@P<��xj j���AdЁI��=Hhl���,���DSA60V�"9�QSʲf�ETDF�)Ӥm�r��b��PN�g����;����(j�5M�R'Q�)j��ꄣI�����l�W.O@Z�@m��t@P�P����� �Ɗ�*��^J� 	:�t����Y�iI�V�q�b`���)�B�i�P�	�h�C�
�jTN��F��)IU@PD�B�'�\�4+E#E��R��*�M�Z�l%MT4���.��I�3b��1�1��裸F�bZ�H�LICU �B(Ҵ:CBQ5��J	�).�p
H����
��6�ZJ;b�Jr9m:U���Li�4'��\��@`����!ITu%mY����JD�'�D3+C�A:�ᔤ���S�y� �p�'�T�#��*r@:�] �B��7��T�������G�NsHX�B�CE�1�GY��Tղb��a��md��4�$MN�O#��E�.������*
)
^K��"����4���*�f�	KԸ���D�QlLN�cgXъU-m�F5��^�8\v,Q[���f�N$

4�.lU��F5h�M'����6���"��V��;[e�1���ɂ�u�L�0l��[����6�8SAI�4)5"S�b�MLR,�;j��I�����Rna4�SDEP�L5D���D�'CB���(��h�cKlP<���F�`�h��m�lF�*[m�A�!H!�.�j
�,m�fճ�(�F�PQ��gUE5QUD�u�m�TimWx�"��$R:t���4%����C��m�)v0H�Y�F�$C�5���;��&��қ�� R�z��#�,k� #d�c44�"�e(#0a�^�JM ��R�Z%��y�rِ������Q�/6j�(�!��䉹�I�������כ�E+�d�V�H�jڜAE��i�`���MPL���3HU3L ��i!����b���(Ji�B���u*p�NÉuN���j���5D��R4G�~$~&ֹ��+ĞPA�� m�b�*3�Ϡ�;��y��r!�;hNL�x왻pS�L�h�r����k,ms��!�8ը��!�s�ޭ��W�5�N�<]Js.�ܸ9�jxz��ܚ�/lm9��]��qەNbCc��Z���v^v�!��)�l"�1���n����P�L�bюl`�Ͻ��aUT\�7   P*����  [j��� � �
� �Gp,����*�@ � �Ski��	Z�  P�*�*�YV�  *�[l�U�hw  *�J�T  �QTR�
�m�Ue U���R�m�UU.핲*��     
� ��Թ���F� P���Ҩ�m� PUQ�TT�  �  �`
�ll  `�4X%Z�UU����q���9� �m�B�{b�W�)�       6Ŷ�W��E��  T�S������ � OX�Ѹ� 
���Cb��M� ��l���n�U   U �8|�� 
��{<���� ���mV�B��*�l� l[h�eUc*^Z�RS��`
H�b����    @�P    ?��_�l�@  ����\�ݪ�c6�-��U�Pp�U [j� C��V��@   �      *�UV� �{��� ��� 
�  .` �d    U*��U�lG�  �AV��T@6¨��̦̊�R涶*�@�   �
�� U  ¥�ʀ
�   Skj�ujR� �   Uf�wYܷ����Rr̬{      m�         6�J� �l  *��    �
l  *�  �sTU�*��}�ԪU �     P��%[ePU6@ ;�d
�      T       �      @ �    ��@   
��  *�   *��� *�@U ��T
�T
� T  TP@     *�U�   *�  V^�j�*�U �J��Cl
�6m~��U,��B�w �� U c��狗�eV�\K�9��� �U&m��wU2h���ѽn���ηncw�         �       �� *��ch�7�,�`:���ם�뵽nyw           U�]=n�ou�k{o�>��	���i�(ٝURl��pv�A*h"^�v��[` �UR��PE� fڪ  UB�*����� �+;���̠�A�UUTT@  [  �	�cn:B�I��\=J*D��(`�݃w�w7�ݻ��� 6�Ϋr�r���;��Rej���������k���ں���Pp���<�UR��  �  *�3l�+(  �V啙*�e
�� ��f�{�-�mU� آ� �jޕߪ���:�Fԯ�����V FN`ʨY�h[j���*�m�EP�ݕ��6z7�t̂����1��*�W�O�����=���� R�pU�*�*��U
�V�  �UAT �   P  T��Sl  ���1@�E��؜]�� �cl�ujqR���+%w@�T*��suɪ�wr� *���T��Jy]�j�ٴ�L�2��3�	꧜�}n.��>�V��oj�1q��1�k���i@$����ܵ���N�v��w2�&G��m�\��-T {z[.7U��6:���#n�㍽��g�3�k��� 6�qi2��on����A\��ݱ�v�GM�t󩗖g�'|쒞#�w�ˠ(�v�d*��6-�w�y���n�#��*���Y9v�����UI��@�YX�O!4��V�zggWFۣ���-�CN�gsӄ�&Z�R�3�;�M���Um�qU�vlQ�=��,���S�2  
�6ӎ겁T
���z�];�M�s?-������m����j�P���jTZM���T��es[m�h m�d�U����eAre3�\K`��
��Yඈ�t�1U^�(ѻ95���kmskP�"upB�PVK�ȁ1M��ų*ʦ���t�6XX�"f�(ә�u���� 1�6�2{N1�/&<�[тY�tұD�nY�9`u٫j�ܑ=��U��`�L�v�c[��������8�C�/R�T�lx��@#�bc&��햰�n���4��q���֨�<1��a'�rs��`
�J���+��Wg{%�t��q�v[&��U���K,*�+v�;�VWccg9qf��eu���U�1�6�&Lō��-fڡ��ݴ��T��أh��lv�e]�]�(�$feM��:�s����!˶8�*�;*�<:�@\�,���QV�t�  j���m�ر�Y/u�`���<�9 e���I` `�ʪ�U*���8�
��� TpP �*�;��  m�`l�m�;Z����  k�� �  ;��    �   �Uz���}|    �r;� � U*����� ��z;s��� ���o��|`��+Ry���m����     UU   �� +2�     T                                 �   P�� �  Y@ ��U v�
iP�jW-� [�`  �` l�    f�P *]�Su�Jۻ�ki�T  
� P*��^��U��ֿ��o��R���*� Um�d  
l*����  P   Yۻ��  �           PU �  U   �        � [�[ U   
� +��9��m@�/T������       U  �C��o��Vֹ�������[��F�*�R� lP*�T*��@�6�M�d�T �  ;���
l
�
��ΰ
�   *�� U�;������\B��R��&H.Zd�@`u���L��=��                ؽ           *�           l<   U                   T     �ܪ �\Ͳ�T�    U  P    P           z�            �        U  �@                    m�N�P
��V��    *� ;�  U�� e 6͚� 
�UVڪ�TUP   @R�qU[��wu�r�@  V[h[-�TlUe�  ?���          @    U@���@ 6�Wue;���   T2 U�R�P ��    T  8*   B�m�[j
�     �m� �>                  R�T�P                        uh   ��         � @  �| �;�J��                        U              U              
�         ��          �  N          �m�           �   � @   ۻ           ����U� �6� *�pw;�ǀm�P *�@x�PT�T�� 
�R�T*n*�PR� �md�  �T�u��ʻ��         B� ���FE� *Ҡ  ������� p�j�UW]�U^��vq��  ��R����u�ce�  +�mޝ����7               
��          ���m�ou����xU *T��*T{�fP� l \���Sl<w%h-� *�         1�;]����W�T      R�       ��T 
�� `�   	�݀����V��qR#N)��w{���{���DQ�� � o�����~���o��K��Y@ -�TT��J� 
�P� ,�* U@6R���Gp0��ջ� l[j���Uo *�:�l����첂p6 �� lN�   +5�*T�Gpì
�UC����n  �T ��@ �T�     � T�Ql�
�  .	���@Se�F44��,�m P /v�g� 
�5�w6�ا�g�*�PUP[d�U�����6\pX�W-]�9�e��*�TΩ�U����6���p��W����UR��@��w[.��@���f���K�ˎ'���-��n�� �ڗ���k�5�(�M�(���g��S����%�˸-����]���W,*fv���;f��UZ̶�i*��7�Al'Y��vw�F��\���\�n��.���Gm�g-��\�� J������\f����g/��m��Wv$;v%ZVYUQ©�6�얖Ul�P9jQJw���۽v���P 
�       @�P 7Z�[*� �<�V �EP�@A�U  P  Y@7V�PLқ�؅P,1PY�E�� 
��ˎ��P  P    �     6�mT*��� �    �    -�@
��Y���aT��@�Ͱ   *�d�J���
�[@
��  ��    `� P+)�     *�T  *�� 
�� 0 �
�  �5H
�[��T["�m� ��l�wwQκR�~�  T o*�*�2���  ��m�  %V�����>����{�����{���o����R��UB�f�)�Y+T��J�q���6ʻv�l UX�t�:TڮR�"�T6y��Q ��2O�`���Mm���]�hc#��$�I�[e�+���wm��r�� ʫl�;�8�sgT�(j�m;���6��UT ��^�`T�Sa� ,�`
�E�[hV�ͻ��*�ٲn�j�{�<
�DۃeAyݷoq�vyCo"
�UUP yU�c�ʢ�����O��*�?����60��B�B�>��g�R��}d���R�ZB8q��F&�m#�R��g������.���P� c:igڇ�	��q�����Kb��JY����7�q�g'���̗�P����ZE�9h��C�=u|З,F%�F-ϦY���^�3҆j���p��L9=X��6j��:"V��{��p�L�UZ���?��Iqև��Q�����d)fX��ZDс��l���ΪK+�P&^j���c��c�U���h8jIˍ�j�ml�V����d��c!J��&5�{ܼ�ܗ�����3�O��-5h?�]oŵ��GU�Gf�c��^[m�!���*�t���	��[b�iHZRA@�Z�,�sM�*�7���* Ycr�U�ۜ�뚞�'>��(R�
D��͘sP�g����af����.{��?�ZEL��D,�ZF��"�^���%��,�+��x�f0�o��/��35	z�Rz��x��v�L<�{�Nh��MP�ŕ�"�+|;�z!f��VB0��3LUhYv�ϩ[8|��T|���ZgJ�-wU@��;��ܴk����4m҇L���+��XZ�X&�R�_�J6�`�f��B��V����Y����D�#}(Yb�u��t:v}57�I��Е��EW>�z֔r�p\�Yd{�E���C�njP�,�!gmS�.�8`3���ᮥER�-�fV"�7�L�6Ξl��ˈY�¦�c#+9�z�g��^�=�(�\BmuL�,�=�|��
�U��II�{���Oޭ(�vw:�.�f�ӕ�i�M2`�z��F����^���Q�h��	�Tn&��(��\v9�F�Zaс�p�-���T#O��k\�!T�7O=��$��[%��s�a8�޻sv�omղ�{5�K2 (��u���Q�KW~'��l�y䶅��H�qlgM=�3!9Zip���4-8�e�5��h���-mh��o�٩ٛ���s�7	���7Ҏ!t�5Օ�i�M2`�_'����qD�8#������D{�6`��gY��\v9�E��0_��<��ߍ�z:������X�p%a �2]�J�,{ ���X��=���(�-p��]Xv�=��s�=��L���!J(*�U�9�F��y�W�Gr��V�)�C��׌��(��Y�0�!�9#��4lMU]Fc��1Tn=J��Z�]�^�*ke@��2�<Є!q�#$ġfE�x�-,>"�q��f��Yf�Fv��\a�S�X���Q��v���V���O|ng���\�"��z���9k��9{a��H�qtt���n�[q�Tj��,�n��7;>�ϟc�x���X�['�w+>]Z_-!�6)�T0��t�����-Đe�Ƙ^���0�����-��VYi|Yiв���x��Ο�c�>j�.֐��URCȧ-��qi|���g$v�rr��oUa/n����t���2�l�s���g#��ݧ�d�m�UQT�6�m�nr�%
ly��lC]��@ ��N��D�+o.���{4��*�$ό���W�p��ǭ��-�zMm�L�2�5Ƣe�]�����wɹ�bFsR�؝��ݶ  �fU�6� ;��Gv2��;��qT
�J�[lV� m�lY@� �*���C����h�Wp� �����m�l��Ǻ�B,�-7]׹��˖�M��q���u��G�ZѲ\�W'驜�e����}�Ϗ��D(�\Bmu[���=��ӗz=Ó�ֺ�Ze��mX(���X�t��}<�S=���=�9�뽳_L��n3������EWC�]�?�_���C��r�/T)�8e�UҴ��3q=:I}���,�	6�Q��V	�nm;s��f�O=��J@rh�"6FV����(��ck��M��#�+4��4"I�I�<h�j�m�Xxݔ!��B0����i��!4m3���w���3�����UJ�c
֑�Y0��u�8�I	ԂF��T�UR���$��ƒ#P6ہ�S���8l�][8�!�
xN,��Bs��4���]n���!�ǎbm�P����܍�Sp��6F>����2��my4�2��_!���ˢ��E���d?."�W�ܬ��V��	FFܒ���p����]ZY�Ȝ9=x��(�h���i�M�6��6p��m��m@�0�#Q�!'Mܬ���'sx�,�	�h�4(�����{Et
���p��k�I�(�m��r:�* �����-i��C˨x�ZF�%@Y�9�F���#��Oim�2��k��iݻk�D8s��� �]�Pb� ����lnwv�A���\��x�y5�/�}^�N�ިw�Zv#�3��מ3$,�K�������ńG��m��:��ވG�$��kB������O�1��#b�(L�U��,#1n%��k�N3��#d�畑��P�Z���7B��M����j��{��d��l����,�]v�wn\UZ�kH��R��^�z�A���ǧ�,Tp��P�Zg-�C�x&OVo4=�Q�B���\��
6�!%+sў������Y��!谓1x����]�W��NG��ΙgSs/Sv�b�KV���v��g�)���G�����N�{`9l�%T� ���G<��v{/|��-�G�X���B���+J���TA���8���6F<6�lx�������+�VB�;53�2��wm�c5<x�vب[�f/*UÇ�n�u,;kA�f�6�0���ہ'YH3Qi��4æ��0m_+��a�N���q�+�j�içK�n�ڎE"��~���4|=�&�p�yn�ut_,:Y�u�L豝&��ە�L�{m������=���n6���#�8b��qii�ρ�DxjfMKn:�0���e!�Qv���um���֙o~��}�e�T���ԛL݋�m���� [VPVBeZ��V *��=;لm��Q8��3}+�����Cf,��&��z�,���9�>���D\B��R-��f��s��gb�(eh�a�3ʄ͌4��'u�\��h��ބ��$j�jc�[������3N�di�&SE���F�Y�mVB0���T]��1�[l�*�[E	R�}5>�O9�����L�t۷Ս����,>�雯_��u��M�$a�$��*gY5L߈g�HMcA�
�Z�CE�!��7�	���Q��\��RII7$v6� N��wvw^�ݨUx��G�lm��p�  Ym���!5G��U� �����u鶕 )Ǖ��#�2D�2A	4��'=�s>��+�oagnv�4�:T  ��J�[�nj���*;�[`m�@�*���< j� ;�U � �e��Pq_��m��ڨ^�6�v�d��i#��`�3&�V�a�]&�WuU�˚)�U *!��TZ*���?��$��m|d#M4F���n,#ƙ:�5^�*j[q�V�El�1mD��Uw���ܤ^�~̙ɭ�۷��H3Q��gL�����yA2(���h�%5ㄜ>"�y�7h֐�:)��4(�G�w�;Y�Dg*�^�m�m���;���f�S���U���(�OE���4x��+{�<}M�-�υ.>�Ar�+[nH�,��m��f�N��뷱a��܅��Q�����7S:��4��:E��S�{nGqn6�gm9v�t%����i^���"�%��b�l�-,J &x��=�{�[�|�~�9k�q�'ǌ<в�;�[!��Eֺ9�C��lo�0���m��1��.�~�|����2�*��5.�˞qW^B/P����	vC9<C���P�Qi���и���%����3f@r�J�(����1��#��<Bȼ��,��	Ֆ��C<s]�fӅ�\�)�GaH9.��Zs5�6Y�Pǎ�Ƶ2<Y%�#�}D�0��޾^�%)���nFCNo[�YD����X^�V<}v⬾�)�L9�y����>�~�8UU8�5��5G�����;��(�J
�T�U@E
��K56Đ���M弶�-���"���Fό�!��B�8E�)^�p���2�	Q|ĉ$���4F�;��+6C,�ɰ^�8l���a�|N�¼��tJ��,����8��y{�o��������^�|<���EЂ ��^{��u��=����=ʇp z��#�>z�	�V�S��"'��� ������@>]B�C���M��|�[�Q����G䜽���������4�f�m�g9��k��Ƨ�u�=kN��\�v>�y}��uϿNv��~������y���o����Q�O��.�i~N�������+����mι��ι�]v%�4�I�>�9箹	�~K���z��/2i{�	�a(���e�i�>N��a(����K�E��ӷ�O�	GpO�h/��'�(z��\݇�t{��]`�3��R���1!�+��8�qDDf8�v�;�>I�;�	�a(����7}&���'݄���Ԛ����o��6�PK�4���B}�<��ģ���4�Оl�����y�[&����O{	G�%�=�UO�՚^eZ���]�j�j�X���\UGq����URZ���6�Ȧ�Z)F��7w~o��{}�_���^y˧��_|�Q�I�M������{݉G�%̚_�g���%���~;�>ɠ���O�	G���ÿ��9�{�/���'�����?�"��}^���&�fF�����>l%@i9&��Y��'N���J>����4�Нl%>]��u'ri{�<�����pNu_:�v���O6�r<�������ԇ�N^H���/���Ͷ���\�\�I	���@@���?Y�>�����G�����y��g�O��4}��{�y���9���G�'Ri|�<��|��a������&��:c��%��$}���	��� ,�����y}޽y��{��|�M����Q�'$�z�^y˿����@z�	��޻�pNI����>�9���	�^��q����"?28��?H~� W�m�ƒq��KG7:�i���<��`~H���ϗ;����O����O�_O��Ο��������[n�:��޽`{�{�tH{������7w�����UQ���R�U)Q��Sr���E�؀�˺p `�U����T2+* +m���~~�Q��������9�J=�i9&��Y�'�	G>|�y���M����0�rI�^w�u?`��!>�% 4�������瞾ohW��Rw&��y�%���ή;��m�]l��S���H���������$}����=X�<����}��}�M�t'�z���N���;������Q�~��>ɠ=ΐ�~���ϟ��S���}@����έ���[t��Gh��@�#��y�~�����#��r��w�����Yw^p{��d�������9'�4���!=�7޾�o߻�y^����H���Ľ�h�!�q�	N
� q���-!�3�.�߿7]�C��Q�����(~��_K�(���:�K���̈́��~�|���&��t'ͿHh���?k߮��z� 9�����z�@~���_�Z�V��~{�w��;ݷ>��pu��~���~����y&��:��Q�����>O�9/�3�O�	G�'�d�{�����Q���u�����.�}��>�i>ɠ=΄���9�� *;u���A��S�FU������lv��  � �(�򇻼6������"�6j��[hnնBQ���Ú"x�n��k�/E����Z]`ծ����vѳ�p  ���l[   �s
�sc���m�ܪ�UTeJ� 
� ;�Pp *��U��v��Kg�������Wr��a-؉p�p��S��@��N��L�UR��VN6������i��o���Rw&���<����z�y��䟤�΄���y��<;������｣��l%`4����>}���o��6�]���%�9<�י�'~��|���O$��Bz�J=�~��d�b���G?;��{������<����{��y�}���h��$-����$�ɥ����v�	�a(�I�M�t?|�Mؔ{��(�������#�E�������?�@�jBd�FKS��{�W��;�.�t�W�/e�6dZh�bXӖ��|�Hy!���û����7��}}��S�X{�9˳����Q�I�\�׾� 9:�oWؔ|���Y4���!<�J<����$�&��t!��=�9%��Ͻn�K��y	��Q� #�x�T��������,�v�O#ap6�6�?G?������Q���>���$�d���<������z�I���~;M�t'�	G��Iu�K����\����Q�����(~��_K�����rK��_��K��Q�_7��s����Mg����˽ɷ]�Jyf�U�UwpT��UUP @.5I���s�κ��`y'�4��>l%�`9'�z�t�_���O�	G�'�4}|������Q��$�ɥ���y��ģ���4�Оl�:�}�=A䗬�_^g��6���/<J0c� f�~��2?XJ>~�rK��_�G�r����������}X�ֹ�:=����G�9�t$s�Ͻv%��9%�M/���O6�;��};�>ɠ;�	�a(��|��,w���9�Bw��|�'�ra3S?��v�V%�cb#U����9��טIu�C����	�����WbQ�I���y	�a(�����/2i|�<����{��䞻��~;M�t'�	G��Iu�ߧ�z:O�:����L4K.4��C$���Uz�V�?���=�}O�>6{-���B�Z��V�pȸ�鞔���5�ˎ����>��{Ǽx�BYnqx�/����;����Nt����?pfo�s����C�Qb6�[F�j�[Sv��HQ�L�]�V�� wR���@R�e-��=��������*W^���B�r�"��q��ސRz�_gXc��U�������q�є6�h� RG��+�{���Z�^s,��	Նj��<^�ohdf�:G�����!2�'�%��x�G�à�E��$�tڷD�Sm���~.!f!>7x���[h���k����9޶����!��]-z��B���R�x�g��(��4�rm�-�cm�P��a�>������՟�P�>�$t,��l��׌�ɑ��'V[�^S��PmN��e�R�l^��$x��	��1(+mUUU�1�v(��ű8X�c�����}���}��4t�:I�^#ut19�,��]�Q�2Dc��\E8����|+<���Ķ��gO��vl#i
8T�<|F�w3���}"2*�m�&:��N��t%@a�B����E�Yme!Y�E����&�����TLJ$i���.��~�J�h;9�"�zA/N4K�X�D�g�>T}�!����ID�D��H�Ӥ.Uhg*,�
��1�Y��"��Z|��o���p��T+	j40m��I-v���;��ela�3T�Ew1*+�*�nݴ�t��ϘbT9�i�����f!/Ck,J�G�-"EG�?/��|D<t��N
���XC��̌a��E5j�uWz��'W��S?�jnl{ǱY�A�3��?|����}�yn(D>�/�a�
��,���s>�Y��+���
3eEF�UX}�c3"�X�խ�4��;���"�(	7�wz��T�ww�w3U*�8d\CfЗ�-2��2--'��mVF{�w�%,FV��J�x�����מ3�#�Q'����C����>u���F������M��Ϸ���Ut�6ܒITP[z�uOWt*��l��45ʬ[    ;�wD�--V�ě����&�C�����o\���Wv��v*kc��9��&[����]�m����u�wd�oN+�z�  uk�֡TTm��UQK�ݣl�;��R�Fڲ�J�ld ` ;��UQTU����@/U������dηE<�w�w}��y�;�t^�HUܲۻ@�
�[iV� B2�eʔ�ULn^zi;3�ğ���(f
��3�W��ڧʋ�yQ������>�@�nF����D����?�|k���I���0�!�6m	d��L�����_��!G�I[B@ێI%�}�x����?����|�,d�?Z�Ay|O������~>?O��~���_Im��e'"J��6�ڑｼ�y��)O=-��&�m�lڍ2���ȓ�t��UQ"�]��)��p�A�ȇR�t<�zE�����F~<h��j|i
�����;?N<��n1V�i������[�e5�]W�r̫�+���V�U^�WI�eS���PZѱ¹?~73���d��^#/�Kڀ��-a
uמ3S#�C�L嚄��8��h�j�UUITwě������X^��0{�"mI�U����-���#����;U�d�Z�-��26K�ʪ�e_���n�]O�
�f�Gyh�Aj��oSZ�Yh3qVV�67Uńk7�E��J��9�&h_���f:��?��S�7�f����qp�������܃?5^A�+^J��\G�{�a��0�I$d��뎈��WWc�"Z�_|����7I}�q�.|li�P�a>M/�����R?���9���͌����[{͆�ۨp�Y��� �ή�s7�ܭ�q��lݑgN��C9z*!����L�r�n�6ʲ�oSZ�|����>�� ~�R�����������a�C��Zd3�%@dZG�{0����0���V��z(��9�ȗ���@q�Ij�k�����vf�zx��dCHG�'V���[w��R��ͯ�g����9C�����J�(�nH-�!����Y~�W���;X�m
)�!Q���E���p�R�,ջ�1A1�l��9O΢���v�^�4�L˯փ�cZG4(ݖ��c���B�f�@R��7M;�b�ό�.����RN���J��4��cY�N�d�U�WNt�u90���Y�L֏F�iش�Eۓk|F�rЀ̕�/�Ev�����Ȇ�pH�Q�BV7KH����y ���{>W���R���轙勞�I�����I��u�ԏ}�^����}���,��(����������{ܹ��Yo߾o�,[V�ZY*9����ۤ>��y�B�|��O�}����1JӍi���}��Z�Q�Q�<�)"�-�C$��C�YfM�Hx�jd6�P���V�d{PfN5��`Fz������m����իT�^��Lv��.����7n�m�� +sVͭ���Ʌl��jB���������G���>"}_5]/���/���a������!�W+��!Ʈ{�AfF�,�!��dw�3 ���qg�����Q����v�K^#�B\���ig���kl��Z+E��3z��n}XI�~���Zh˃�k�CD6�fw���˯{���<r��kH���T��:����[�΋�߰w�2R�=����7��J��ܬ���E"X�%2[�HQ1B˥����Ϗr�;Pg�_?����m��/�v���G�ï�����o����ڨP*iQ��#�c߯����G���9
Q�A;�R��D�
i�P����"�EҠ��ϹO�"��H�>�(� �������ﯯ���Q�����j���B���P)�6��بm��6�  6��`��P��M�H���z�*l��=l��T  
��T*�n��!� � �*��@ +(  U�.�  -�*��j�[j 
�
�� 7���  mP�
� *U 6��  � �T �   �      ����*�ed��[�{�N�]�    ���Ͷ� �Z������ʠ��n%R�KdV��xs����@��(	�5UU*��B�AYM��N� 6ZC�Ayj���Z l     �ESתVJ���W��ю�&��E�H�Y��f�Ɍ�5�u��`ݍ[�|���Ɩ�R�Q���� 8�MAYPR�J��\�2T:�� �1��P��Źv�ԉq�T�C�Q˵[s��^v�1ͮ����\�]�'mir�I A#��R-�-����	�j�Cʦ�M��l��}�}�ک�z�ܩ��;�-��+(
������{�6- �P        *�*��WX@Ul���P�c  UP]�      U��
�S��l�  mu�����S�U��[� �l�J�3��@  U    �     
���>    <         *�U@@)�� -�T �*�  U�T*� d� B�T      5�    @� 
� �     @ |       � � � � ]HT�T[+�Tͪ�PmL  T�ڠ�l����:��  @|��6ت�3j7]�  k6�  T��U�ۥ�� 
�e�v2�R1�Z����w�����U
�  *��{�k�zBĮ�Vն֞>�7�|'B�-HR�zd��%g]P���.����4u':��1ݤ�`zZ\� �CM���P �l�����V�붩���;��l�l�� �� �T�P m� � �J��*�U[� �U]�z�ّT�9sS���[�MKF�3;Q���e��dm�k`����Ɵ�Њ7q7����ǧ���ڞu>�������C�A�`ĸ�ʮH�#�����_s|�1l�W-��I۽iHć$g����[h�_mW$o�߅��IjF��5�Fk~�'�?$M!h�_+�sFeΤl�����	I���P+m�V���$��6��3��&���H�F��Ƈ%����ѓEz��r�䍤IÍ���^Y�W��OP�x�|�P"�m�F���-;~˭k�}��z�V��{�wy���Ʌ?7�'����"H�*	�GU�(���&����f���r"�"�����}�da}5�u���|Ѥ����/��#�l������~7��H���Ϊ0c�+�bZ��)Bc��UF�W3��V�p�*��x��*��uU@U*ʀ�0�����V�}	�[#�u�n�������I���>�&ʴ�#����4���*���"R�dH�E�9#�v��RCmHc����!�א��|�V�׷����"���&|׈��#��ե��ԃ�=[�#�F���(�y+9	Hn��s�r{Ӽ���)b���'>N��#��%Ag͟�l�*N>u�1#����.U�D�#X_p�yrB��l�6j��@�n�r4�m��1��rT���~�]���=��u���5��/�6J?$m!�^�g8�W֎��G�Ö|�<���=�ē��jI$P�S5��~�:�p�o!���frqyQ=+uB�#<��7�~��gu�h�K���p��q��	)jG1��j�gP�7����V�m�w@ Sm�Tڅ5kiVA٧��IK�d��[����*VI�G����%�6{�ɢ�ԏ�U�g�<��E���tsd�\��;ؖ�e3o�.Avyc��g9���z3\��G�8��y��w���l�+|eCG�4��o1��l�h���8	����	�rض,q��!8��l�͓E]�ʫ�1#�61#+����h�?��_�Q#�%��v~HZ[�g1�j��C\�K�|��[��~�2�[j1[�~3�1Վ��s$��1���7�tkx}�R��~C�Orϑ?|�����q��B�eY��ê�mJ��fY٩�9�{��>��Ըk�sRċH�5�n�Ts�G�z5�'��MO����[;���mE#4��S�x��
�W`�{-Ӄk�ԓJ�� y���żwu�ʈ�wd�V�$q&�q�f�%t��l�+a�Y�*�$bC0�1w�ʢp����|+����|��l�I,�d��UX�U��!<a������囍�EbV�����#I��6��TO�Ģ�KX���-2�:	Q�A��e�q�O�E����6M�ߍ�{E���VO-0�Z%d���9�~w���Z5b�2`+��"von�'�BXӖ���������1F���S�}Y���>Ua�aX�'�ۓơ�&�)l�З+WY�0���*b�Y<��4�����/�|��w�W�}^o4}�I���Vߌ����U!¼�E�j�N�ϝn�U�U�� �R��\�@%���-��'��k�t�WE�5�S�z}^�.�����1�כ�nzgɞv��Q$��U�_˵>�Ͻy�Gǵ6p!,i�L�2��!����{�����|G�Pșh�$� u��5�����¾{(|E�b�����x��yL�v�T~J蜾�rG�:��A p�\l��j$�4;*v<��'���b���=�5�S�G�*�v"�80�[�&t������$�\��g���6�����o���{�א�"�����9n ȹc�Z�Bbߨ����ڍ�nI!%P
�]+��w;�5P����Uڴ�p*U �{l��n��K�Bڡ���1�5�"�������2�Zݪ��s&8���T+u]�5I���aP�HG�Tq�o]��w�  ۸�6�*����m���3N�6�� �*���VS�l*��w   w �U[J�z=N�*������en��0ۗHD�q�g��I:6�ײ�ˣ���v�[6�e+�I��mFU��3�'�{�e�<���ց��y(o/������5��,��yY�օR�Y��6[E�[�H"K����F%��qC�]~��n/^����q���|e_o�%����K�H�Q9#hēQ �����뿽v!�z��fL�׹>O�N:������t�t������MFcm��.:�Q{j�k�N1D�}��Y�}�,@���No�Y�f�p������2��[F� �5���t��Ԇ��J��N0x�H� �z!慗BedC(�K�vEM¢���w:�ӷwev$���S��z�v̓OT*���k.ͦ��4KI��ϗ�_/�}S�i�X�!U���3ƞ#6o�h_�ؾz��l�^�Y�ϙ�!9m�d��<j/�gt�g����汶լV�l�y�<)����/����z/Ǉ��e����w��[��3�
86дVM{��<�v�w��[>�ɢ��6Z�R1S�l�T|��l����`���>�$�:�`L'�*�*��L���ĞH����N��U��TN�Xfp�7͂s[>�ɻ�Fk��	<��}<�#^��ܛ�6V�w��~l�ģh��k�M�C$B}���~֤��לl�˚ϡ���KK剳�Q��UbGR���W)~Y�d�]M�o����D�U�;V�9�NzSOm�n�v��U[[  R��iȹխ�M���=g�u,^�f��p��$�F��MH�6N�tٰr�:��i }�)USd�H�{Yh�$�!�HT��I��	��'!{�vk]��O�	+������6[��G��v{��־H��>�ަx���cg�S�>�kIS0D�e��n'.�H�6O�z�߾;Hկ�6�&�9g���D�U�w��j�Q��.|%ߐx����f��D|N�H�����$������[Y^ˆ��o:?�{P���9<��8��L�BEݵ�O�V�x�۵��Q�ْIa��U_?��C���P�N������������1q��duC��g_$��&Й	��,��&�Y��Y�A�P(�UR�� �BX��K�L�18���#�TŎw�|�T�'��UA=tl��$	ďq�	�L+r�$y#s�S�~�E�d�Wܭ�%)#n*��[G�%W���͓Eu7~l���u]�H���Z��5�ߖ5�H_d���d�^�����m�#-�m�
FAn��h2M�Gﳺ�B�ĚG�%�P%��n�J�5��͟�?$	+���@�6M���$~���@�Rf6�$�?$	�V_��v�ϻ�3X���&�d�ޖ/�>���b]�֍�M�	/rF�x�L�G�休�@���L$n*حh.ɬ���l���X�W�O�T�֯c���	��,H����y#vو�tF�$$�A��}�<$�	-m�q���[�ql&�1��ʫwb����e*�w=�[m�9���}��N�Έ�(��la��o��)��5�;$��2����-U�Ҷ�ha��§c0�/��6�d#��m�6��;jCԏ�0��5t���I��ft8�\E�c<Y�x�AW�"b�t:!~O�
]������u/��l����qƩ>�̣M3���QQ'Տ�"=��i�iI�8�#:ð���m��I�,g�?�N�g�i�X��!��Sy�TYbaݯj�7�M�A�~�I"��;�+���6�P��l�*�������U���p�_���[6ޞ
�Na�d U�ehkK��׵m� UHrv��ڛF��Wp{����]�  \�g��@6�pUQT[;�m����M����   �@ m��*�P������~
��� �J�J0��9x�Vۖ�þi5�g}��-� l�(㶴((.U��V��Y󹑘p-�E��C�D��H��hSO�#���\�Hg1x���;I�H��GIZF�
8��o���/?����d��b�"�����CN]�?�*-\M$	�#$��!x���4G��s)�"�r�+�<d+�v+�K�4��5��*BQ�*�����J}�:́T|��.�?����"��;�M���~?�+0AU%��'8ng�j�X@GAɬ��vYb/�G��	7^����ӏ�<[�  ����X��ۋ��� Cd���]�5��w]�R�́�Z� d�+V���f)ٙ�&fඝ��3�����F0�}�DTī}����#�I��	��m�\���G��.��]�3�<p8�q3N?B8���Z?�Pв5�臲%�YG����k�0�@R��c��ۿ7��;�_��2��t�	�+?��YqUךA2Cm��\��.9?|{3`�"�	 YU��3�sX���Lg���ܝ��}���6 W}�0����]i�*�d��������a$ĉ$ݞj�Ү�ľH����T>�MR�UW/.��(^�C㶶�Zک��I�΅Pw9[՗��U�DU�:I�Q"x����Y�"IiM5��ef7�|����_��$Č\��m_kx�$���zۅ�c������1"x�M�'o�XݤI ����̪i�,��"O�'�T/A�ie��>�;����P��a�j|1w�w��WM��$�F��(�V��^H(y"���aG�<��!��_|�뗿<����S�iNI��<�P{���0܈�  _�":EP:�� �D���":4/$@$ S��A}ڽ�h�GG(�:���6"3�a���#p.-����5UI	�)�ϩ�or@$�ݾ����I��I�x�	)xĘڪ��K�x���C/%�'��?[7iu"x��1|�g�LKR7�ưĉ���~�wo���I(I�k�𸥐mEH���ߗ��N���:��u�����&$I �f�Z]�z�$�3E�OBN������2��r��m���Լ��m�7kъl�
� 6�6���`U��]WU/s'�����"W1Ԩ�Dd���a_]�K�<��>�G$�ԉ'��//����"~+�����$�P)-m[\����I;���ah-ʯ$I9^/(�1"�'��'�*�䉉rD�~��4L+5�H�]�I���m�!G.ΤI%�Oi���c~H�m()�R��*Sg��I�"I�6�[(��I�J{��Md1�KQI�$�걆���Y��$�"S��aie�w\���vn��$ףl�O��떹U�O�Q}�kEc[Dk�Д$�+����FLH�M�ನ�*�H�i��Iĉ���J�rD��Yțo���i@Z�
��F�-��iW��6����»k ,�m�	���� ��4y"YY�<H讼�:�$�<�_Bk��1"I�PSd�H�*SgA��D�	$����~+l$JX�j�w�;Sz�$�$�I>H��sV$I8�$��,-"l�K�^�'��_:�RE�{���r�+2Z*(Ј�f���uJϾ����H�V.��Q�I��$ޟ�D�V�$I1�[O�"N$N��/yDM�ی�ػ�FM.���_����4W��'�LH�M$b/%��ĵ"O.��=y���0�H�^���#��d[��h6۷������ҭ��I�J'�>H��q��T�$��%�V�'
�#�B��.�%Vڤ�Bc4�M����@^�uP��{l� [j� ��Ce8�i���lT����wzd��e>�T
��-)��}8a]dwm:VT̠�qUa����]�Uu�l��e TU�2�
�d���U���`�U�UU l� *��� @� �J��Tm�l���l/T*��-�r�f�YV�^�s����7P�M�(�d0[��G�_�o�|z�k���x�D�$|��]kR��I>���q��"h$�	�r؁"!5��;�읇�$��n�m��AkF�%l�98�>*��U�DR<�&tz�H�+�rG�/r�1"bGR4��f-ik�,�M9�e��[j�d�߂p!%9���F�&�fw;�A��#�@�KH�D����M��HΪ'7��B��6�Q����I:�z�	� �1"bG�7&�3g�sY%��?�̭s�Qsij��%&6�nFa�:�!v��(3��=ľ3K0�Ԭ��<X�v�C:D��wT�Y�n�j�r�pA�l�+��-7e�T��m� lԲ������%mUN���GC���?�Nw^����:�#��cNئ���j4�n6�M֛#�w�W�R�n"P�K8W�<D��!��ǚߍ����/~G����	)?aEq�~�a�p[Ұ�&�Gq=�M0�����y�'�C$qiP�U{τ�^Y�G+�х+�Rx�R�u]Y;^G����~���#$��Cy����gYs�B0ȴ��r�g��`��a�����~��	�"�ў&��&���&�:�u��u[B��uU�L��PjD�jT*����S��u��2.-�
X�-CL�d6am��^�4F���`�
r%$e&�"�;o��<B�w^8��:,��l�j�Bs���u�p�u�6���QȔm8�u���ZJçH����gN�x�p�eb�V_ ��M= �a�������v�Z�UW%*����k6�X��qdo�ؾ��8�x��0.�ME��Bw�.���,�k��2"Qƙ�F�&�U�����_�sg�{�|tÄ�A�י�k��7Og�"�l��x���E��
ⶡ,��m���v�J��Un�d�*��뻕�f4\I��d�%~gI�;����Qh?�����0��}k*�~fϨ��5���r�~�0�K� ��
�?~5=93��W�*"EX��kM�:}�o���K�Q�d�޷��ѿ)C#��K%'3e�����������咳�2�]�J����>8~8B�>��|֝#�cPТXX�Q3$jHd�6FuK����w:�$��H��	j��Ѫ�adʮ�T���������P�eZ(
k�5��ƴ�6a�<��E��R�A��;��}��VC�q���7���FF$�VA�V0��K�����@�*�)9ݭ�R��[�G�-w=�	��_֏�uc����-d�p��O�ϫeo��;Wڙ���nBNp�X�%)!!pmB��_t���95�s���}'�y�^���f#��ڳ�����3�[�~<Fb����!3� ������r��)�6����\kAy0Cf"��+;���j,[�;���K乂	~25"nGH��E��jݶxi��b�XZ�>�f�#9`�1+��:}fcX��w����R��mtiFܒ3� 反8B�﫮��q����l�K�yh��g�:s����:�#�����{xҷ�%D����n���lf��*TVz�ûq{p2����� v��� m��dw묞ղy����3� �b�v��y�0��b�|m���e.�^R��X�Խ�f��~�� l��l  ���l��;���T���wR̠
�b�p  p �PT��S�6��� <�qW*ђ�Ur����bwL��Kk8��O@m\K��HL���m�.�X�r"�mE�{��������C�*16���\hhy3�0�&�p~��u��)�E�&FӆI$l�idw/b}׎�:h�ҕ���L��Z}X͖Fr����g�:m�W�)�$17#p�%i��àˡƎE�)%z��>�v��>?oh��u=���<�
?�f6܉���s�Uxvcλ��oa݇4�=�2�bSv�����&�-H��ҥr��7?�H���^�-�7՟��g�,'c�n&Z->���N��|oz��Y��UUU��Wq��Y0�ݳ�vVU�oq��T ��uFۉ@��I# k��4tNUθ�q�0.��gRJ��?��2fx��[���ۖ��T��*����x����s�c�H ���a<}�s�{�Y߾��~_����C����I��l�Z��=����~}\կ��U�G�su����ex�L�J ��h-bJ�_���S\��[Ư�B����U�ѫ��,&���H��='&���յ�f�s��^ݗ+~�{��5����UUddIYP�0	vlmL����������W��:#�dUj2���.N}���߾{y+^,{6��e��9��4�J9B�n�=���=�O"���z3E��m<gQ�-�L�IiH=O4����d�k��m}2f��0]xo_�V�LL��I8�NI&�UR�;��OQ��7Z݇v7�J�ĳe��m��˯��m��V�9�K���Y8sw���>ٕ������봵�ˎI#iU)9(��4ə��_��W��� ��  e���iض&Zxg��g��}{��_٦��*�r��3���޺�\�\N��H?~I�ܐ8c�6U,�쒸��GY�_�Y���v��ȟϻ���JZ��}4	.@B15���u����]��J�G�cت,e~��:��j�?����Hم9�3$l"گ��c�{އ����ŵ��s\i�q�?�N��v�I��\�ϧ&z�� ���J���C�%-���|�n��������
�mg�b����Շ�?�����"Sm�j��<l�˽�������g%׆�YͶU�]���-5U\�/����{�X^NVC�E����}���_--�
�idZDO�G�5#���~���q�"JF�H�a5����Q�������P��>8~?��}[w���j~�t�kyy�A�i���d�K��3����uN\WRھ0���Gk!��Rj�#qw�]��O��+*�Q0Y������z:�����S�\?�J��&w^��ㇼR�>4�O��˗D*D�[��?���p����x��7��=+���:%m{}�s��'�x��rn9�n}d��g�Ɍ��⪫m�؊�́n�@  p�*��.cm� �[� � M�T*N�U��l U����l�ٵ�d��̎��*f�$ݸ�  ���l���  r]��*��6@U T�� �PP�[�{w;l� �@[ j�P 
�S2         P�@  @UfU�Z�EP�6�q��of�  
�v����PUU��b�t����Ic�b�[hw f[�i;5�4��Zy���[m�s
���[%PU��Q�b{�R���*v�J֢��P  �6�VBn��xؖ�:+�-s��Zc�y���f^H��*�&�D����Vա�����1��wM~��j�C���Tq��P��Wt;UJ�v�:�4<�6z�J�4�q��e�`1�2q8ʗn ��C杉�pqW\���^ѻ6� va���Ѹ��i	r��*���[h�\)��=l���P  ]z��u� P           +�Cn£lAT�  ����� m�  U *�Vڠ���� �M��@ �[%V�P�
�1y��R����w�  
�        �
��P    �    �   *P *��[hT��eU   r�@�� UP+( `   �    `U  ��@    P         ` � � s  [+d�m�m�  �r� ��� 5R�Y �Ʃ[-,,�@    mִ]��^@5�*�   VPw.x��`
�� *��[j������lY@@��;5B�  T���y���t��ƶ��-�P��V�N���V�c��׉%j���Pv���)<:\ٴ�Gv�Qʊ���lq�UUUU*�65���&�M��/T���UT�Pm��
�[rP�PUmT �U)q]�6m�� � ���7p
��Sh�l�t���cv����j�VH�Z1��ImQŬZ��5���ng&�k�{~������?E���5nx�GƎo�d���Ǝ3�D�2%�#���*;y0O,,���F���^�\V��w�y�u�����󰤔�s+qUV&�֟�[ΰ�0��&���F�W�}��3���Ĩ��˫�M�R�D�Q��Q�+1x�#��3|Nl��ثʨ�ן����O��+�|x���Wg�D��W$%���I	m�JH���gf�
��6��l��!��reV6����OA�/�L�~�}���A�[j����`��Ԯz�����!��V��w`�f�V �%�`��W4���������L{E��Gy��4Q��ޡgO�]ҳ_�n��#H���E��DNt�'�ԗ�ӗVi� !�O�i+sv[���z�{�����y2قB܉7�6�w꥛����h��_�Y妠/&l����U����Ԍ�ԕ��*�a��?��33ҕ�w:�9���:�ŧ���0�Jx�&L?���]��C �KP)Fk�T���u�߰C�ECRZ�l�ϕ�L���^M~�ϧ&>��V�em�m���nUq��yU�=y��d�NM���<T �+��d�,����u���雚�n�����w��d6D8}Rr��k��HV��~<O���\��7+ib�čK���Y���R�ѯ3v��8_��c�Yg� |{�צ�}��ki_�I$��F�O�Q���ky}������'��d�+L?��'v��_�����m��A�6�h�a)�$�D�~_d���Ӛ����I��@��&�-q��JԈ%Aq(Hd�+�:D=���Y�D�r�O�׊sv�6g�ʙ��n�{'�/�j���j��U�(�.w𪋉���ʰ6�T�s���ʷ��܉H�Q�Jr���Z�A����f)�E��� �A:=�ekP�#�L�S	>i�1��Z�OWP?��H_�%���:U�o��o����D|�F���j�_Ə�j��~�����J8��!��ʆ����6u�#���Zb�
ڶ0k��G�ל>��4�&3��%^&\@��=�d,^h�(�.}�rf�g~�׬������W���۰7��xKזx�q݌�1a�kM��D�*�D��ܒI"!����B�{5mD����s���w
�Scd�[[(N9��R�S\����d���FZqiZKϰ|l�#�'�X~����f��;��Fj�]���-���%��]��� ��,���ъvC���N���t�iɠ��ޭ=��,��`�J�W_��3�����ӓ���X_ ھ_a?o�������Sk�(_��m��Fr@�R��5U�S9�o	\@���s腙��şo�!ZF�OL��g�P���[%(��2T�k\������z�ղNf�Z0d�~��e�#w��\�
�\* �׵fc6l�*�s�w
�����l��@  �m@힚��	�V�����ܯwe 6it �svUDyW\v�nZ��ѵN �&����`�CbJ�k3or� c�l�T� 6*檪m����`� ��  U-�   ;�  6� w ]�*�6�k�ٰVU�c��TP yV�p֍�h��������[�r���N�����UmK����؀�wMuja��^�+���L�OnFLɍ�L0�31H�M�QO�]gVs��m���f�Zw{ʁ����J���-�$fI$'o*<D=D�p"<n׺��q��aYc��^:FQ�{��j�5)�!B�$�Y�ќ��5'߳�^���P�{o?aD~R�I�{(���˽xί�-�v�d�K���y;s�|��7�ݿ�>۬wW[���ELF�L��j��E�;�ݭs�ۼ�UR�ۨ���� ��v�Bޝ��L�*@�ff���ٴ�}�f��n昢�J����0I�J�I��oI��J���	|!`�	1�}�w�L�=6q�N�z�]w���v�"�h�ւ�]�ڌ���=�[�/U
��3��S�;���TX���y���O�����M�{�u(s�ᜰ�e�����e�SH�q�d	�$��Yj�r��Ȍ���~8a���'�P�a�>j�i�[�}�^��鹏�_+B���Fj�F��x��ci݃,5�w-��
�pU*f+��Cv�TF]�����ߛ�Dܶ~��HE�'�̄C��1^֖[Cf.션F�ϲ$*(�}d���Z�V�Cӻ�i-ʠs�W�t�������Ð���E�a��~4��mE9#�?�"s�����Ǎ�/~ύ����/ˬ�)�a����Cu3��<�.c�UG*��S���v~R�3���y���=�NY/l��2�׵��jN�L�����h�E�ش����R�x��rE����0�`��'�L��Y���[�r�Vj���|������ym�^�� ]J����UUU*�\��5�]��U�h����_-+��.�"4s~>0g+:l��-���4x��P��4٬��Oɩ!��p8����c�45����,}VGG3�#1U	ʝ�C��Um#����2I#.J��"����F�v���6���I"�"�2��vzjzs���~�v�I#lJ�(4�q��8ʿC���L6F��Ϗ���l�����_/�K�g�K���E�rI�k4i����6��j���s%���߷�W-	��k����S�xcR���6�R�U�$ wP �l�h��4*�kK#!~>���#w�������k�=\�fA���DIE��qħ��N���߭��M��fY�WS.��i�3n��nڌ�AR$�qFdIɵ2�d��K���s�
�ɕϜ���,�@�_��I$�#^��w�Y�_r|��vK��-�w��ru�k�g_6�HV2�*�Ūv��}��o��m6�/�	���<wU�̔����(`�w.쪣b����*��W+Y%�tQT   6�x���s@�;�u淑\7;���*��V�:A���藤��Y
�����K���%j�s�l��KGb�UUU��*���AUTm��Ue*��p`�T���[%ͮ��P�  Wu qT)m�?l޹�
�����;��TpT4pMT��OB�Q; e�yf� wu�*� -t��M�Sr6⢍�G�5d�ӎ�X>���8Uw�o�^ٮ�e�VEUR�vgfa^���A��l���B�<E��`�a"o��Q+��v����0�q��q&T��#Z���*�*�x�8æ����c4Y��lĴ̇�qx䵈��=A��d���Ǝ����q�j�0�^im\0�3�`-��=��Q�T�������B�P�%�6Y��jc?F�D�kHmq�%��g�}�ՇM�'wz6�m��i�ڧ��q��d�x7\�7=R��ky��w@m�+��i�U�
���vnvnn;���D3eI"�EA���6|p��֮��#"�Q�M��MD�nF��X]���n�uq<�ƬD\� c��Ə�0�g�)��\�|a9F(��#�|�"�Q�q�B5�3�wO�V��Ζl���~�Bϥ�.��l�j>��:��}93�����A��K�0�#�N}��w5]�-�;O?h9Z+fV�-��)��n�m'̿�h�T񼒆�]����k>�w�7�����5I�^�ͼ�[�lm���&�f�,�[�
� ����d�FQn�m��&���D8��8�"�2/Ô��"��S��B!}D����Bj��ĩ��)ܒF�$�Y�Cǈ��}�E�qM�~0�7S�:^C,���5���ّ����%m�H�D�v0C��"���~0�5���+�r���~ZۧV����~���,{���vN�%����01�$	�d��q��Wcg�8�A�rWI#Xdɣ<Et����kH���ڶ�ˀ������k���$��᳚4�"E��q/�us��n揺��h�Vѭ�"���j�'������뙕�՘��W`��ʪ��e��J�iE�-��+��s��*�T�UJ�6����Ȭ��9�����E�&�Z5�~ͤ�/�&�k(fF�U�ee<i#�d�rI$%�US�J�nˌ�h>�������nK��r��	kj�ѯ:��r�((L^����v�z�׻.��I Y%�E�6�,I<��ݚ��{'����?l���f�j�
��沉"�."�nF�Mm����U<�|+n\d��;圚ޞ_�|�
�#��Un�Ë��`��Zӽ��o7v� TY�U�h%��m�l�ʽ�w;�߯)&��L�7��W�v��c�뾆F�n8�e����[s33^I���/=����CL��(�*$��������w������D�׷D����b$�R4��ƽO�+3EX�����>d��������y�����[
"@Hi�$��&�w�]�w��ɷ�G���k��lK��z��$F��$�� �Un�q�3�VZ@^�W�T�Bv��]��TUT�a���XuA��uԫTW]��*�=8���f��}cI�6�a	U[U<��7�A��wO)s絜4��/]����j� V�[[@w)�U&��{���;��m��
�Lȋ�*��   �U xJ��UUm����JZ� ^�*�2��^����l��α�)�;�� T��\#����P�F�r��x����3۷z�4��S�Q��\x�+�7�s~h�J�I#$�|al��ϖ26әB�����x�>[_c�4�-������ձIWͷ%DbnFۍ	N��t����꨾8G}��?p�S��y��!Ҝ�,��� ����4��B���r
y���D/��U�%C���%���UʦJ�dYgif��(ޯREW%� �"�'j3QW8~7��࠱�t�xު�b���`�<B-���di6��P~�XԪ�J\4N�{\Td��Y�WiW\U
�� ��)�[�]{{�,Ȓm����#u\[V
�YW�v�wZ�mp�����.X��T� R�0�%��K[���N�������m�1�W�6����7����mv���Ffk`���"Q�#1siǧV�>�yd����8r,�i��3.�;9;>����IWUc(�O�f���#�Ls�=��%�(���<��'���^�a��g�&	&Y����Ě�IB��F���"�z T.���p�nmV>A��V�ZL�x�?~;�������* CkmnU�:���Ӎ�<r&��Q� F�Uj�VP�m��c��m��I��+����|p���!�_�����g,�|´~���E�����6O%�bF�k�Q]t��'���VYr��3G�]�p��6a�3'�[[�C�c��UM\��NH$�����C1O��P�8�^�垈n��;
��!�r$����>Oߵ�~b�1�-E�����_e	~��i������O�*Ëq"�?.W�����"�i3��"?W�ߎk5W,i��3����	��]������ݩ�\�NUVL�J��I	[�wk`�ʳ���L��lN3JN�/e�j�j*�l�����o։&�)��K޻y�۽�O����i�y�������
�������m�ˑ��M��q��Vx������ԇR�O��d!b�x�kq"�;d0�,�K�|�fQ��mm�FA�Yf=Z|�[?!خ+5	������G�o�?WbE����.�x��usIXm�I$�ԕ�3�wN�_vs��������4}�U"�`�m_���ڽ�.��Z[�%�(aƜ	$�0G,�hL���܇�!��R��_5�d##��5c��CQC��*�����z��6F�e�/a�9on��+��q�j�v�cq�9U#Ht7H�C9f�V(�=X��:��%;/����r���B8��7j�-�����i3��vB)().Vyn!�y���#�fԛ]p��è�Pl��h���M���`����\��V�Vj�w�v�]k��O
H�H�ե���~�8������d�	��+������p�=SE|.��w���@@�kG5׾9=3�rws۔$]���}ןg����X[����&_����i쎘�HڍĔ�ql���wz�[��U
����m��<)�T��  �������v���m� mKK��gZ�8W�+K{&��F�n�E<��`#s��N{%��3�3���駝��oF@ 
� *�� ����2�Gp`� 
�P ��@ ��p@ m� ��[[*U���^ر� 8�&�]͞�����VVU�vϴ��d���2�srە�1��T��C@�$%Y-%�_�������;==��i� ��z����'��|r��%��hw[�]�<�%�8Tm��8����:F��*�t���P��7�g:�=��3dC��������S��SI��9�(� ��ȻCs�T����藳b@��Ȕ��E�>�ΰ����#�c��K���q��&䯍ş'�����[%a�8��{��47L\k��!�7
ە^��s�=�r��k0�֌�Nh�������jǢ�L��-��3x���
�M����Z�%"F8���+WQ�����(p�l=f�s�ݤ�{Y��UU;�����V���7��*8���!�����C=Y��L#��/f�[�dJu�R?�ݨ�J���̒Hˑ��WKN�3%s��埒���wW���L��HgK��g����j�`�0��zN�Thط*El�Ժ���X����g�+��u�!�C0�����2�ٸ�Z�yd������ی��U�.��>�*Lq��x�
��~�3��T�����w^��z3�9�}�Z!%�@8�h������wNt7�Äof\�#��X�ZX��>2��{���-�����
ecS���)Ψ��ܶc�v���2���R��I���U�UR	��ؐ"�E��re\�.���[�k���TY�1������6�}T��"�E��RD\��7�/���
i�i��eV�rR¸r˔4�B��X����l^�_��:M$�5w�nPqv-p同0��I�X[���{םQ�.��;�6F�3n��a�� m��rr���S����F�7xP�����n���G�d%X�A�{)��!a��߉hLb�6��r6��ޏ'&�a�C|�`p+�ȇO��������>��:��4�޶�iF�E��8�|�Q���;���U��ڥ�U ��j�����ej�EUc%k�뻗��)��g�t�nؘ$[�'��4�ϼg�y����R�+jzng��Y�꘸퇐b0ن��uVO#��Y	Ȼ!�;BE��g%J��[i&�m�J�,��˾?ap���|p�%�|~9����F���eV�{��sw�5<�=-�ۄ�A#��������תg���8ا�!�Ru�C�s�S=W��u��:�*\��(A�(�2I���y>���}��~�?��_b�Zf|0F��G�l�ʻbZdϓ���eBZ��⪪ⶦ6�slq��Nym�꫻�6�M��N�dX�+��KQ��kӼ��'�=�lz��,=���+�C���'�/��'���'�kM��F��\i�S�)$��#��.�R¸r˔:g���|����G�d;�H���B|Y��C8Ȉ5V�!q�{��z},����ܼq�x�z�G\~��㧙��V���?S�6�W�<o�{�����m�#l����4==3�;��4ݡ��.�/u�#L:|$�8�<FQ��d0�΋���S10�[m����8k�".���=�ST�>�t�܅F��O.0�6)�{jb�Ҏ�:��ؿׁ^;��;n#^۪!_�O���� m�
�X�6��UN� VR�  �U ��*UUJ�JT�i[fŲm���*��K[*��f�Ug�YUUg�4� j�� PuJ���   ��T� ��V�Y-�T6�m�@AT.���  
l*� �Y@
� m�      UT @ 
�  ꪶ��,eP��]61�ooK��    ��W��~ݺ  �{���z{n�{.�1�� ��� UwSv�7E����5P�	{F�a�Uf� U*��Ų�c`��:X:P�� �fZ�2UU�EP�
�l�e���横 �z�r+�g��S�����Ņqf6!8:��5v����;sv.���$�qZ!�%�'.we
�����%[X��J�Rō�;�&�2�b����H�6R�^[r��V��^݉����C4��
�6�b�u�b��U�[ne9k�[)e�<�8�h�w[��/6 �&��Q��6��֔�� UwP
]�(ٻ�{]��@         R�bٵ�l� l�����-(T  �  U   *�T[���P �۬�l�ͪVPUM�U��m�WEY[6ι�   �     *�  � �P    l    <    �l��U 
���� 	�0P
�   ���m� P�0   �    �
�  ��    U*�      *� 
� � �   ��-������`ت]�  ��@ا{����6�@    �M@��+u�@ � 
�
�UPt�n�;�J�  Sj��b��Uݔ*�uiz�˪����R�J�ڂr9����,[��L���Oe�Ca�*�۳"�e��iS���e���ٳ��o.;��wf[��]�M��t  �⪩TYwM���T[j��6�� eUPUdr� ��  � ;���J��P�o^���n�uhB�r���Z�'Z�`��5ͻu�ٻ!^���©X jT	\��&E��04�"Ϗ����(w+��=ٞ���{ʧl������',�J�b�7�mm��F�+��Fzk��}�؝g���e*�|��6-唸u��\|xæĜU��.Շ� ��SH�n���Y&1_?^]`��N0�6s��׆!��^*���0��ڛ�.0�My7m�JrR�V�qk�Fg���>�*^����L�/�qC�&�m�4x��}��J�dq��o��[k�$۪I#WY�R.;a�!�8��Y"�^#ضD��8G��)�Ex��4å�~�W�% ���%��ٲfxWв�ѧ�� �ګ��f��]�M��ݔ��E���2��-�a�.p�����TC1H�U-/j�I����=��"B����9[�ǈ���q��˽�T%�B�2�Z��ڶD0���"�P��/޿l+��s���>[�cd��(6�zng��Y
9�EǬ<�6a�.I�$Xa��%��8C=��Q'��*�����	%qzt�g����t<j�!P.fGf(���zM+2�T��@��G6�B��_m��}�]R�)��l1l{�a�.I������#����^�C�[e۵*�ε���w�U����
� ۻ6��s��`������tzf���Q�OL��՞��fE�,<�(<x䓗���؏KD?	
1��p���4F��Ѵ=/!g����'VskH�&Al����[\z�Gƺ^��h$���e*���2.*B�k:Y�9/�C+6��lS�٣㜴A�_��
w-R0�d�̒H�qК�-���ݜ�c8aT9(�0�tʊua�Y�h9c��k�=7=;0v��!���(-��V�OV�CŰgU[6D�|��/!v$]9`�n�x������\��X��:��x��v�l������\�]��� 
�U���j�
�t�6�ذ�%*c�n��o�iv'�1o�v�Y[Z&�x�V��ؐ�CR6�ҢEX��J�%7���Eg�����.t=�v�s�ޛ�� �'�6bH�C�-��ʦ�c�tꇫ;�o���m�&�Vv]��I4vH&H�i!.mg��r��⟂���������ey��Z;�4��w^�o��a$���/Ն�?U^qږ�eouY�+>�=���m��[p��U#����D,�n��]�m�emS� �	�k�b�3�-��ݷ��=�ԝ~�*��Tɇ��y�x9�~a�w
���F6�Hn��7��΋�-|n!����`����{T��߫!���*���0�H��m�vm�d&I#2#����������ãj�O&x�L��8��0���[�p����}����U�� ������}��E�k8����������s�V}���`i�������ًQ�4�dȋq�����t�����v������#9{A�d?���Œ�������w�=���������-m���@�	,�+
�,�2�+Lf���p �  *���
� vR3lk��gH:��VVU��둝>(Mԅ�i�.nD%k`�-�v���[������jۜ�� ՕB���w[�\�*T�n����;�@U*T ' m�T;�������� �U�� Um��P �p Rɕu���j�#`��	�f�fGi�Et5K��j����U��`\j<��1[b¾�MϦ�e��y���ԡ�^3���J�}��ɞ"<�U�Y�;?��mÖ�&�K�t���L���g�8}E�Y���:�.��0CfMp�{����G����RB8Ĵkm�&�3��=i����p���+9h�_�Y��k�v���&��M��JI MH�ڿk�Y��|9wP�;�T;U�L�:lv��wW�~,J�������o� �����+V�����������R��!��QsVs_�'j�J��Ǝ����{$iH�	��p���Nݲ9��ۧ[�@;�m� 'R�j��"Bedq�U�kϼ���W	f��_������t��5����ໆ�9��U�ۍ3��\I8�& S������\�1]z�	2�7%��
����;�� ��ZB��ݽ>�>9� �ċ1�܆�U���#��ۯѪ��p�\h�/ǟ;����G�޵W���5�ܻ�6�0�FF�F%�Gw۪�D3;6�?���x�������~����o_�X{2I/�fF�I�6}�����O��y@������x�"�����כ;?���m�(���]�xڌ�zR�n��� �PVڥZ��hA�b���F��V��i��Mg~���#s�ۯѬ!yåi��_��wq���/zz̙K�km��s\���j6L���C$�����l�k�E�ix{�ϝna��S�C����EV��8]~�a��w	���~SJ�R����s�
�x��&�j�q�p���=H�Gţ#EH�n[���Mں837���W�w�2M��bdat�y��7;�>��9�b`��m�X6\��=k����44ז��M�g9s�밪?��x�&��19|�o�nJ*j��R��p�ʃ���W�/T��t���@����um�ױ�͊�0����� ��C�R���
�K��l������J�Y�ڮ&vb�p��UU1!]g���e���{�C��	:��BEz�=��#~m+�l�����yI��5���[��<��T��+��0�2j�hnԼ��퉽�M�s��']{c\z�{:��¶��a�7hwz�w�p���3��0u°H�ί���_���������S�'��ѯs�XE��,�n��7�����'�>8~;�M�y}y���M�d7J�r����s�qߖ��*�BT�b��k<��v�/_�vJ���B��n� �)e@] u����́���R��������4sP����W�h�2j���x����n�pþB^�AK$��F�U{�s��{'���e
����=ן����4�+��8]i�S���뼑��(�#n\�ע���Bken�7��PE��E�BA|�yq�e��]�����)/�ځ��2����L����Qګ�Dv�kt7U҇��ï���Nmz�!�E�89�v����S8���e��a���5�2I�Y=���Zza�9����,z��.�S�f�r��[�]�U]�e+\ t�w9��uFڨ++ki8T�׻j�Ve  U �ݭ��̣�{�.X�S����*����ob����z�3��e��p3a�۶���+��lZ�]��[36;{`  +��@*�@ �\��sTk�Gp;�ݶT�P++�xY@[ 6�� ���� �*Un��n�pک�7x�6���MT���댘{j{P��*����wjw *��
��cy� �UB����m�����!�!���Vz!��/^��s�t��c��g4P���d��jn���)f�}�;�>��g�<3���w��m�OV��Hpq�6ې�\�:�K�2pײ���[���h=5�H��=א�0�c%b4��6h��r2�RCy].���Dx{8O;�^-�^�Yq#�O���nP�Y�|��]ip��v��&\iLnH��']��?�<��,A�ٙz��-~gu�>N��]-8G>�βz��.���F�m�:�U�m�y���n���n <���.j ���V�ng�t�ڮ��҈��dՎ!��.;A���7�K�%��"��g/�b��f�$�C"Q��r~-�\q��r�j�jb�bX�a�Dr]5f�4��B�]�
��}n%Qd�-q�z*(��e�P��b'%6x��>7�o�#�]���FEִX�-����I�Y����ٞ��'�WWUȸ��ٍo�oغE%�:D:]9c�n�1q�/ ��Om��K6%�>�e���	��q��p6��C�z�u,��p量;FkC����[1/D3�P;|�_#��V��D��b�F5�2�[mx�6n�cg���S` ���V�m����J�f����7�x�^���{��6U�P�g��w2�ɋ�l:6�Z��%fˢQ.L�&�N9�t���C\h�!ڪE��M�t��z�����L�����������v�cJ�UhT�xji����U�W�����y�\��׬�m^*:&�ǔ�8�ˎf뀚Ռ|�N���)���oT����84n@0�P��:]�9K�5�g��,��G+��%���I,�r��S;̺�Y�	^��"���bm�gK9�T;//���������>6��$��)?I$d��u�Y��2��P���cᒴ��'�*�!X�9ʜ�m���ԝ�����݂e&0�Cۧ!��9���F5#�;%� JήZ�6{ww=��)*J�*��,�
ۋ,,����p���{�x��ΗB)�7I�#4�q�n6�f1\l�*���f��L�x��Xȣ)qL4&�t��s�[�|x�7Q%h$=#��h��gHeb�`ڶM(i�$��o��g�z��p��2Eո��!�2%�5Q&8�m��)8��h������<ag�&�|��:���p�4������u�����=C����⪭+��8!V��2��,�J�>�VC�3�dĪ,�]-,9�o��<Bsz�)˖z z��wcw�+��������+�,��P%��������^�"�>��6~;�Ԯ����>0�Ϧ�ag�ʇH�����di6��ɑak�UTZ�����OY�zk�V*kL��ه�!V�adu�7����S��;f@�ihV�."��Y��E8��L��f�X>�W���ɉW�9��R���U�d��I� ����n��w��iE.d8ΐ�Ұ�El�Y~A��u�]{����"��-EKqz��n����c����#&�x#��u�=��_���VV[Ti
Uy�峸-��P�R
�����m�R�UP �ٞ{ ;�U�i*�vi���̸� V��j�wvX��wT��Z�y��U�s�cYɻ�K����~Z�  9��P  �۲�*e���6�� eUP .�P� � w   o�}���� Wu;��(b�ۻݎ��Vm�˩U��p�Np�>�v�m7p�Wwu KR���u� %K�"@H���	�s&_�նp���g��x�T{���di�[-���؎BܺUd���F����,�	�U|��r��gHeb�pJ�4.(|F��.��R[b��U�z	�ɝ��y�f�#L�u\8C8z�ز���X{w/M��L��?ͱɁR�D�5ܔ���]�1�U�g}�������"�px�g��v3���RV�W$��\���4��i*��GO����0C��0ˇ������7Y��gO��	A�� X/Rh�\�i�[[����TƝ�� 6��kR�k���ۍ�]�gO���_��G�Ϭ}yt�����=mOVF>w� H�F �ɕsY���L{�Ծޝ�f�Er��s8E�h�O1Y����digJ��4���"�ʪ���I�����
�gH�9�+L#O����VB0bg�0\���g�M���Q݉Zlȑ(�+M��r�p�?�K0��&����x��D�gK6���X���l��m6W�q�2I%�t��!Y�(=�6\ZFK�٢ȿ-I�0���}+H���p�I�Q��G���g	S��w[�փe��[(m�&�e����~空ޛ�6TQ�U��5agH��[0�0˕����2VJ̈if���y�,���~�#A��e�MN����~��܃<pS1\#�!�x!��n�K�&��gz��&%(�Iq&\M�!�>v�^Cg:e�`�ϝ��+2+��i�ҹ����2kH��0��8�1�ZE�~��G<9v�a�Ds�-5"ʶS����/k%l��:,�ClIm�-k�W��s�^<v}Y���K^n_N����UM���-IMUz�`�F%��\�$���rm���r@�*��;;*
�q��v�L��V�^Q�9�N�MC+F��f��oפ��mZH�ѭ��u���۹�u炲��t�ڄ����aU�N_k4x���4�a���6�$�qt��"�Y�ώ��*�pߗ�	��t���C���NL�u��ed�#V�j����'	/J0�>mu\8Y�\同,��L�1�e�,��&�Y7tnI$17igHôaxh�>��ZE�7�r�z�7�f�4�z6�Dbp�7w���������ۉ(�5�J��O��UK 
��YV��u�ڃͥw{�a��BV}Y��x�z&�t�:���oV�di���<E>���i!m�0�WgO���C�:x��J�p�4��UÄ3����6!���C����?�F�(Y.�g�>8E����,��zp�8x��[�8�Ӧ�1˼hq�M��"�q��f1��g3���)���d�������C��>!f�[Zl�fm6�AzF�QƋ�D�i�4ь��4�:|o�w^t�\��%^4dͪ�l�j&�Ͽ������� �P�Pr�mΑ5�RE�++̫u�W�2�;���U  *�gwvZ��z��ۘ����[[[�*�[���3����ϭ�]j��4��N
�p�c�lv5]��]�;[PZ� �h���r  S�cmR��U�L���U �[�[T7��T
��EPj�*�l
����<UUUR����Z�F��o��q*��T=K�'������n�!ҫ�����V��X ��/'l�F�I��"�y���0�FMޕ�G_���Xp�:xc{y�,�fZD��.ZȪ�*³Y�g�S����Sn�NVq�<x�!+$���S/׵�q���.i8܍��0��gD�0MA�2Z;VȞL�W&^l���߯H�<^�x�d�Kr�rD�u�{�s��20�fP{	�[��i�H�-�G �0���Z�!��m��I1���:A���ȉ�Dk�H�!O
͕���+�U��B��:�ލ�릭�P~w:�z����v��hU�U��r �[�n���ԫ�;�H�i##��Ȳ;u[�h����c�oiz�T�:h��5վi��%"M�"1F�H�!��nq��ß�IU�Uc�=FI��,ٔ$�"ȭ����v��;��J3#J0ےa�D3�¼��#:}B)�6Y�=XŲ0�X�3]�Ha�}<�6�&Ir$l�Y�6��ζTu����<m��l�da�k�:G��1�"���om*A��JI!i�CA�����6s�O����d�af̠���p��yE���MU �iC5ن6���[ӣ����Q��UT�.�*�1	tm0�#m�������G�?k�ZFG��i��J>6D��gg����(���I.J��>�J٤2(�x��`�H�#kjŞ"Ί�{�� �7��r@�'m(�����E�>#*wL�x�ԫ�7�;;7���ϼ�|Fg;�x��	�I���Fw|�6����G�BٳS��0T��dag�˼j���}�e�lC#%��E�c!��0�v�3D3�=�Ue�"��^��6t���m�ψ�_��Q���>������ٽe�ܰ�ѹT.d;mI5TR�UUuzSs���]�����2�����o!�:m�*��ȳ�o'#��5:���BB���՚��Fe�',�g��l��0�#�7Ҵ�KK:�w�M�XJD�nFXJCC�:h��W	���@�v�c6t����U/!Y�l56�<��Lz���	Y������N�v���!�!�c�Y���M�a��ݠ�{D��w��&F�p�[�ęj���#���g7mkɸ�c����;�\����*F-,[����݌]*��T�h������ 6��JU�m����� �l���j��	>�͔2���{����^�L�J��k}ʸ���Y��W���s��;�7_b'�a��}Xΐ������,��y�'�;93�w!����U�D-צ�#L�U3g
�gV\Ap�`�:h��«M#N�D��8�q(�q�J͓G���Ya�W�cL����=��᝗S̓۴}�n[JG$iȔ�FIr=�m�%����b����YS+х��s��u����w�,U
:y��v}�����z���j�����*��U6�H�[Y 6��?��mTR� uUP
��UUU 5H݋��, �dUVeT�󪪋oYJ�� ���P�
�m��تx 
�
� �p� �0�ClUӐ
� U� �WV���  
��U
��� M��   U  �U    P� -����-��m���6�'r�w���P  ���;ې z�/YGWv�`
��� *�����qڼ]�5[*�.y��n�� 0���d⪃b�E�*ʨS���4�F�*�� R��U]˹�ܪ�٪�U%"ݰ��Lv7�UU��3NX�n�/+(F�N�$v������;TVt��bTŞ�;*��3Ӻ
��7s�VQ;�UT *��i������jس^)[tSrvױ��;m�e6�qɠ�q���b�wlXs�6�.>?:�C�^`^��:Π)����[o0�@�:���S���Wp6��ցl��~~]uޝ�P   �         -��Ԩ*l�E�{m@�@m�ت l�   �| ��T��  X�n�T ��U����U 6�Ku�m�۰    T T    ���Y�     ;�   
�    U�P *�� U���U   ��r� �U B���@   �    �U � ��   >�@         m� ;� ��   U*�nն�UU@  [� P�� �0w^���P^�@     �U@�*TW^�@ ��� U   ���ݻ��R�R�� ���]�M�ud�UGn�Ű�ik� U ��n�wJn^�YX���7@Uj��#J m�������=uU��M�ni�٬ ����8]�<gv�[X�-;*lR��홙�  Vڛ[ U ܶ����*����J� �� � `U
�6���UJ��dm�:�s�6Ͱ ��*�Cʦ�_yC���ӥν��
��Wu*�@++mU�m@�+m��5oNj���ߞ��w�֜�[3M$2�c�M��r����_x�|NϹ��4����L>b)�6|p�C&c0�4������I,HԈƔ(E �0�9ZJ�u�Q���jm��K<Cv6���Ýg���Y���=�QEn�lBRq������K��Ϗ~r�����F��#M�=�W�Y�iIs<	Z�Ɖ-��t�����������:|<�����=B)�6E�a��%Yx	�g��ШR�I�w�o9�7j�QW�=�\*� ]n��n7\ت�E��t�l;r�Q:y�J��E�Cѫ�P�g�΂�֑�Q{܍��Fd�1�Xl�4`zw�������@�ѓĊ#�w�,�!��!�s1l!�n�KY���̍��AU��a�3k#����W�����֖G��U��D/	�k�F�B[nF�
8�qT�Doq�4���A�sq*Ş"����/���<��DR�j�N7�E_�C+���a�0�T6���FewJQصz�eLǭ��t�UUPm�n0�@�ɯwv���OT��R��]��U�����I$�A(lCH9���j���C�B�_½�"p�%�<C��I*B�I��q.��C=��x�飇���/h��	O]{�߷��-؅�$�I�'%#�9[��C>gVma���2�����E�G�R�ib���b
�إ��}��9ϴ�s���Su����ͬ��<�z�x�eV��-�c%%V�0���XEe�vqY�Q�(�/��Mhx���A�m ��`w,�k�uA�u��\�5�q�Uu[ &�ZئK�s���q�Q�ku~a;9��>�j���#�Oy�����͈YDL�)�Z����k�����>���kjŜ<Ac�,ؿ2fetn��y+̅��jE?'�Z�u�3��*�y��߳g��9�s�hU�Tfiu���J�`�$��]����_�V.���}�7���;GfYi���ץs����ũ�ō�,��סl�Ҕ)+T�]U�F�%�@�ȉ�'�.͡��@̭����ˮ6�-��!�C�0�/A���l��4�C7���<|E��6�K��"26�d ���<:�٭0�#&��Jܽͣ��v�fAOޣ31[t[���i"K�:�n�����s���ۙ���9��X����M�BEj6ⅹ�Ywp�a�z��?{!/3���5�V6��Q�D��n4a)ŵ��h���6�����2<�ëԽ�[�-\m��nF���!J��Y(�f�a�T;�T�;� @  w9'iF�vD�J��S��\X�<G��� 8m�el�.��_lqLڞ���t<X籫�N��pt���ռ� S�dn��TU�qR�c�h�l� �*������  *�w   m� �+����*R��R�r����;��{����p)\��*�.+T��U�K��޸@�[iJ�t���hܑ���[�������N��������r�}nmS�:u�#�[d(޿?��{��L���[�lX�~g��A�I#���2H�!!��'&���L1�74�{nY�y	Y1Z��V�%W��$�qG��%6nU��կ��"Ϩ��`�A���2j�E�rR�-��Ϧ>w!�U�WU�i�L���ʑu\8C8}���P�,�'�l��3�u�<G�I��EI$�\f�%��Y۷�u��m����+��R��T�D˃�/k�--F{'ξ��.U�,Ç���`�q���A�gޗ�b�N��äC��G��*�$�Ir:�B�q�}�e��2�E;��0A-�2�ڵ�Y��Y�yw�!�BEƆ�5f�+<C���%d�QEF8�t;��8Ew/9Ər�|ת�X�0����D7S<rX���9�.��F�%�!�I#,:�Fr��]���W��6�Tz������v+<k�P�xUq�܇jr�ͷn�n#$m�B�:���Ī�]�].>>Д�^�:�>�muL�>\~#�����o����~כkd�UqUUy�.*�X���jv�Ԭ[wqd  we�L��[�q�+u����kҕ�o�Q����w+�z�"?_�������5���rR��
�F`N
��7����M#�P0�;�H�`�=W������ΐٝD�j	������r4&�
���d%d�����z�����{���=��nzI��7�?�[+�V%n�oPy{���y��JV<l�!�+sMՠ����Fo	�ivҺ�&�Uu�!�bA�!��kUɒv���߫B�u�%�S�m�ND$�UV�ř+m�0�pp�,����@�͊V��Ц�q�QuuT�[V���=���ɔ񬽭M��/ʴj�{��_��,�� ��T^���t�yRa��mM{}��^���5n��k���i�KmA$�@�ofA�V�ݛOX{NYg9�I��q��Yj$��W.M1��n"ā��(�{ٖ�Y-Ł�>:E��٢�p<{X͐�e��W<W�gsx�-��܊##uwhXUWx����Ҹ�9��'����!�j�M��Y���%+��L�~���TZV��T�Z�A��]�m�:8�l���T�,��T�� 
�GU�-m�mm�m����r_ߎW�D3�
��H�r��T3ՔaF�3��_<F�m.)H\a���"�7hi�b���E�
g�`�I�O��G56�_��]�B�p�"2K�Wf��$Tx�Ǡ�ٽ�5
�]2�Ҙ/���K:r��tC>9�s\���AU���;�]s�&{�J�p��in��!�	o�C9C�9﮽95=7�w��Ƣ�(�֔�U�"8�&�o)g�
��f+�롆��њ2���������uT�C��U6��]�3J�Qt*��plJ��m����*��̵fzA8�Us ��ʕܩ��"�[wb]ً[v���0J]�Ӗ�T���kt��󫻦:˱��dN���	�T�UU 6¥�aUT���u;��� m�U@ � �VR�w 
l� *��������7�m�u�� �P.�U�V�J����Om��$^����s�wU�\�@ ǲ��*���h��G��<x������P��3چt�܅F��C���/`݇�	�ބ��
F�%+e��Uק��93�����qq9:�hƆ�=W0�U�C����zc8�1��m��Ja�9Q�T!��pU�"/%�U�(��N�*�ܰ��*�RA7�b�##mFD

��r�/){�v������^H���d+�X!�^�vZ����g����jH�I$�.A\n��\v��VB,äL���x��u\8{���mc��f6g��g��%"Q�ڪ��Ķ����ڇ�d*� efd���+��L�a��isu�!���'Xf�;�gc�4�`�㺆�����E4u�>m���6���=�sӑ˝�z\��J@����]o^�MM��7բ���n��k�s�l��Uc(��w\$�0��ܦS�t�t�)\��ڂ��uyq��ě.Gr={*���w]eV\C/F��=4n͗4�۹�[!)(��d�7�1�kȜ�[�H!�1g��=jx���E�e�4��}N���2��ݐ+.Ԟ�Un^6��d㵚���v���eZ�X'h ��<D��Q��9,|l��;~P��Q�uo<h6��͈ag󼔮r�Y��u�Fܶ�@��3�3{<�ϡ1�+о�D3Ð>�6E��	]��skY���q�q��j��7U�*EW�������?xV;r����7ݯX���7l5{�z[+�MU#m����\!���;cT�@s NےA1X�^WSv�����! ��By`{9�?�^3X�Z�TSfI$��rV���UhսCT��]S5���m`�A��Y2j�"Οػ�%X$G�I�CuQ��o+��6��s:���^�F��gNP�����xf��S�V@(amU\�nTTmK�-�JX��5mMU�ܬ�2���\��D(�U[Wzjn^��s�3�qL[�y�� �xIY	�K?�!#�D��u�=̣,*�b��&n�0i�BT���L����4Y�C���l��N��3��j��1��D$����`NPh����T@{���s�'�������W�Ǽ������mx6TH��J'r�#��t������<'�D=�☹^�{�F>&g�5�8��H�[R6�7\Y�C1X��:�).�%"���^#%E]���ݡ^�T݇�~?����#6�j�U1�ci�qպ��J8\MR��d m�Y���md�ݸ�3ʴVR�]�џ|rm�=�fvY��*��uT��/�Y7�d3��@��k�Q�K%8����Eǽ_����է�:'`�!����V#�S�CT6�f)��ً�;�Ɂ�H�2����ug�#Oz��F��ӆ�r˯��Cx����%8�-���]+��t�ww`�b����=��f#6���t���k�3�*Eݚp��rٖR8�d����!�:�=��Z��/Jg��ď#j�bd8@L���.^�G�}�[�@"�mqUV���6�4&�e���U���*����@�   w)����A�xM�ʙ��u�mT�(s� +����l��]����֦6<���θ�?�ϟ> =r��R��q�T�@ *���P
�u)֭���]�p`�T�Pcd� m�p� 6� wT�mP<�k�ԫmU�n%MC
�Jd�Η��Ҧ꘎ɶ�k��F5 �`�� )��lڵĉb�[P�ڽϺgf����]gz�ȿZ&]�E�����=]�*J���9�ӳ�����-cUU$rU���ku
�Lt��/`�w�k��Jl�4����a�[���.>!�a2�n).'^0�v�{��=�v�w-�~�$f,�<�I%t�*�]U�Ѳ��=����1����u�� G��-=H�+����/gslO��I$.��Y��;^��e��E�����1��wmu-E���3�T���Y���`���3d�ƶ�^��t�R�tKh��*����n\�w]-����5�����gk��z�(�B���aڭ^6�vՐό�8����T���n2�LJ�D��~9��O��r�4�\'�*̗�3g��H�H����7���Y��^o�F4ҍ�)Ő����R,�e�9�����,��Ն�㫭�����U�m�/�P�#mƋF�tI.���(v�'R,�ߎ�I�@��ǫ#1x���m�M�!��K'+gM�����D��~:Fb���J�"�Ex��=�t��څmZٖ��㔪\=�[Z��7I"S2��Jj( �T�T��֭�m6�P�ps{�}3�5�}��?����VB2׏�Ԙ!F!F��i������a�ڑ$�%'q�;������|t�Q��Ef�hڶp����x��q��iR�EȌ�Bm�U��Y�f/.��0��c8L��ӂ+��0���]�����x�d)AiF�Q�����{�_�d���NX-�2��pb�y�ǎ@��_OMOM�{�[�42�UX�]^?���2"E�,�6��:D�8P�C��ܩ���XG����)�� �U[(:v�0;;l�v�J��U�������e�UTb��l,��D�w�����&��f!�B�`��8E����D��ƍU0��kd�j�P�rI$(̕��GY=�C9?�Cx[��^r)�xU�ז��I:�2�����m��nk�⧱�,׵�֥�ݚ�z�7��gk&���pB�<��m���x��f��3������^̊��Z�ѭ��N��w:i]��-�٨�"�w�u{w�&ԍ���-U�Q�ӡS��:{c����*һtlL�U��T#�ɂ��QuUy�?Q�:=�vl;���E��5��n��[O*e���FS-�q�#1����*w�빇}{�ݤ��37i��f�n�)1~���nH%?_n����7S��j��i��|*�ڳ����۬���O����ɑUj�1��Fg�o�%�>�Y�Tp�O��ᇈQ���l�c8����3ι��(����RUw��><B�Ċ��uE�p���R5�d8D8Tfuf���Vx�r�����ϧ�ښ�kj��IR�&�l�)��<U��z�    =l�=�%�Z�c�5�X�r�ʵPVsR�l��K�ڶ�r�Y�ԣ�m�Ղ����6����Et׭�ͮ.  *s-�*  ( 8)fF����*� l��6�� *��p  �U�T�V�5}��h�Um���(zf�a3�-UU�9�kk]�CcwnѪ�7$݁o2 �J�7w-��m��H�M�����|a�V�����x��<vJ�脊ʂ.�Έqg���"����>�7q�#l�lV�sP�V3"�gbs-TY�b�R.��>�r��:G�U$���ڑ)p٥WX���aVKɐ�,�	��h�#�U���b^��Єa���.��$�q(��Vj]����T4�گٛ2yG��HW�ď�Ҩ��'xj�֛-X�[mX6-�vm3DX��[4y��`�aXdx��˕�\B�D��4pݡ��ߛ��#nF���S�m\�L;!�^�F��*�tSlU�V����j�͉�4��+�"�g�[�7Ha���.�q���7����@����Xl��[(��K�7��)�Zh�6c;��9=�Z>4�1�$���C^�*a�^B����#�b�J�c��q�G�PH�N7b)(�x��:�P�q
"ųG�p<Ĭ2<t�nT9}�cL��kT/+T�UT����ל���Ɯ�契��%:��ۙkaSא�0�ܪ�I�L�aR���KqG2'\a�B��^w\l���˼��2�Ք��G�ơ=�{c\a�۳?��(�&~UT�o�ѫ[6�N�o\((��jڠ
��7ucp����it;�F�����C0�B^E����e�l��l)��_�q�������mHV���'��>�u�ώb<�L�\a�H��d;�6��juk�ޜ��GS�P��*��g�kGyx��;�g��Q�Wd:}��8.F�����&��,�����䐴�r�%A;+�o��ZSݛqh��7^!�V���Pcek[�u���-(�q�t����"�ۗ��⽖����yq��\�\���C�e,�n7�6���ܐUUWA��.�;-z�<s�,���
�Ъ��!��h��5*���7V��x�I�V#[��FȽp��CuG����#���D;T���ʥ�D�ۍ�K8��:e��\:�#��l+�^�Pfׯ!��BdY�5�L��ަ�X�D�%(\��\Y�C1_Z�V�?��M�~�~���b���e���J��^<o4��!��J$)�\n���^�������
H��be��/N1�快��V�N�\������w��$��nm�`��Y�W�W��|��zh���Iv>��bo�����]ҵJ�iET���mȰuG&ӵ����ue��K*�YX&`B�͔�=�EU�Ukk�3�h���G�����<𦯚��☷^��0���y<B�}b�V���]{���_C�tΌA�g�6���!N@�F���2x�#;�7���:�AVA
��}��N��C�Yӑ���Y�B{$;ս�'�~�6BH%���pI$�ܙ����k�M�gH�A�f�4��ȭ�Y���R��o�Z�H���TnF��%~gMRO.�x��E�[Ҹ�!���T���49�uQG����D�"���;��@)P���
'�eQ;%@�!V�D�D+��EAS쀠�ן���A@���"�� )�AAU?�������"���������������@QF �A�QTUU��d��?��E=�����Q�G�g���?�A@�����Q� � _�PE=g\D���;�~��띝���E?q��ӿ�E?�E>�'������oG��|� � s��<����QQ�6�Q����ъ
�2�� P���� ���9�>���|��*��UR�*��*��DI"EU"	I)%T(QU
��P�J*UR�QH(T"�U@>z U�	%(P�R�RUQ%)UD�P%�*�EUD�T�"�RJ�J��RI
*�R�UP>�"��e�L��	�W���B����Ի[67����f�����4��\�*<w�˸�T�+��{-�[4���Rsa*;KO{�RΊ����w�fJR%A*�R$�
$�R��x�}֧�I�׵�r��g���ӹ���c�CǞ�+ޟY�w^�/�gj�gMT�*�����Y���ɷ��.f}�Wbo_>U�	�C�j�|��o[%��c��{��ec_,^�҈�Q ��7M��L{Vn��JO�T��v�m�[���:J�>�u�ں]�c����n�]��z�C�}��2�l��n�f=���{���v�͛[I�n�cz�6�K��i�E����_e��(>�uI(�)J��� ���(T���}{�t����>v��^��.q��[���_l��=����ݺ}m�Ď��ﻏl)}Vد}�x���7Z��]S�^mE)K��d ��}D���W��!O�Xǜ;�r�#�y�kCG����|QHR"[��T���ڟX��}H�|�ۏ�]�+a����:p{1�u�j�vd*�;��������%/_7������=���/��/��l
Kٯ���D�o��T��;�;3������ԉ^���_;���ٗl�	*U)
G�䊤UE!E*)���]Rr�5�u���mD�|�]�ݵ�;h�7�*�Ͼ����k���2��q�g}��|���k˫�{"�-�����M�*]:�{��*K������Z�h�_l^������*E�_lg�IUIAI]�f�׽�iU���*s���}�UJ/w}��@!���y�
��w�}��M�tz�H���^�U�t#E�:u��kZ_c��(�į!�{n�lw����U�ϣ�*���Δ�$���)I(�U"�T�US����_v��<�z�U#�K�޷��k�ݽy��|}=��Vv;���g|�-�[��{�uѷc�{�}=��vm��s�����Ԩ;�}�\��v�����t�]�����r᭩��{����R�"QU����}�=����|�����|�����}�zϮۋ�ۮ�Ow:����mi����������{}��ު�����z��М�u���{��ѥ�<�t���%�g�� P�JH% �IR�B���*���G��<^l�]����=aH�MR����kw%�J�{�)UW�(U)Y�ěkG;[f��U�S�qJ^�9j�յ<�D���:�DS���J�� h2S�&�IJ�1 ��JUM4�&C=��F�  � MUQ�@ �j�P�=@h�~c��_��I#� _��ɍ�u2�~��L�O�Ӂ�[[]��着�������}UU�W�{׻���w��������w��w�������w��w��������w{����w{����ߏ������o�C�D��~�&ߌ0Է$���G��*���|�X�)
�`�`�>���
�~��t�L�Փl�A�聪��S���tj�ȹ#Aq�5���l���@\�bc����f�����:�`�����MAR�z�l�-��
7v�穅�R��m�:�!��z�Aʱ�����4��W�������X�k"�2%Du�IցA���+2���<jۈ�f��m�%@�.Pd���d����W|�b-�f�k1>�_X�fC�yi�r�lЪ���i������7 ���Z�a�ě������5��/cr��{����.�$r K�f1WQ�%x+U��l�Su�U^%O�
�,a��#�,Y�yR9������*�Z��C��(�A.]�Ղ����!Cu<`:rб�I��]��ͦj���}pЮ�����h�e�3���\ںY����kv�!��K��v�����Z`s��^�*Z)\{Z��f8�!��)Q�Jc�]�Ώ�:HCTv��ⲥȘ���(���a-��!{vA����Y�6$��ڙ ]=̖R*�ђd�s- �ؠ;���5�z��%�u"�3j�K[��!�Z
���&�ء�te�f��-�x Y��Y�HܺM��F
���jlcu�ǄZ�G6��5l	X��Vj�=������ӣ�+z�D(l�B�{�����N�����`�#5¾n99H}ue����jC�`ch��7��V�2~y+L�T�o.�3 Ȇm�.c��J��"��+2��.]�R2�ma��Q���&��ZT�&�Nٷ5jQ�2�2BlS!p����KX�GԺ�r�w`�v����J6�|[	ܽ�[l�j�V��q*!�e��P��1I*�e��NHiMӪ�XU���c)k�pĝH�Q�9[�sL��va�ҥm����B�`^1sO�˫wAR���\�l]:�e1��Z+�&�9T���� �Q7��P5(aVR��^�[���Ĳfp��-l�a��u��¬]�ѕan�� �8�Hgĸ��b&շJô4ħ¬2������@���D p
�7 q��z�`E�h˅K�71�r�h�2�B�j�FM�v�INR7z6�0��9��!!���M�˫�)#�%l�t��ܷ�$Τ�С�����j�]{uD�rvZys_�Q��]��/���u��f�wb�EF�sr`���w�.E	0��"g/RR�:�V�wSZ�$a��*l7��Q1is�6������U���ބ�rN�+lo�6���S�V�!G�lY�,*ʷ��q�G�vcƨ^��$��j��X&�,zC˚3e�iT-<�U�nV3.�=Mֈ7p]�-V�sw�9곹��qv�2�6���% 7V��n��;��hr��z�eXi/'�����R���3-�4�ۃeЊ����E���"5�3�ng��+���SL����:�.�_0�Q��\�HJ�v�Cv%�+����8U��h1�� +Y;cVi�4͜/gs��3�B򌗕?���y���镢��t�:�X2�S��VJ���h��m�5��޶ҝ����,[�G:cRM���4��zQ�תβ32��͔�9ał Fe޳>8E`��\W|B�z�G��U��2�2�ܖ�S�	��$L�He��>׹���7����-���C�0:�řV餬U�]���
`STi�A:˝y���VIoPM�!]����}�^f�@btj��j�t�j�e+n��;G]��[hm:YN��	%F�U��ٔ]�����F��,��E���%1Cj���0=��� �x�(l��f���"6�Y!�d�Ø�
n,�U����Mr(�46�H07�E�we�@i,�رcQ	��
t�3n~[%d�䔫nTu2�,�L^�Ǹ1�g@)�z-��o��<���*f�pږ�Bgk+i���z��&�cFX:��[Y��5�.G��]�ii��4��mH����s�
�op��1Z�+v��:(�K´f���i�ϛk4k�	��������깦c��Z_/��P Y�҉#Ew�\20�g8ԫ��u��[�*暍�xm�V����}p��Š��e��mڔ�Z�t�j)S���1�Pt+%Ͷ�
q���,��SyZ\���U���A�;2=�	%K,�iI*�WW�����r�f�@k�?�U�joM� �QTɖD�%1.e��M���`�-+U�r�^˦�ͻ2� �V�����ss7k4~>��I5�	���`Qn��n3��4�û��dhl/e�4�\��si���WX nc����8�uؘ��n��K�^J���5�p�o,�t*a%Ff���^4��vOrT&�����lj���-��q]��)g��mfL3��8�k� ��r�GfG"i�c���V�kʆj��I�:�c3%C3C�[�W���n�3�ur?!�2vT���YYќ�z�輼{��LţQ�짆�>�,g,D��*�����7,*�1[�G1^�16�l9R���(�㉛b��a(S�t��R�Lj���r	j���IF�[܇D�]n�w]��RI��X2�l���nf����8�0�ۃC��N�t%K۷�����v���nۧ� �U�`�+fޓ
y'Y�.@����-4j2p�ә�t����� k0��AD��	����fnC�M����\mU�Lk[�i��n#�h���e���6tE�LJ�L���g u�+r]IY#o�H�q�-�(Zӧb����e$^�|Ʀ��h��ݧ�����V��N���-G!э`��[��U�y(��0��T�-c��#t���5�`Ș�wr��V��ܘ�ű�Ee:�v^���3�w�C��$׵(j# ���D��#A41b:��ѕ{yMPƫ$Ua�X��{����w��7�7�؍֋ĭY�a�fh��8H��t�]K�v)��l���<�XR< ��7�+9��Ln�̡"gӢS��mZķ���3t��-ձn|���r��T�Q�����3�'�Vk�����cD/�;�|�RR��������1�7f�e���mh��wh�q�^R�Ճ��]�EVa�̧Z�#�a)�c�ӣ���7R�V.ׂ�JI�m�\�򃄋�PU���WݺR&� � ���]B���6	T\�u[`c�-��v��ɗF�M�ʺ�
��v^){��o1<�+C�2mk�D3[I�܁P���V;֘[K~d�-dL����ʐEX�m�ƀZ�h��ote+�8#{q8�PQ���pnb�ө��ڥd�[)��p� _����])�+�����9�7��,.'���c��M(��7��вP,�J2�Ň��0���!�gB�����]ζ��㫗f��A�Z�5�Q�J�Iv٠��o�}!k]]k���R��ި;(�[6�f��(P�x�nh��G�7oxm��Hqn�̓�E5��PR9yq\7��nA�l^����S�����͛GN����'�jC+tX�G��u�nI+ �P̢��%Mܥ������)���x݊����ayP��S
�l�f�ҳi5ch���)��k@c[�;Ⲧ��Z��d�$�
P�uoU=�]�IVd�E���>L^�,䛭�Sb�b��=vj�w�x�CG+&�5�*gn�ˁ
��H�ŀ4o�#f��<zϣb���ot[���G��7]Ƣ���-�P�Z�l��-Tp;m51���f�v�V�(4�-��:��2��>wp&��;8B�f2{)��?:�@:]�hɨ��5��d#)��ڎm�����a�4h���C�K`�p���Y82���Щol'Rd�vV�ù�VX5���۫�T3�Y��M|N����Zss�&.�	�kw�.VedU��nG�o�^U�͖]7z�h�<0?���.1O���^J�3����b���T�eS��#�kE���SYWOv��2����1��?E5�[,ÀT�ᶓ���"1zɏhS�PŒN�yF���Ke�KKÃkn�Ha��7D�AJ��V���'�saܫ��8�u�Z��k�]M��a���6C��σ�Ѩ�@K�n�Q�)��/^�7!�S��%x�������]16��I���a
�w)T�ً^S�xa �-������Ь̵u���L���D��W@i�d2hύ�7*�2�%�`]l�w.��A{��h4Ua�M�w���gfT���؎�yXj��k�좷�+0�E��W����7��B�h����0V�Dte���Q�.(�V[s�4Eۖ��@�3�ڽ���$����)������VU�[sZ�R!l���b]8֡ ʘ/M��UkT�E�)0��2Z�ra�
��;��j�,D��⓾L���	&���cm�==�Aw��[\����Np�Vh;JV�^&��v�hN�P�ǻ�U�������@>��}�]�\����98N��L�"����ޚ��umƉ��8�1����R�r��i�[�'���p㷅^��z�#)���Y}kl2�p�oB�]����$��ts%��[���7��\���j��o�0������E��FU��N(MU���4�m,�d̫b_H������ךZXFs�U�q�bl2:0g�p�x��%Mx;&�a����S/%G����	�X�Qƣ!��ytƻqu�k�nM�^��@� ����R�,��V��uo	��T�:*�s���9�h��	¦�陑AQ�U��G�޶7E��Gϒy��%���n�$��眰�Sh@:O���u���ڭ�m��U����L9{nC]v��Rx��˻�س��o9 y�4��CS0̹os`��b��]c���M�_Q���b�=�Nm7 OQ�$�N��n����V��gp�ؑV������m��2��C��AV��WGQ�F��KY��f�AZmځo�e��S˼�[�5����DAvtB�
m -â��3����R�#�W�?w43"���Cpt�r+:F�{�>�Y:f^+d�iV[�c��z�/;.^B�Y(*�ﺱJ�'4�hj6�K�O*���؉f�bno$����W}^���K5R0�����(8��ݳ3�����:���� �_l��L�l�ZYg`l�*�ZD�4�^�f�f|���DPaM�`@���WSi2Єn�`�@�ư�K.75T�y[A�A1� �5�P��Kt<&���B�ι�nM�S\�Z��ا��*fɴ6�h2�H5a	�m]&7h�6Y�kF�vH+�T']�sO\z`��Ty����3c�F͝Zȕr�t���w��P�,:���nf>Vn�؉�PF�d�{����Ѓ��a�55鳑�dn�j +r[7:2Y��i��Y�#x���)(�`�^KUi������e��`6n��H	vR��Ud��/��/]��D�
�M�Yb��V2�l�NA5ԛf�����j�<@�DI24����Կ��K+vn� f'�����ݼ��]�(�M�8��a�nZ�wz��a�{�E�%)J�;���V5�3S��$���1%e릊E^��^`t�21����aH�V/(TT �siӴ�)�;f��J�YB��N��\kEWNQtW׃2rX-�<kg�|y􇻲dݳ&�R��c�������H����E�ݕ��7������;?*�D��U�[/$�Z���� ��;P��7/zZ�ck��sVI�^�s.����n�����r���ŉ�Bܳz����ݙ�L|5���pl���rzBp��nk�E��8N�m�T(�ڴ�%����JŴm=�u ����,�_f_]`�/c��X�!�H9�Zɔۮ��s��~�S���6���%�#.�K�nUЏ��`,�}�T������zz�g�6���y�T���5|��7j�ʟ�u���Ǯ����
���c�#*��e�wA�"�\x��u7����ӬU������o�7ݺ�uw�ߕ���n`�y��w��!;[�q1�S+�1��m-�9�����T��^4�ӨOeH'a��.v��|�9Hu�o{��Z��63iw Z�%p�Y�ɏ��%ӳ�s��6�]d��a��q���Ё��Y��|��ec�R�&��p__];g����컙G;-�pW{Z��Ʃ��e.�En"�(F������骎�=(���ٛ���ܙ:��͉��X��tFn����+G�iu�+��su�:�
��Xy�NC���<�uwoT|-��m2�F��c��4ok�>0ҫ�;1C7��.v>��A9ֺ��P��VMV��}���9.Y����;k��)A��M���ۻٹձG�[/��Q�qT4�ۜ�p%��ؓF��f
G�-v��:������75]p�j��:�o���\i-��M*�_C��%�yZ�6�u�0|�u�~��a�,�e*�2�v��hzd�]�	��)9��E5������8��k�-�>E_�Qy@�b��S2��om��E3	����" �X��-��l�P�r��G��u�&��/�S6�,��{wK5Rj5Uɯ(mٸ��E]/-�s\�e���]Լ�-���j��N��y�D��hkv�XY�ׁ�����A�{p��	jI4i�mrF�R�u|vuAǠ�I��n�������t�v)p�)(��t�IP��;z��.�c����jsws0n��#�J�6��U�T�}�gթE�����.�wz���(��c���i�0Wv%���%��,��/c۬O7�����X����ۃc;Y����������1�̵r�f�+r������O�����paݭ�����U8�E|���e�vw�z��C!)�: �Ҟi��`'q�b�/`⫓�7Fm�J:���Be�΂���j��1Q�.�H�C�����,��P
-�R�TR��R��UUUT�D�R�*��:㎸ �U.A�J��1#�U!��¨ .�^�)��l"�K]+�m��^T�d&�ny�kQm��>Q�dW��z�6������a��h4V���R
�]���`��Ke�UnvP%`*��$b���ePZ��U+	(�2�š�'�N$,uN�=SZ�"����(9i�2r�c\�aΑy�h�%6���v�M�s�%���ɱL����N�mJ���nkg�^t��UU[����U*Ԫ��J�*�@!5U)��`*�*�I5U:�-[���iCV�Ύ�Ñ�SÊ]�Z�U�8.cbz��T�����..�<�M��.5����A�uݝ��'
F�n��ùu/�n'u#�um�Ε[7Ǯ^%뷋��̇W�6��9�Sب���Rb�SM�{]R��/=CE�B����7H6�1Y����f�xtWHa1�&y�hD<iW���=lT�L�; �Þl69���oß2\$�!�-�����v�0�q\�=���a����7s׶ݮ9��u�{��M�%�9�&.��y>wc���S9�q���;�3ۊ�a��#�P;��`�mZ&�n��n=�sw^gep��A���E�g-ƹ�+��OLsq>1�ʝέKŮ.���{2=c���m\�!��k�yǜ�:�pu�Ɍ���=z�wK�`CFN�t�3�ӗ��;<�x�t�f�NT ��{v��Ⱦ��뱊jx�'y��Bh�e�9�kNQ�Q��v�cp�g.��<b��џg��:}]�^5�j�@�q���9�}���H��u�^��;t�ט5ݍ��=�s�̀��NF�1qڹ�)5�s�\�{x7met��m+zf��(06������O]t�.�<uP�@p�����9��Z�
9�+8��e��`�m��X8��J��s�hN�"wf\"�*�lv"��	,�r=dKvq�����F��E��]�nۦF�떻y\\�9��v�h�ɶ�{����'�'>����d��yz���⛦�r����ve���$/[����T�u���9ܤx��㞗����7;�1ܙ��t�4t�M�g8���vEZ[�c�z���ۮ�e�mȫ=��N�9v�^=T����ڃ��r2�^zB����Ս��Ⰲ�m�s��si��nM�l�H��+f��������L�z���c�Lpɔ�&)݈�R�,�]�*�@�
w,�Hw�A�kU�#�k��';�ϰ(l9�q,�r��7,)]A"�8d��s7A�۰m�ƣ���q۷6��e�u�9�������g���RE�� �&�����9�9�z����g�ގz�UF��ޗ����">��*c��[g��N��:w��{p���,���Poi������x�A��nh��g�[ݻ��m�S���u��E�qfl&�z`G����]�I����'>s[[��g�c��n��Xu�\\�˸KX��y�s�j݋�\�=<�r�����[�w	�{r���=8<��q�a$y7=)u�m���=�|c+z�ݞ2��u���z�7J���;��=�� �{m�6�89�7V��.��*�㶩ǶR��;�ԉy�G���7��e�E׮]�n�{m�67�:ꇺbp+ K�v������l��sװ���[���.Nx��z���R��۪�]��c��^#��rx�ח��Q��܆��8���n�v�g�2rqÁ=��۞{Y����˳VE�u2v:Bm8�r��=x00����xa��t\��-\nw1��]q(�ls�y�n��rni���V�s΍g#���Nwh�Ng������v�t���t�;�����)����7#�|C���e��<e����0FϷ�p�a�y�SĶ�[��r��ǳ.�YY�k�s�B�B��c��#8�m�;bMN�9�N9-���K[����mvA�s>�[�<��3�ObP��b�A�`��
��v��mcsn{[��ʆ�B�l��v�ޜfD�s���ϨHR�0���\a�]ݝ�\z�W>�mx�r�����v\�w.�#͗<j�뵎6�3�Ȉk�,dr��.2�֥K�ݕ�Y� B#�X��GkkY���6�>�w/Z���v��A��*�ݍ��$+н��#�99���Iv ��.�s��p���ɣK˘��㓡:�幣��B\Վ^qc���A�u㎓�a�t\"���9�m�Jg�x��;BG�E�v�!{��'^y�vp������nx�ۜ뷶	c*F�]�n��s�˷�N�m���qmAp��$�s	�vO���ї�[�W��V[LE�=��wW]���˸y:^���ݎ!���s����p�s��O.�=rV������݇��n�\lNA��X@�e�@�7���3[<��63vX��f^3Ϲ���g��{���&{��uc�>�B�!����y�j�Q�s�=���������<Kh{Y�فt)���T�ێny-�k�[�yl'��98�9�2�;�-��Ӎm�ǍBg���7gq��F�7�M�,�du�Q\8��;�<WY\'Y�vwt;��a�/sQX��N���ps��2.w;��#p��sp@���v��`$�gӆx�(q�-��E��v�v������<I=u"���ܝt�R��Z��Ի��Ϋ�mĻ�B^P�K��|nw��ݢ�zw9ص��/bl�upo(
��ִ���83����O\ -5��c��]�Gc��x.���r��6�k��9���E.�&`��]r�7Wh*/<L9��J�mv6�ei6x��g�i�\Η�"�;��n�b�S=��7��8�\F�ƽ���̙8�W����{;a�W���9�:v�B�qnݕ���`!�E-�V��JL]s�p&㢹��:���r���G\8u�Gg.(���UѠ���#�E��a�kN$Px�W9釋��P���5ѳ���X�^��O=6�']��D,�S�}CM��E� m�K�T����-�ns�yu��g��m�J�q]���;;q�7�B��%m����E�9���0z:���-��
,��r1���eF�t��M����h�s��҈p�gz���t����Qσ�˻m�km�]�O;k��X��� ,s�y�W'ul�@���7(v��b�n�sV�a9����rYٽ;��n�#�oj�:
�K���ld���㣋>���)9�@���p ��˭�"I�zU�/������l.�kvz	�q��7��6��+�9���[���u��L�jhx����F��G�N��L-�WZ��a(2�[��w\c�$�#b�wk�u��6`�K���+�^v�-�APMu�W�]��a�`{�{�m�`���c�:I�<�]���GW\F9�s'nH�.|A�O���h�c��s��rE�75]�Z�.v�ەdhK��Dtg�ۭ�MZx����
x�NDv���O��ە\�u��,�6�ۓ�u��A�����Bc�]�..��콶랍M�=^j�7i���-�9����\hgw.�)p���ڎ܇5u͗����{���9=��7;/\���ק]9H�닗�Gm]nx�pk�p��u��^K)�-L��%9������/gH��qt�m��p�9�O�5��	��j\���a���a�p��uv���w9�u]�=u�y	N9����u���Cd:[Yi�vLݩ�=� 9� M��Ź�8��ŞƟw��k��p�@���D�Z������|���Kk����vm�:��FiD!���>-ۇ%�tt��n����+Qu�k�s��x�v�Mu�z�k\�x���>6�M:��H�D���g�8,�<<�c�F������Ç$2�����o]��;���W򮹉��x�6�^�{p2H�i��X,��nBv8ulU����1N��м/7s�a78B�u�ۏJ�R��nx'`!��|�g�P�&ˌ�%�.Ri�\�<EmgռV���c��5k��{u�gGW����	�e�y��g�c'Rz]nc�lb�C�<�w �ً�����a+���h�tj.�V��9�ͦ��v���g�l!x�9MZK�W;���Qa�N����z�f����\n�r��RF���s�*��2s�����3۬�͹x3��wf.;�Y�p���vnD�Eגz�Gd:\l��эt=aqYy:�e��KA�{�|\#�׵�g�N�8l���n<�^lO;q��](Qq�p�6�F��/[�\u�u6��j0l�]��7=s�a{m��K���`	�=���l�V�nf.���4�`�s���rp�����u��<��
��z�q�z ��m�>���ݍ�qu�尜�W-ٱ���T�i��^I��nxvg.Ջ{e�G�79�[,�N�n7#۠$m�8�aNSN�h�*z�F;1�]�����gP��M&�#\��x�X���ٛXv!eݺ�3��OB��cW��Wr��`�e֬����������S�s��h��ܛ�y�nl.6��rP�dݝf�K���W��wa�4\����neN��x�7*��{Cv��ADv歹���t�n�:���vQ;�dKI��:�u�u��A��ca�X'r�d|&yݕ��3\����ǜ�r�8T.�wU�=�iup]�xKl:� �:^xpn��'�M�4�빷n�$2a&W���%4�q*t���^�3�*�]p�N׌\���&R2Z��<����S����s����]𕛞�+��yR���㛵�C"�t\yW���hB��{^�nM�f8���+��n�q�
�n]�ʚ ���wiB�7t�qtv�ۂ��9	�`Yi��>L�{'2d��];S\��I�t���gkJ�kpe�Ѹ$�ǰFV��˗��&a��(o,�"ƸSd���L!����ww���{��������w����~�w��{���������Gww�����^�ww���x���������{�����p{�������������w�������;������w�;��{��{�����w�������pww{���{����ﾈ���>�>�#����?��&����
߃�ƕ[��f��Z*X]qҺىw\X��WkW���Tս�/���l��Ӡ�	ө@|we�������>j����s=�����״����XCc��WW���S��uWq8�^��d�!�ǵe�����G͢��H]��{�	�q��h-���J~�j"�*�?��K�yu��F�5�T[�4`�g;(��j��3�^�!j�ْ�5œ��Z�!{�S���t0�Ne�\:%Q� .�Ԩ<���o� v)^S9�oo�7�NB$A"!�
����\rvi�w^� ��>0L2KhC�io/uj�S���ք/�z̤=B����v�g�L����o���sy�{��{@p&�g�A�����`��H
�G�0(�2�=���Sޮ�]�����_<+Ma5��X�,��\��h>^p@�5���t����{D8����@9�� ��%���3r�����)߫���Y]���{�K�t��c�j�o�;���H�p�8�zG��{��|��z'���h7M�m!2+Nҝ���a����"���ǰ��]̜=1	|}2���U�b�����B�c�|6>�f>c����X�$�;�,�q³wyuŘc��@�A�u;i�Ӕ����K.%��
=�u�	b-4��Q�Ƚi���b�4*�w�n]� �fx�%�;qОptF�'W5�sx�Xy)y����x��?t�GKy��\�Zj�p�Y퓎�9f�웧����C����g�69׳��X9HP{�sp��!���.p�t�j;li�9p�wF��e�t�盲�Jq��]K�����:��H���Ğ����θ��;۩7`^�8��y���W~�
ֆ�O�����,�)Ɇ��xV��:MS�2if R�6ݞ��Ѳ���Sd��`0�1��,���°U^B�g^v+�N8�Y֟ά�{�ؕ��U�A\���"���/v!�",P���8�&�JNcj<�1S���W��QP�	6JFZ�7�n��R���"k���G�U��+ef��DSt)��`�ic=�!ۛ�n
�9.��scu�4�<�\L�.��zk��-vM�]�G`Hl�u{b��>ۆ��x��C��[l�@h�ӌ]Y�+�II�i*W��Q�	�svLXy]�u�{+���:Og��B��vm�N��u>DIӴ���ÚE��r���Y���]��p�f�dכ4<Mޤ�m)YKJ��9�nѮnw)����=��[��{YG�@�Lg�S[m���w�)�Pn����fJ]���W7��zi+��<�����Ȳ���Є{��8��m���)���'W�7WZ�}���Y��9+�9�x`�)d'�畆b��2����Z��v�����p�p���^B��6D%A��1z��Ua�5���zMw�{:��y�WJ�n-x~Lrی�Îԩ�aI^�Poh�s;���q�u�c9������xT�v*���Ql�hS�y����]r L�@[ݤ7�"���wo�~���S	���t�yT�74 	�|�&�T�*��z��w�T���Ӛ�qZF���JB� �A� �WvmΖ���tn�3�.ۃ��3��uu�D����~}��{n�ۦ�f�Ze�s�iï�Ir��nˌ=�7^�Y2��D}��x��zc�
�(�Ue'���s�41�LR{�c��z�ޙ=f��V����J��#��s:�^����CA�=/{_��zz���fk���귺=f��b��G���纻�j.��̓��/.=��e�B�����=���pDX���ƽވ��HE��=Bj�Gѕq���A�v�ظ��J0�0]L5¯��&�Y6jʕ��-�{+.Fz]n��/iJyv�����X:��p��*�d����n]����8�pkգKa K�
5B�>�=����S\`����K����
�g���X.��:����nK�+�k�=��qR��%d��s�JvX=��I�_Y�����:eR(0J�G�{^�Y6T�zV����̘~?�"*\�qK�k����)�@pM���q�{Gv�) B��-$`������MBZ]Êa����5�T�{F�loʤg���ю���2���A�{k�(�a׋�.��p��#�����bJ��Fۦ�\��x+��Պmn�ͺA�^a*��]��h\�ר�MPiңN�Ky�ǣ}�@�Cu,^~�2�]��?Xɝ���	v�`�^�U�`�dEXu�,�<���0�8����_rp�)��`��E���]-����5����7�B���F��tܛ���-;�Z�}��Nt^�󞓎L��{zxe�.�6��Ic�u�V��s�H5�@Dݥ�c4sܩ�=�_o�x�}�^w�V�Ϗ��:-�R�[��jJ_*���`n-xk�:���B<}q�A�.}7^/{�����'�4�T]?)Qm�쮠��̊����7��3Cǹ��t�{�=Xn�=n��5�g0Q��.���{n���{m;��Ů�-�����SQ�� l���3��%�c�:nzzT��v��Ί��t}��G����+�x�֪�sJ�Ƶ�w\�97j\����m�"k�Vfn�BI��ۂ.��4��3�"��p>�ʾ����.:ˠ�x�F���35����0P̏l�9T�"m�:n����+�u��on#�����We��W�'����m�?����Sپ��i��������]�Y�]2�L�ũO�KRi"p��7sm��9��8�)vዄF>�(]�����d �]g:}Nus��x{�oeZ��d��V�0e��b�zǶ{ޚ���]4��2R�Xx���W���:��jM�n������<�WL9��`�S��-���VM6 ���Ad r��B�r�3fe7+v��xy�܈knR�P�{Y�ۦ@�͞�5�Yp}��k�zd��&�\>�=Ǻ�Y�{+����	 ����xw��Al�wV뽹d22�[�?n�l㑙�c��.�T�Tw�:���חJ�-�Q��H��H�Yw��O{Ex����21�w6�#�ʄ�fK���7��
��Bw- <m<�o�S���LDt�7 q���W]��㓜CMAH�Xޝ�ͭ�sf4{\
�Bph5����9�;;���t�ǡ�.����8�	0�$�*c+p�r��mz��x"�Z�5�8x����g�%_�-Ɗ�p���N�A��q��ηU��@�\��hF�b����Z^J��@�O.�y�}��x���I�׸��W@�>i��Z��Fƛ�t�	G=b7"~��n׉�d*,�%'�g������~g�2h��ۮ����
���cHR�Yȭ�
�D��3�~|�5��S���ov�z?xu^6x�������B���ҳ�l4"��.�<�e���֍�*����`l92��zv���m6���g�ʹ��{G`��*��c=v����}��5���Y�����ޝ/s���PK�kX����6(;p\cT�sq=�d��[<6s�WO]J�tY�nβ��9;Jfxx���Q�qd8��6g�����r�v�q�Co �Y�\��3�v�.��Ns�	.N�~�-*�5~�mI�ݟ���1�UR�i����=��ȟx���ҀEh6����o�y�g`f�s���&�������|<]+�K�oϯ2�d+fݹ��R�2���f���[/!��
^�A�;�]^^��LM�O`��R���2+sw�vJ��굁�{���N��#���I�n	�;R�^״!�ۣ�%�zn��S�qPqLk���+�!ʌӋo*��s���q�Mo-Ӝ({��X��H{�#�q>�i$�`&k�4���V��&>d
�x,vC��Iϲ���Z(��d����Y��,�:j���<�#����N�l�f�@�m$�(L"�G�(�ۯ?{��ΣØ��|/Y�����V��q��=۸�w�#نL�s+}҈,m�z�$���V��2�׆��=���ȦJ$�F�I�rE�S�k�"�����v�5�l"��Ν�k~;��:3w��6'd:7��F���yY��<�_��c�-��0[e"޴Gx5�{�<Ǧ����X�w�����I>���s/�c�a�S�m,�m�����eC[�Rfd�Ǚ]׽z����n��p-P�7V+]�l�;���ѳin�n(���	^�ڙ罕���+6bȫ�ᵼ¢�	Pl��N����*>��XmN,{�����sR)��|(q)��0�@ӎ�,fm�C���ȩ�Y�-�Y)�"^�/ۗ��Vыo������Y�咊[^*��x�_f{�f����:q�W�g7��ӗ� #�]H	��V/�ݗ"wt֑L	�݆[�lq<�,*�0G��]l01�S;���{:�<�}�ה�C9��>�;�S~��ȯ�L��V]���e��sN[�>�L^���C���V�`j�5Cջ�{�Z�R��=��e���V{k�#ׯ�]���kΏ�X�=h*J��U�4}93q^z׷����wSs;>��Hz]ك�Z�`�����tO�ɕP�ˋ݋�k6��3�A�	4� ��5�?no�6�������ٍ&e���k�J��]�N�ނ�TЙ��=7���A��/��<Ն�l�-5RD6�o���3���k}K��j�M�^z��[s�]C�|{:�^X+[�G_z�,��<��||���O^�s{v����x�O�^(U*I&BC��D�$����L��ywuM�1_����NeM�������*!t=�)�����k2�v,�Ƹ�n��.G�z)�vJ��R��nh����L�芒Pj�U��sESo�x�8��9K�wy�C�i�D��e �T>��/NZ�#�W�Y��C�`ٻ˽�p`�-{o��kԓk��g�t��v�^��Y�NZ��p���|
��ks�t2��i�ʾ�e�����)�m㵆V`��|��;�Y�ku����ٰ��h.�&��/�	pK��NQ�z�h�JhM�H�ۺ#INf� ��'��맙�/c���� �t> �b�k�ͩ��OW����.)Śr?(�j_�Qt����g������W+�7�?����e�7�8gP�᳽���<���ͷ��M;�5�ې��l�����xx�LPme�=��=�����"ʽ��]�������x�:y�b��r=n$,lvzS�[[��^��b]*B�?�E��g�Og��l�����)�p��n�~��t����v\�j�Źƶ�V�#�%l��* !j���ޡ�k����������$p�¹�?��S�xʭuΐ�
�a�qvz`�wfP�;i��[�M��8��,�)6¥�`Vg��x��P��۞�5�}��.�h�٘Կ���i�z7c�y�$����k�3���@�1�~�L�V"WE}�Bi�F���J��w=������詤|ݖ����n�"MY(��5��!NP�y��8����߯��\'�4���l��9Y�m���{Kv*Gx�S�e���n\8u
�vh9�V�,t^�ٚW�޵�L�yMni)��E�����~����\3�F�w�:U��L���<d�;�K��w�}�)���:~��/fv�J�/U���]���7k�d���iR���{�GG�sz�,�[^����f������H2���C�R`�.�bMF�E{w�9��ru��N�����)�Ӧ�G�r5�~��%��[Rܥy��}������/���J-X$�=��D���3��p��lJ�_g��G5��W�j��g�����mz�F��\K+�B>Ĕ���G�ў�����k�{���k��
������!%�y$T3�2Զs��	����{Q?A
K�B��3P���b{u�.��qjO1�?V�9�#Dϩ�E�_�eIv8Y<I4��4���[�U�@��~��v���vzӜ=nf�)Չ���t���x���gB�i��\�4�<�o�����N�Y�ZB�Ro�I���o0.�[�m�4n����}�1&3�s�s����\U���铥2��xE��Cb;v_k��v���y�=�c�{p�O'!�냲��Fte�k�xW���O&<p�������M�d����7u��[	x��t��U�i�k�.�㛲ogr�n�K�YN�ItGny�����.���iM�ㅍՒ��K�.�b�*4�M�Q@T	�{��f�i>Q
)����:���P^�R�Y�(��Y��bv��=F޺��,@;v)��F�{�xQ!�&w�<��'�'�N�E�~wS��{�v����)��{��G��i�K����s<��>שqN�u�
]�ݐھ�{��&�t�3��^C�X�l�j��|���Z��T���Bî�X�Gh�z�n˒�+/a7"t��e�+�Z�5q5Vq���D-��F��_��,�qߠ���&T�[x��x������8<���Y�����w63b)��q.�m���/v���1�B�w�v���4�kvYbNa�t�^(�Ð	I�`�[�Q��w��dޯ,�i��d�eJ�1̔N���d/�"��]y�4��t}��ڽ;�b1S��vZ�3�ޅ�T��i'�}u��^�����uj�[rE2�ί	���o������)��_�en�r�����kFTC�;����k�%�_@6���m�teFv�܉���^;����5C �ki�֛�vW��}�@������ͫ�M9�԰WuD�,��j�:l
��
�p��ud��z6~}];��f!F��]ܥ�M;��{��v�6+xrX�Q��C���e�>�[�wP������;;���yN��@[1Cs(a���6i�� ��Uם!0�g��Of������+���V'�Z��өk��Y޶3KU4�ԗ�t�Zo%`�;5��M��X5����2�^PU;.d����FSڷ2�r�;���v���N�`^8�3����,�.�NX�Wj���r&��5��]ZE	DV���w�{j#7�Iw�X�B��p�o*vu��Y�{�7FW9�����3b�҉��HX�@��w�OAG4�'Z���q��dW`���S҆ujn��l�k�_SV��f�����L��u���"�|ct�Ye<֚"��YYܸ����_��7�q���N�{�[�w��m����KH���cp8(����g���}[v�_�{�ޫݛ�y6\V&y��� yD�9�_]b�`cѬ_U��
k/���ֺPBl�`JS�)��wK�ɰ�L��֗[B�á���WS��4t����.�;�J����L5h[���R�a,��������W���;��r�ɺn��Q$;��ֳ����t���w{O��{ך%_�h��\��/�� ��4�ج��6]�nt�V��4nU�2��,�)�T�W��;t�4[AjX\o��f9Z+o���uC� �hI��U%mM��kF۫�	Ҳ��:�R�٪�$̪퍞aѤ���.���ꪪ��u�1�M֪N�2�gN�d��ˮ!8$�NQ�rnd����
�U��1�hW��`�k��yt;��r��m�z�}u��g��Vsu�67������\U���H܇W9:=�\�^�Cg2�@;�����v�mQ�kD��+�Og�tD=91�i'�����G���MX9(7�lDo�5��yۮu�t�� W�v�N��d�V�;�ĩ۵�����7V�p���A[�JZ�|��:��<Ic�9��zZ�;<�m=������9�o�5قڶ�˲����y��ûs{O��s�^{={fO���gv-
�rvន���Z�"��"Qb5\����3n.�6D���Y����v�Ґα��;��Pwd������u��)��Xq8ݓJ:�]Gd�RnDTv��<��qsګcB�����$�V��e��{<�W3�v<�I��#�,Dlqk�kX[��t8�^��s���\n�۱�Xv�%G�]�:�rr�����Eӱb�^˺�1��A��Of'#۝乍�<W�ݷns���#Ϋ�\BХǪИ^8<��ո��78m���C����݅��q^d㺍��F7<�yq�ݐgt�c	�:�������nE�r/V�C��Xۻsں�:��4xg�����*�Vn��\��!�Ge r���a{u>L6(I7�����oc��<��H�͕|볰mp΍�����<z�)P�8���q��k�8���]ݬ s��9���wj={{j7����l�]9ޯk���<�n�A�v�����q�ln���J��˹y���uٸ�9v݈�>z�,u�B5�$<.��S�<b�r���laxm�V<��2[euR�Ľ=���N�1�۵��e6��\8U�<�ݬn7&�6���S8��t�v�n�sO٢l��8��C �(G�#�b��n��wQu�>gr��<�x�|��`n}�@	4�a0��*<3�l�J=~��˕;��B��gdZ���!g�nx�4��-���I�(��p�BN��7PP"L��5��8���^[����u���2ui7��.f�u�T�{Aq�}B��n�3��MW{�,W�n��y����H6�A_"��Q��SY�T���3N�
�GYy`��ݽ������73��)���gt���9ʍ^]�����U�S�k[�y���s�W��Vnp�6X��8(<`Y㧓�aq�S]��`�yY.���|����ͩy��o�teؕF���k&I\�3����W��O
���S�L[�J����FcV�P��y��fd󑝞D�0�I�p� �o�T+�-:s}�.�K���щ��>=�>��)��	��݂��5�z�����t��V]�S�K���f3ȏ�)���A�	T����<������79��������1����^_]Z���Yn�8<Y���: �W�3Ċ����W@�P��}G�������2�mq7�?�Ҳv���E���Cq Iس�=�������.t���D�O,����}��������Z�<v�n��=B�K�x�=���Aq�}���\�FEp�i��F�����c�_j��Oc��6d�e;�~vy���M�Zd/�D�I�7�54�D,Kg���\�zr�ŷ���X�fVgMv�gh��-;���⚵���2��Iι3]Kԑ����QB���+\���]=�t"}���aaÂ�:��H֛^5�s�QPo��)٘&�����	�^�t��1V�Óչ)m�#���2}�ؚ3������lB~��PX6	�����M�Z�a�{Y��ߧ�̔�H�RWr��yO8�TŒf�͖�c���uE�]�#��fa����VS�tf���Z��/�����^f��@O�ǉ�|����+�ߍ5���Y[����t3����WG�Ln��w)Yq[��Pk��s�vkKU�+g�@��,�oď������H��Y,H=��b�&&k����}�w<��u��G��J���ef�L������c��ܞ���b`2N���'�>?���-�m݆^i��~���t0�0���Z�ƪ�WH�k2���`�ef�ށ�����ߧ6C��c��rj3ż\Ngj���N�.��e��D(P�!6����ݻ��D��gLb�;���3r3�Lv.�E�
�W=L����7��:���vKܪY�^]7[�QY~ a��I�'< v�/��f}��'=ٶ���w�D�f��!�]w�eʷ(�`f�`���+���⾘c;�kW)i>�K�݋oNy�>�4��|iӽ��Y�ja��M�y�,<��ꠀO{���/g_z#N�8ެ�F^ɧ�E-��5B��iC��l╈Q��N��Z0�Ԥ3�6˳3W�<��X�9H��J��_��*�ݻ�g|��~ӗ2��9�ޙW�����(�y�}�emmȷsV�C�YyW�3|L�w����a�	�%�%�닓2m�ϯjE=�S�,�z|�2���~�V��+Wk~��WRJ��b�Ϲ�aaw��PSȇN��Gw�����h�t(	��}�Qe����HZVf����S$d/)�S]|�WH#��`��Q��;:��7o(�k�����Q�AΜ�~,w�cY[��x'K�W�Fv�ګ��)G�Ew2s7_��,3��>P|4�Թ=�ٖ�F? #DRG/7o\q��f�k#�5�̭
:�ԑ@v���AA�+{;��j�9����{����<�Ź���4�+����Hkd���KeULY<�.�x<@1Ѱ�p�6QƏi,�廳�S5;#;K�n�<efx�G��}[k�Y(�h��+j�gP>���B'���܆u���Z}��)h�˼��xq�R����Rr�4��(���S�y�v�/�<�'��`r�Ι���5�Vʿ,��	��:�sY���11}sҨ��D�i-�wP�B�vƘ��+�`À�2���p�M�M��s�}ܬ:�CU�:�bs�c��N{�����Õ/����#ʜ�c���D�z;�b��%���V�V�p�
]ƞZ�ȹ��\;����Ͳ��lt�ǭ��<qnG\�N�����k��:< ��zx�g��:,:��޳rv��n^���r���ٛ�w�h4Z�vG��:E�����<2�`w�#�v��6�������3pز��X㗕�Dn;sŶ:��(y��Ɉ���B�)�SL�ǝ�7'^l�m�5�m�4����g���NZ�]sG�����n����᠙p���zj����d�ɚûIP�Q0V]�M�6yy.�oE����8.-�m�'�����c0�^�s�\읺�zp�4�hB�]\����.߅�RI��2��TKW�l6����\zgn2��ͫʕO��|8tQ뺩�^��|�.p�AZ����N^7�rn��7��qu&~�|��q�
�G
���ܟq�f��tНH<��e-XAv��u�c�����h �-D6&6�-ѵƨ�'�P�G���#{�+	�k�j�P�cʑ� ��rn=�m=h�\��N�u�I.�e��~�xhl��|�߽��������ĥJ/��W��ͯP	qh�+-e��OP�k���HD�}xT���i3�R����dS�WE��l�}��̤���6�
���۽'��%$�Lz���sd@6o7=�J�eֺH�1]�F���hs�j�3��e_�&O	��tQ�/eQhue{퀏 �W�
B�]���eO�MO�z��7]H�����˿\�:o�����t��ir绰�
-#�D�Y�[�^mi���s�Я%�p�~�u�sO[;� �e�uj:A}��Ϩ��V�uqR{�V&���0yVQ3k�诇��o^*ћ)�~��wt�}T��w�gn�;؝�2�+w�ƛ�d�#y���ójޑZ��_Z�K���U�t�WU��"h�(�j:��m��Օ��kW���Hf��,y�[L}��NN��7{E���sl��N�\_��}�{|��,j5�laKh>�0V78~<~��KRa�ad�����8;U��ܕGA����8��`�L���=��"�w9�
אt��:yܯN��D����d�?yg�j#��p���k� ����Q=��"��Y��J�|����S�^d�V�!�FT�>��	�TV_��q��~�¾ t�nvF��m(�Ʈ�K���9���ѩ��b��b�p�%`���:�=��kGg�<��)�n-g:|`d!��{�V���	��u��z��g6�q�N}w�Z���C���7��L��0��;=*��Y��öa�������ϐjn�z�p���P�Hk|��F�08����Lq�����f}��rsE���kG��m�&{�{Y�f]�����$���+�~��ĊJ�4WfL�PW�e�P�+|<��f�w�
j�#���D�����@<�ܝ7޵���}���7=S4�zm�"Ѕ��`����=��yMs�EJ����q��۾\B�!���3}��y�%q׼��1Ǵtr�T���aߪ%`@,($C�<��f���/n8x�����nθ�@��������ԅq�7�ٝr��U��q>0�Ok�.�]�v񪇯���:ҝ:G#����3,��qb�8v��e����ZOT��z��y*t
���I�W��u�J�i�D>�My��uN�W�m9�Y�y"M@QJ�S���'k�w}��8�<T�����\��|�t]���M�R�s���[93���y�%f6��$Ʃ��������:0��P؀�#�qfO ff�nb���Po�F��+DR�[�FuncRjg���	^�CMڛ��߭�����0�#�욞��]�-\r8�D�Hhq�r<��}tU �
H@��|��Bg�o1�Q�6p�/���gJ��}�Ӈ=?w�gG�>�W�5�m�tga���;-�˕�g�Ya����hly��c�]�ۮ�:CE�[E�l����|[�9 �Aޚ�ҷ~�ށ||�K��p�=�щZ�7���1S��H�)P�{}��Z� �X[-��J,̚�됷����9�DgB-4H4!��k��&���s/%����������y���|���u��
��sQ�����;\�y7Ir�tR0�)�D������EyL,2(�n�<�����?M�{;��c������9x��r������V��
 �(R%U���Ȕ�jl}�}��h��g������n�`�S߆����.sH[̡�Wu��<��km��њ��{<�fw&G���Q�d�mw���l�\@.��*�{'_g�7����o1�D��zՑ��/}������Ï�����h���;Oq�X{�U۸]�+^�v!Y�\2�#�Y��H���W2���E�{��r���Ҝn�������l%��l��;�4.՘*��ñ8nw�/�J�7�o8��Q~zG2�U�����JSq�zՄZ�{~����
�2v�R�h:B�6;:�O����[%��LF_;
[9�����(�-�	��Ѻ9ZVO3�^� �w�S ���.�5�YA�ft�;ze/�s�=���ܲ�/Z�hw3�{�N�y�7�D�,�] �n�N��>ZZ����B&�	���=享z��X�G(ȹ��u���B�$�ۀU�x<9N�5=�ꮹ19S�J��D�z�����By�B�� �(2�T ��{qYQ� k`�X�ypDI�R ��I����^�ҝ��e��|6�l)���Llq�Uʵ�P��u��Ut��"d�t�'ޭ�V]����8A;2�m��8�I�Y٨<����ؓŝ)a\�}��ǵ�;�4F-j�'��ō��� �JrE�a�~Z[��e?'�{0`��/7{}Q�_^��
(��h<��x=ܟ.�K�Ɍ��[�����>K�x��L�a�}f�'"���0n+��69Z�õשNLt¤�vL��'a��g{��~�.��3� -��!�lA��Q���p2;�=�o+[���hk�-{z�����6�#A{�>�bp�yF�R��qfi]����#o����锠JҜ�e���ұ��^�f�Mhl�u������U��ûjyc��\YW]#\z�냧a��x,k�ȩ�0��<�n쀙�(Ɗ��������۾�P���OE,rY�Dpܼ�/��;�ZD�h2X�g�v�6���i�Jv}�lvN�L�7���FJ��,�k�d8�a1�ijώJ%���f�2%U���n��KH[�nUu��u��N�ni����'�ۓz\��P�t��9��@�m���5��9��~3�$W�헛�Uq�ڧ��N(yh��=��]��Q4��D�Xz�ݭ��D�V��5G7sݎ�}bt-�t$�������V�r�8/J͓\�rF����#V#��Q�jP�������4���F�o{��P��hN�$�lJO�R�F�+��Jfs`��ϒ9
��٫��S,]������_��pI:l�'(Q֭�S�v}��h:Cz���?����� �;�����K�
2j�ɹ�V���!b�N��n[�)g��V^ض�g��]�`�i� � �՚�O>]=��7Y���0�+¹����`�KFغ��=�ظ�L�x�,�MOWbbB�9]�J�D�e��1Tǻ:r��܋��M�h�G����D�fs��Q��)OR�]|!V�m�=�6���)=6\[���pV��zJ�Y��E�
��3{�<F�'����2��q��u���Xp �'���)���eM�,��j��n��YcҚ�k���r�G��G늀{���o�x��<��v�c�j�3�%���y�q.��~��{��Rp�0�d�.�{7�����=�H���2-��os'���ln��{��dg��	�l��;�5��}�x�߫�k]y�2
�Q�S�������U��,�s5�����W�ۀZ�7�KvY�.�|�w�������'
�|~}�G�����A��c�zMr��m�q��e��p�j��h��7r�ޫ�Id�*�5�|��@���?~ߡ�׳���<9i�;d/V� �]�+��D۳H]�T��������}�W�����K�+���{w3���3}������|2=9{���¾��Ý��Uv5��/E��C�Se�DI<��I&"�θ������{W�Mt/�sFONo�kY�e-�H���n`�W8�Q�^����D��=3-u�f��eaK/	r��P̾������Й��Ha%��#y�=J�f��0��(���^S3��<�����x��j�:�T���//&Dߕ���~��&v37΄��|��x\̙��=%����) ��γ%I�j��e(�S�ї�Yo�]\:݊���(Y��S.�+�����f����y�dݿ]9(oy&fҁ�
;�!_l	��$`��[H"��Tgh^��u[�ٮ�fw��=��X���S�,cx��g���ߏ[�=ri�R3{ۚ���kl`�M6����g8�E[�i�HZ���s�N�*η����E�)3sEU�>J^]�wl�
ֆ���{�}f �b @E"�9�u��Z�%v�ey+�-碎;k���ۛu������~~��	��/Y?	��5��ȹ=ޮx�N/�"�K�9�f!93,�z��ˋQ��n��}�ˬdC�bFm�`r�w�r�y���e_t{�������u|�$]
X�=m���>A�e��V7�����Ë�[�		~>8���h[���w	2��я3P����}�rإ�����]�Z�^�-�}ﳯ�����p?�?O`��z�i�FƐ�!�^���	�=(�i��z��	j&W�#N�y�主��$��@ǱG�*�EQ�U��۶���h��~�� �3�y�43����>%`b����z3�x��E6YP*3q/f��;j'�&�'���yت�p�g@؞�} ���M��B�]A�����wN9����x�e��qE�f��&�o�f�5ح�؎�!�! !��	�����y1�M/p����Fj[��.�N�^w_���R �[Ύ�̪ⲑ���{��[φ=�ʾ�;M��w�$�J��@�C`��p�����Ưn�yoT�y$9��Ec��r�:��`�0a�P҃�.x.3�g�<�y{c*mÃ���f�t��{\�d-�{�˙�j-t�I�Pq���Eu�[�ѩt�$��Nn|�q���t{��wϯo��c�b����}v`I�ݱ̀�m��-$��>fΧ�����\}Ƿ�i��[��A��֞�}�����aA�0a\��':���,}@1zvA���V0������_()�a�5rw@��|�nEws��D����H���:�A�f�φހ�T̐R��[�ݻ�5����aȘ� ��U�\�I���Oa��c)�=#��Vj胏�«�F�n������Y"u�
zI-�t��J�d1YqK��ؘy�
�,�N�fK,^��lGh[��yǳ\=�،8�`�|S2X�ũ#����u'7b�|�t�Ӡ�N�J�z"�q�6AY�n�j�l��ܙ�V'J�쬦*M \��S�ͺF���+f��khS���d��*#4�7��2�V-�/Um;|M=���]h�4�Qa��Մ �����A�XU��C�����g@�Ɂ������`ten���\�4袟�Y� ͻ,6�d�pv��6^;pr"�u���@�cqX
l�Iގ������k�z���鎮�X�m��6��.BH郷o�N�/n9%��F��پ=}��#:L����J��[Q�s;��)��1���"���i��Sse������U��Sm���L���_u��� �&i�����-�Ş��O'��L�"V�8���{�>���H]Qm}�3w�	���%�:�*B^�_IuX��eQ�WS��z[��]{����-䚚�,@��ۖ��I���_u�ot��b�Ͷ�
�*n`�����V���s��C�7y�;�IV��X��/�-m�h#sTRl��V��/[�Q��U�[���s6Ľ�٣���=��a�J)��Yۆ�2^:����2`�P��A����'�N�y�TF,�z�Qq�d�ó�'=�EvߒѼdd]�y���h1ԗ��sçr&����|y %�\a�7��J�n\�2a]f�RX���g����#}�ˌ͔c�'�\@���!��w,S5{�'o�H0���B��n)~���x_H1�~Q�4�����:���ɸL����G�����c�{���w��{ݻMA�#u� �@�Y8y���4o�^�K��I ԫ������Hd#N _Μ���;�P��[�S�1��l����<���s�C����pi5	��H��ȉ+���+3-�>�q#��R���:��@(�4�Nn8�yv@Cn:��g����y.qՊ �م�On}�a!���/2*K �7';yf�c� ��
st����9�饞����HQ F��ǠǍxZ��"��j\�e�l&�����4��i,��x7�;��D�xm����Q\͸���*�E{��Ce?����n�i�r;6f�S���X�pA���MX�>f N��+�d�h�D�����(C%���{M��	�;Ф��דf@�wǔ
��>OПi���U=��5�H��u*����t�S�*���7fb�D���al����������ݚ��$y�� 
�		&�1}@AI�G�`��˻}�{��@��ۃӘvmdc�}&�ޔgM��u����[����.�[�wY�Pi�2�����m-���:R1�*���������i�{���R���N�7�k���S���h�F�����tu�3�	v�F��,w,(�f�=�֔:���-/=�\�����[t�7K�|��#�c���3�+A�*jn�t8)�ûk�z{�۫81+��.v�Wn���_}�
��uq��^*�e����9��u���с�s�<���Cۡ8�$��5�Bu��a8����ny���<v^,�ʧ�{�b����pv�{0���e��H�N
�y~����	�*�k?"g�/j䙞ɛ���"Ae>��K�{�A�LA_"D�ƒڛR�.��� p;�^8+$! tĳ��Q��y8PQX��x�c�3�	��۬��!�6����YYj���Mw�"�-O�ӏ&%�PVHF�^�4sv;�m����� VuL�^<��ސ+x��k�V(�oq��r@ Ƹ-��R{p6��6�Ǭ�K��<��cu��xŸ�u��H�;�;�wT�)2�Ұ���4�w�}�C}�K9�lxVT�Jvϝ��z�'!����^��r�{a\��N+�4��t$+��
2�(��l�k��.Űn�"GW���'ދ��ʍ��=	+ۧ��2�:�M)J�E��Dd�Ζk�kQ�j��#fYyG�M���9�[�K� �7�#���ܣk�}=�'��]�FdQ^��uL̏���5|�ڗ�1)��̸�04�^���>陊L���h�B��vuv/g���1�,9��[���>��Z���Ԭwx.�2xj��?���w;�M@+ۼ�������"�1�)����x��xl�p���JΆ��)9�����^p�Ax����"�Z>��P�M�o�5祱�~^{["�q��eY���|�ɺK%�P���~��޹����#3�B�=�JZ�_��Z�K!��:�:\�\���.��f��WMv�p$�����q�3;*4�M���}}Y!nugf�o���}��֝�u�i��{I���������E�)��!�g��3�	�u��N�B�6P�:ig���i0!��{��v���`�^:�Ť�3n���fLr���`����w^!������E�	91������ݼ!�V���^���^���7r�����
�n��=�m��';!U����0����E�lW����`�*�#B�H~\F{S��k�+?�E;�X��&��ia�Gr�XP�V2y'ݪ��}nNT�۸�B��7�Yv���8�@H8m��A�HjkR�
�ۓ��ov�~��M9�a�Z�cb�<�7�s�:>p��O��S�ܙ��[�-Yx&�E��[���ެ9ٹm�}��E�k�UT���JOfh �9&�8s�����$���fgח�'g:d���v�.l��*�O]˩����]��%��=F%Hj0!��ʇ<�بq�5p��-T��=�)ܜ��1��}TPQ1�3�OQ��Q���jd���o ��㈬2��6�|5`��<��.�;x����3�Q���.8N�t�N��)�{�Vf.&�p�|\W�wƇ�w]z���V�Ka	p�D8�P�%�|&e;&��|7o�^v�/ m;���;f���a�Y�ܑs�n@�F�ʨ���Z��4񰚻���0.MC�w���GvqS�u�]/{�o�_Zz�׋W���n&2�
���w��vE�hP�(��(��fN��㍋�.L�]9Y�#���\���k�L]�1�;A��� ��⽆�l�Ly�p���ԍ�à(�0C��/=����r�\l]G�'%뭳{k���l!M/v<��W{}���ŞV*d\ͳ�cѵ|����"����3��S��bc��%n��k� ��S�^oz�E�֙��gh�������:��PA2�L��ogU^�fwDu˳�;.�֝tAs1���2����N@����L��6
�����@�w����5�� p�1��}�&���&;��$YE��ŕ�7ޜ��3�T��\�5���#�L�؅!��*/���zĮ�'>�N�j<�L�6�L+�س�T^���\i:ک=>����`�؀�X�}��ku�ٵ�'�*M�c�����UL�>.<�R/��
smJ������!g��͛/�<�V )I�q�l{��"UMv��&�Q��~�+VT�O��ߎs��6�!��Ou�l��\��3Q�xp�I)k�u�!�������( 8�s��8$��Dڻ>�y0�!�X�Y�a6�P �'#v����V�����S<�I����� �Ù�9U�*�濺O��v,�HsY����ܧ��FF���^����P F�0�d$Ae������,�'�?�ȉ(�.-$�Y�t�F��	�Y;���9:��G����z6�=
=M_q	�\��G/ALW��T`��~�D�a��5�=��:%��i�Ɍ	{�'=�<uD��nH&��4#^t�:%%�\�i(r���*���/��3i�w��Af.��t,�U�b��c+iU�f⌻��j�����oBq]�/f��G��+}ڂ��=�rru\/f=m@i`�/],�0�:y����||.��/jg*�k:��q�|��RE��(E�ēbb,c�+g2������^^mM�}5�&�drUu��X�;�xˋ]�
b{��$Q��-c�Us�U5iV*�����}䠙S��t�wt 9��̲��HU�lq�;7gv$�4~g��M>(]�Z��T���B���W'����z��b�_̼�AQ:�4�D�oI�,B�o��Q䎼��鼽�}=3g��g���̝���,Mou�e44�%�.s��Iv��c��wE�|����Ǭ���s]V�H�&�n��S��A3u�0ֻ]&�cm8C���p!�N	e�RB�b$��'�w�֦b����~�k,�t�:�g�zqT�(�IH���c�H��+�=˹�K�w��+X�cyD�L6��߂�	d����Oq���B��6��sL��ۼ��3�ـ=�q������r��x}�CkI�a�iv�sٖݯ�Tђz��;S9}�P�=�z9�!��$�>ģB�.�F�=��z���F���$�x��G�:�=P�'��jX�P�Fo&4�[��o��q�[���^	���M���V�J�{j�����-�c�tlp�
l��paׂeg|t{��[�����kN�2H��\�4��z�^ĺ��L:�P�O%'7L��5��7�ǈ&�]72�.��u�ed��S����=_0qQ�R�ao�cm�%�?�S��^^t�{cR\�眖[����s�����c�8�\�̃��a܁�nzvgy�pmѠv�͉�C�RpM�y.9�osדoCU�;��5=��}�ڗ2E]'�v���j�vl��k��υ�2mP���s���qɸ��1��Z�a둞̄aʺ�U��cH=:��.�\s�e�u��Q�Վ<#�J��=�ĻL.���zT��$�,�&n��H��*V�ߎW� ���;K\��"�}7� ��&�k�n��4t�c�LR�=�=��J$����a�v�_Ob��R�p���L2�}��CF�b���(�v^>��0�b~��О��d���Â~����I�Nƚ�=�L:=Jk�U]��	�alZV�.��/ r�6��$��!�Jn��~Yy�n���r������WVn��{�?�]�Fcn��q����.�7�3��u�v��÷��H�1�wi��Ʉ#I���hh�����(}9��#A��:E5�i~%�"3fx�#eB��mt��u�n���T6��U�ĩ�dˆ;L?n���S`"�qC-�M�ᜬ��
�r9�U�X������pfs~�b}��_M���m����C�T���������ar,��:oē^&�2���~Q�k�_ԝ)�4қ��e��~��V8@�6B^�� ��{یNط��;2��3�޴��gW�ʫ_I9#�D��t��si��Ji5�˗��U�3�Ǖ�s�9�Nɹ�uM�X�Ut���r��Z7;}�04��.~;p�W����KҜMvm^Ow�p�7�j!U=�.^�j(�� �$�۴G���_�a���rv��8�r{�цO���y��r�&����;��V5π��B1�\����_�����������5X� ��f�Վ5�	&��e��1�ࣵe^��j�&���3]2��&�l�mR	�9�h����Y}�S]2�e�o&��)��n�VϹq@�6�P ���{�=J��mm�����u��9��[n�)�glM.�h"v,C	@��I4W�qc�ѧP͹���jx(�:嘳n��+��=�~hg?s�2FY:�l���3�{�����
�P�G������o�㜇.�e�Ps�/+v+o{����	0�("CB����V���,N��)�� P�DQ:���uW�:����m�x��D�Oɓ ^�����Dm'�"V���OO}$�xwa,<�%��������h��B��fzn9��NsM��&��`̝$/VwI��K 1(�w}xUqWFrn����@|������N&R{r�`����s�P��m�]�b8~�o3���ڛ�to��@��eCS�=�=����o���v�z	;շe��3/�n� f�=�����N;exN�]Wi��ꗲ�Wޮ��7�Wkz�}���w�rd��E�
�8�����r��W�F"M������,X:�i�J���vcun���_�ޯM�3f�jڨB���d���!�;.�6�[���Hć���컽47t�\�2�h�7���RI��皀'��2N<W�ߏ��;��ֻK��g�N��K g�[�Jz���������.(0c2$���xdZ�^�L��Dڹ�sS�e�mmқ�.�Y=����%Z������`���d���v�e*��4�.̛�.h�
Q۷�G:�8�̬�Z��6���cs�I�;���':ù�kyv����*/7Bh�n�c���Eu2?&�i��P6�ٱ� S���{�7%���Ї�ȣG�\��[�ٓ�5�CF�i�l�>�c(�B�t!�O��v��>���i�T0�_Mc_/�Vz]�w��y�^��(W��S�?jP
����kr�B��3��{��m�Ώ�>�W��C�a�:���9�I"�f�w� �1ɱ	��V���lk���y�N�wct!�=R*V����s~/8n�e����ᠫ���q���p�)�M�l���#p��n��u ���yjօk��^=����sm��m�_��;yz�;��20`oހ'��>����vx�-%B3y����׮�%MĎ�ϖ�lf��\�5��*�WX�p5N� ��Q��;��EZ�W95���ٹ��bV�GBQȷG�〰6�%O_W]�<���D&�?��5�I��i�g���u4%�l�-���+v�=4����Ó�s�D�os�2�1h3y̟�ŗHO!�4V�-n�<�mGhp�Дa3�<<�d�Sc3�{15��Г�%8)$[7V��)��¾'��.{V>�(c�h�#*��M�0AjTa����Ν�51��+k}?*��~ Y�GI�Ce�]�D��������L�!�V���W�
��fF��$��h�@[��ꇰ������1�_#�3{�򛿡���2�̲���g;f�':Mپ�4�Y$E�*�.�N$f��EV��e%�����UT��(ḙ��!�8h���Nh���k�r�%.τ&w�r`݄uhxy}!`���+h������}��GK�dǷ}yJ�qtHC��j	N�^�C�DC��T���	6
�	�&e�b!u�#��ﯮ3JԾ;��ӛ~�y-�V���#���C;;�`ܪÊ����]�x�w�h@�P}�Cy[��&�c�bB�@u�6`dہ۫6L��=�^��2!d�wTM}�u�xN�lΓ��+
�`� Z́�5����2*t����]T��1��;>��h���&=W�0�_����y����e���m4�*zP�ɭ�^f�\N۟P�J������G8v\'g>��@oI� �S�ٰ �����#��C��g�ﻔɓ���a� �?Vg�ߨ*W��e[bܮ;-?V�n�}��|f�][������T�ew558��󭞎(���~CM�:v'��$�\5|�'��瞹��|�Y�٩�����/��պ�{��2]�j,��xN�Ws�Tg(��]'e)�����8�~hF���VT*�WO�1ϔ�����7��g>��/��AÆ�mtg��=~_fV0N���g���[��>��e������ݽv���^Eo>��y��Cě����龏�ٙD����u�<0Fi��1�W#%��p�w�!�C��e(-q� �x�.57U���%�TH����A����<��!q4v|��ue�=���㣜�+:�w�Z�u��K��d�w��p�^_^�Bqw������:�M�Un6�P�#��o��J�k.y��8��Z-u͝�u�W9O.C-��pnn�o \Y�{R�7��Nr�3��@׆�u%>5�ݸ�/�o��y��p�K�_h����ln%���8�Q���bZ��q(A�\���x�����׷U��ɞ#n1�8ێ�j�������q�)xv9ٔ�;r ��m�g�|��]�]]@�J9�*4���ӎ0�9s��x��0�#�$��i4c��H�(G����c���z��Ƌߘ�;s:�\�>%����u4׻�t�!�	h'Pz*�{�{�x���|1
��L�J~�2�%YF�vl�99ǲ���}�[gַ<�;��j���1��26.w�T��/|��ʬ>�z(Ɵc��rP�$M�O�;���8&�a6A(�qD�����H�ǲkkw�-��/ޡ�d�U���`���u����t��lc����I��s�C۞�r%�
i��9��������l� �gB��������x��Z.?��K
�n4Mz�ͤv��_e�dxL��=]���CcO(�a$Z�$L��=;��m+�Y�>K|��m�]�3yp�F����v1��V?wER���+8���������$�P�
u�Q Q���AЇ$�D�����Xr�*�3�w.�ݢ��p<&�3L�/�wl#��{��U%D�|�:�VZ��&ˁ��׏��a����R:T�f�(i:L�g��75��&Zl2�-8�#��}kx����a���m��2��{'ʁ0__�e��d`��)a��^��ګ�/��"W˛�<�	�Z�V9⨌�<@�1Sٔ�V�<�$Y	2�pM�Яk�=+4�}ep��۠��t�*�۞�m}���zb,r�	�b��~:�:���M� �c�D���~�����ϵ,%bX�����r�x�O��.�8�|�fb}�@�G%2.a��5�}y"���S���4�A�6�Us�2t���NZ�啷C,���O3n�QMژp�+l���=�T���Q�w�X-�ڃF~3�$;�^�����8RNR��R��ݮ�'x	��_^�4L�Fu�Z;0�r�w����5�%�6E:��6K]�r�bm�۬p���]u�؞<쀔�Y9��}��@�8#+��܄��z#�Ox����ېѾ݊�${ +���w���_ܿ9�w)�P:�Ea�dU��Gw��§v�sU�EBV���iWT)��Z���Qs˭˱ն�".:mFe�msC�&�s�n�3�qR7w��U��b�*�Ν�X7�X����)	�����jQ��fQ����U�n!ۼ)eN�e��kqв2RY-O�enc���'{�s7�I&��BN�+DyKN��VV:���{3��������K�@�=zIs;y,�kB�֡�LU5P�E�!�S�Zt��O��aw�H��2�'d_��k@x[p\�rf�e��Ym�}�S�;��9���N��ڽ�E�b��[�]��p3�]X�#��{t!�E��M�B�\��[��CP:3�f�vN;չ\�R��RYsv�.�l
ѽ� k��c�F-@�̛�T���y�]�t�EeA-Η�ݹ����滭#g������j�%U�uW!0*���7g6��hm�)Uvh+�BS�W�k��nTT�:�0T���ی�u`6��cm�W�7���.�F-�l�5���:�(Gl7WV;\���,;��\���l������÷�B���1�mz3������
��{F|�z[��vpq�i��Os��=II����9�5�'W[9���V�ۀ��'
5�� �p�ny�Ɠ6�d�^�f�A�ӝ�<�9��#���c��70�ݣ��O*�鶗k������k��=� q�ۓ��݇�����6�뤮����9�����]!�q���Y�7��<g��f|�W-���ʸ'���p�,�=�y:���N��{�C��&��n\];<Cp��r��=v�_k�}3�uʘ�;��8��Z�ٯ9c��]����{n�rp���k[�&�r����t�ȼk8�:=�lX;<��L�>�ncq;�y���X )��cv�f�]�.��`Y�t�k��f%��^��W���xkh$u�#���4u�q�m�lonÄ8���2/[������޺�N`^ݍ�k^s���3���k��LDj���M��w+'0�������{H[�kS�n��ݎUK 	s���F]��%���5ծ9�]�8�p	JF��Շ)������0k�zxPݼݛ���r.�r���q�l���(�C��嘟nm���NLq�D�8�̸��c2Syz���<�Du�yz1�������ɳ�n��
i1�(N��Yw;��8��yFM�vʕ�<j�ݺ(4.�p��v���^��]���2���Qѹԝ�������\(ǖ'�xN\]<Pb,���[M/4�\�,{F뎞b�{5���nXw U@�9��g�-��f����{!����j�.�y�nw �.n:^������A�N*5�����E#�Ӌ�wIB"��fz��$1�q ��6}���bF�?&a�ʇ�#����l��ٕ�3�'�g!�z�{{��"�-2�a�v9����1�Ho3�ƌ�;�P���7}OW���[�SH3@
���l�9�rq��N�� ꇜ��@�:���OOh���z����n<�i������A����O��k-	i�,E���.�y��K�@��Ί���d�h�����a�� D����R����M0�R���1Ol�cݽ5�2��w���䋛��[���5,������J6��@���bEK\�"��p�&*��z/�i��?q	�E�lE�(x�\�2&�
����5^xo�vU�|�\���H��x7W��ّ�#8�5v�f֫�߀�����i1Yu�Wӝ1f���F�~>��+�D���g7��F��c�I�,��[0gB!@���שP8<o�>\�6k2�/��c+n=q�8����i�z6�(ߐ~��WQ��V�y���ɇ�ZHb�Rח�����Kޯ����8P��:"O)�Ov{F�r�2�;:���.3L�Í�חi
�vk�(���T5I9lY]جJ	g�gb��������'���M�d n�C-��/G�<�ټ[R*�|:8F̨-�&���Uže`�sS�@gd6�yF�7���F�����e��z�x3�MX�A�h9�/�O]Z͝/sqyt�������Q��'!�˯Q�]R�
��i�v���u�q�b�C��fj�F�E����і��9��#�
k����93���fӾ���d(
�o8,(���r^>=�3,�U۝���E✻1�{S��������w{����=�rm�6�S���5{�2+��绗g'�=���G{�\�'DZ0p�o|2�Ʈk�l۽�i#�e*>�)���6wdSŝ�O�IL���?{�͘I�Zi5�|q+�"Gԉ�������Y!�X(���t5�kV����3��5�P;.|��~B0A���b��ւv�T����؅@�q�^��5V'L2�wge�;6< �f�����2�X�nK�r�����~-��p��#�#�8w�݈e^PYP>�&'$���$ƈ"N��Ef]�F���:�nP:�K��ϼ7+��,��oA@��J��S��s�F�ل�;�
(#ADC������Y��l����}���0̉���(�.I��*U�:7`d�m�5]ߩ�#�a���X�"�>���4F6��(Ƹ!�z��h��B] ��sx(k R6����
��mW���5B�p�.0UA�<��p�:�z��d+�J,q+�5��te��@���T7kx7f㳫����\h�;=rYۂ�xr7\��0P�5�{�շ4[�}/�I!�tc�UQ��쓎�wZɫ�L���,YO��U�T���2g?��$잟fq�2�dwˋ7À�"jI^�n����7.��C��_R2xuGg]�y˱�,Z�
�S�a�����=���2��,X:�D�;9����~�O�]?����(�f'ۺw�����:�R�\�3��iC�W�H1��PV�}.52�tYwr���]-t�?�^
?�~�d�X&��#����k�:�խ,���χ�|���z�R��w����ٹ���s�%��@6�Q��R�����qh7�;^x�5�zLZ9������z{����G�i�H-��!k�O�^١�t��qH����@�xe>{s��w�oڎoY��\_�4ǽ>�p�1A����R33�����+�F�Q]��{Cc��$�LA��Eɂݝ�T_E��v�C�ۣ(N[��n�������D�2�r���Lق�v�mzL	?Om�\�����䖫���?J�?��N<Tϻ&b�]� �.��%�D�/���>�8cTne��1.�O���-���';ʏ���I�Dm)5s�\��H;����~�tϙ�\�t�;��3�������	�o~�"�Jtr`f��vY�dfH���3�1k*���r${s��y�����ߓ�9�#ս�_=?v��� ���7r*;'�D\(}(�{�Ck�2l�^�Nϻ?v��^RH4�oz��v{D��&k��:S��~�am���	�D��Us���X�\��ECf8�|�e�UwϽ1�0�b
pZE����=��+T=�l��U��� ��JhHU�=s���xVyk?xj�1�niD4P�T��V��j:hE��PP�,Giy��:�?Ӊ;vr9a�Z� ���E?�U>��SM YU���ʦ{�gk��M7tC�%��>�Њ�BX\���C�诪�4�ǌ�>��NL��4r��\��aR>�Z)�z�͛妁�8�S�iKk�$�jh�F��um"�WS0ֈ�7_��2��  �������c%�����3ܝQs�s�g&֞x75��\!)q�z��c����]��r]���`9-���W	�?�����i��R���׎T�J�Gv7]�-�[�{[�E��)'q��a��Ю��K(c�L7�D���; �[t��/�N�S�A>��*���rp�e�v��˶qIM��oe�&5���I��?��="$A��������1㫫Є����}�R��sAY�e��L��R����ÿ�}���(��!7��w;�}�'��bg;;.��Z-:�2#���F��W^�,#�QkO�x����Bh����?c�~*h��=�#�c��ٟ�O��֢B���r�5��rBH���!?J,R�8�:�@}��W8ٔo�����[��_";h7a�j�D����k��C��w�8��V3	Bp[l���D_�}�o�N��ZXu*�5d)1��"5��~'}���o�/&5ܜ�<��ފG���7}�1"*o���2�0Kl%�٣���Ay��p��\c��q��ye�!+�s����:ڗ �� �\���Ҭ*�\�����k��L��6 �!H~��$��̕G=�{�p�L��'T�n!�e��Aٱ:̬;�O��;�
7�(
/F���wZ�L��%V�@q�^����Κ:H���2B�}jv�z�+dӝ�������))~A�݋ށ�Lqf*�Z������#N^c�t.�;%��ڤLz��ڻ�.�&)�wx)D��}��{75�@��3!���ۙ9�J9hb,�J0}�fw��{ ��B!�@�Q��~���q�h�[���M��
���s��ޗ�~Tj+�B��	t�=6���W�[q�0DEA4.ʩCQw\&�a�[63��A���>��sy�l��{Nԑ(�M�'`�}��6�p�^�G��<��*��Q�.�ƌ,��Hy����H̞�[�u-v�#I�#P�U�/�:����A�kr灌x�u:�����.fa!R�1�]93/��ž���E�7ZIx�:7H���������`!9�^���f	E��(�S[{*�kx�Xb�8�մ��6��I����e�_Q,b�J��_t\��?b�WU��7V*��0idh��\6�PS-g�(�%�?!_g�������TGڭ��ğ����s{&�1�t�	q0���++�	tǽ��BT��c#s�����L�s�?1 }�|�MBۇ�ٵr{�O.`"II?�I�E��ή��L:����7S�V8
k�3g
k�:_eG�A�G��Ϊo["-|��J���,șU�����
�#���י����
̉��G��H��od�y���&�2ܮ��ހ����e/ �@#���5�u~����߮g������ψXh��]>u{��`K�C��+Xf�;eѾ ��#V!{1�=�"R1n�ι����d%0�t`/����g�0h�V���#}�!�փ֩,|����8���#i�p��?h::������H�����O���)��]��Ζ-���7Ӵ�������%19��	R��}�lК,�!�����D���;�j�gA�DS���;�\�+���
h2/�,@JM!3>PqWu> {7$���˺ۂ땎�[�.y-��F+=��R.��=sY��>&<",��̌�h�^�q���v;s�$���>��?{���7�F7^�zr�5-x�ܘ�A�Z�6�����Uv����ͩ������=Vq��Y�h]ӭ'��o�<��%����U���m0eE%��DW/=ޭ���ʋ`�f�A]�h��M���ٛc7<n�/���e�H���f�R@Ў&'q��I���3�׳�l*՛��I9'�4J<�y��ԒqaD��l�>�	���vp$rp�E͈%���L#���,r�{=&{�	@V�"��"ܤ�{�n��#�������5M�ur盛��"&���f	��.�~��9�S-�jo-U�!Sk��������9�z!� �	�-X�P�o���Ț鄆����~���R7s4�/�J��vb�$���������H	�H�J5����c4ט����pp�*e�9�4o=���EBpm6������_{����
&�{Em��g�Ʊ�j��� �L)*����i�E%������<!�ٵ�qF �除�����m\kQ1&�b�b��j}�^j�3�D�)DUkܨ�^�ȣ���  IV�������n�)g�<i�=Ѵ/�'+�G�C�y�Y�[�EBP�S2�n����*c�{	�Ӭ��Ld�Nךn���={!�h��wT!$b4 ��\z�ˢ`�U����HA��6�;��+$�"�(�������dŎ�}J���������+�dЍV��|1�b�v4��mK�bYBnTɌ �ˮ\�#���B��>�3��+y�r�@���^���#J�#b�w���ӼZi�?0��w!f� ~�����7��͟�`��'��8>=�B,A��9Ү���5z/z+o��t2`�g�qS�KDn���Ԟ�33��C����������s�*oen_c����Z�d `7������{���v�||Ϭ�䪽˥T��P�?$(2:��cH��d�f��!S�"6���wsё��K�u�R��>ӒOIL���̻~�@� ���h'�T� �Qf#$�O3&�g�a��E֠͑䇄gg���CVج�rb�]ӿ{M�W���]\ԑB#uDY<>90��O^���#�~9�#A�򌓌����o��PT�$�ٛ��j3c,i����DœB�*����A�V��L�A�#��K�^F.J�h�G�����t�ƌq��RM�#��Ѵ���{�/�ӈR5�Z�3R�)1i���u�7�.`��h�E��XM/�T��H�����}v ��������F:�m����Z�GUn��V��|u�F�s�t	��8��'�m�ø��A_�q�~ף��nl�'f����p�dD�Ol��H}��G�`����\�uM�'a�b0���Aڮ1�1\*%�nT��*^����e�M��V`sP�V/\�bbr�`W( x!"�ϑ]޾j��{��{}ΛS[���N����ghr�V� �|������Pqy�#�Y���ެ�"#�=��/��Q��\6d��2M�D}��&�a��sBi�쟝q�Fg�����DG�ng���5�ÙM�<���L��J�1C��	e�����f&��a
`n]��Ύs���!#Ԃ��~���cѝ��Ĕ�A����!�zz[kYQ��o7v��4�7�KQ�C����qrk�K� i�WH{����;�aH���t/&�A3/��}��=��.�:�:LaU����lg)��(��3!e���;���F4R��:T[e|Y-��a�/\�v�9q�`�ls9��Z��7.pn,n���n��=����S�̖�2p�%�z86��ײ=f.َ�,�R���}m�M�Wg��U�����g����j���zt�m�������:�5�ɸ��s�a�pY2E��+;:���u�����s��-�\պ;a�#u��d7t�o\��;2��B 0�"���1B"���P�]���q�lZ�1��b+W��N,�f���,�ӫDk:���{w2������l$:��\Z(zc��=]�|~����Hb�WT*<)X_@V��g���t���A$��jRb]N�E뙩(R3�n�\���߆�������N��LE[��'�W�ë��W�9:pഃ�(F��I?$b�'��N�7!I��CY���=~F���3t|hп'-�8�N�.�J�st�T��a܋�[�e�y���!����s�D����T	]�Z1��V��S����{�N;��������o�3��b\`��L@H";*,w���c�T�
��0`� ��-�&Q?=C�>�M�y��H��0�Y�N8��ڊ����/V����'�ז?�P���v�o�h�L�."��=������ܶ��<L>#�g�d�g�&�o�Dy)��%��5�Rl~�pJ�`�{�M� 5�+8�#��P�������d��#�R� m����\�W�/��F��&~�������om`�!շ����C VN��#�h��I���M�hD�@��\̺�A3�C�A�#���Xvb3 ��{v&48G�3�!�V>�Ǹ��i1{���x�60j�z;3ʈ����O��|b5�	=���D��p:y� �a�$Ě&���w�m��G����? ����J�=Y���ZM�BU�S�+C��Ĭ���5shP"%��/���I�QoCtf��Ыo���ݫ���ݦ�봆j�%;���նݝ�GF��f��%�{��=��A��z¬$-�F�7� rE���� �A?T�6���֣�ᰃf1�������Ȇ���p�L�$C�z�viNn���O`�4�J���ۃ�?�vNiE:�h�),��vM��5�K-�@wV;��pD% -���
�n�Z�;�UH"�%���(0U�=W��P��Pg�d��(`�Y^�\j~���d�[���*�3*xצ���&�M@�I��-�t=���5R}�]+��?
��r?����(ӏ�)G�|G��S��@�F,DB/�\=�w2��&����#�\��	�M_U�V)SUʔ�|'�c��eF�Ȥ��6�,4�Xz�kQ��վ��A��W#p�b*�o�LL�]pVD1��B�nʊH��|��2��n�?vd�HP$ɮ����Xb5(R!	=ݷJ�����E���bw����x};�$E;�D�!�p���N�frcn2�f�7"t�-A}��&/'9*4Cg D۹�|���6u�/�	��?�n�$b�ēTHc����5qZ�0XALc���w;zl��m�-�PV�m�Mr����!���n��kOB#I��Oe�Xu"c�/��_D���зj���`�N�`���E��������D1�0{|f�AL�ڞ���~��Μڛ����CF���1��ɶa��0�4~ZeU�4��B�ĹGez:h���p��>@pbݶ3erx���Z�r�l�g�+�u��v�'��<Z'��Z�{�Z����O^����B3J�}�����u ڸfG��e_,�.�"���lj���z#����P�����.���c흴���w��ז���;�K��v:ݢy���@�#�Xx&���1
��CD�)�m��Y�n�����s�$�pIa�D=EF*
�FD��sQư<G�}v��gVVo�q,ƣ;����{��l���z��=#��/(��H�p윱�z6f=J�P�!C�EV�J��3c��|�(Kr��9�U	�³)���="٧�)�s轏���\�DUOI&��|5ᖈ.z�/���w5���|�b'}�&�����G4Gx�J\ ����3ي��;˒i��	�~�=�f�Ƶ�i��ӂ�|P:|jі���۳"��,�]7YB����3q�P�a)LD�#ZR��ӕ��g���l��WS�0�=sR��":��@:�ڨ�d�e���#w�,)S��hZ�W�\h��ϳڤV��r �p<���u���aQlU/_w���j'��n�1a7�j�� �>��uLF�Glw��j.�������e�Vfݱb4� ������i�����61����q�y^�2gp��{�*�Bp��!�Q��C�Jq�0��96��M4c�V�v{^�1%��<�*h��3 Fn��v��v���#$g�p�tP����]�Bbs�#�A�I��Ÿw	ɘ	˼�u�xz�m�0��=��<��[�8����:B4j�Ѩ(�'���t�����D�0E�b#	Ȥ �wg�I�e��f0޿3�aK����\��+��p
(ӂ�b�䠏֊��;�n��b;y�O6� ����ܗ$���n������m>I�;�T��M�8����3�n�׺�]���e�ƫ�a�Z%�鎍=X�Gى?�VU�J���m`©���Cv�Q1۾���[�_�nnY���E��|pи��ÊC�{��ko%�]��tR�H��c������C6�MA]��oSTh�\���Y�gGn<Ԓ�rP��k�;�ީ5����+r��W߬�γ�5��M/�X��lz���!4��	������;}��m=����y`%lkG`��r�����b�$��Zk�_[���1a�Ÿ�ܰ���̹��D����]�zȊ�5p�� 8X�N���/���)`�ͭ�ʏy�}tط�8� �e,ɹ��ݙs)ۛ���ՅbwT�U��EԺ�l�^�=����tof�K(��̅�}�Y�N�V������N�{rB:�p�80I�s8�D�M��w���Z;��[9t�J��:�Z����/R�:+*e!t�d2���VV���@zU�T�T͎�b¢�����A	���35�ѻw��>����C/ ��E���1Vk[Rs�)��չlI��A7���Y���e�8{~_F톞n�E�(d���3&�p2!��0>�H����˚ ��I�Q����8�l�����m	��=�ӷY^�Ī$|������=������K&����.�I��#��y�����&�8�6=is������2�2�m��1���iJ��C�禳+�":�V�I.H�v(I���6]��q�eT"8¡��ռ��H/�	�SL�P� �y����z+7qeSBp3�m��:�H�z�.-SY
�̌�tf��~��ե���y���ɉ*a�G����s��iHn1}Wt���(i��-�U�q3X���k��c���*���d�X-ƚS���(�4�"�������@ƃ��y�Q�g�+=wDЗ��썜��`>�w��wo��F�27�(d�ze3����u��-&CpT&�%)�Ԩ;��7*Z�����W�ݸB8x! ̺Y�i(�ކ^2�%{�����]�Lg���p ��w���3�&��,�8�Jf~�{������*|��w�_Oo���Ҍ�iŢ< �ia�ډ���t�`�/� 8w
9��m��tP�x�IÁ~@�5+��	�ݻ�"^3D�L��,�>�̮�#[{2����?]�����:W���W�׊/ɸ8!���9R��X�B̷TR}]�R�ǔqp)(p�u��_���=���״k3I�{��A�t	�N�HX��+���"��#�T��!� n����wŁn
8�zV�����=ln�����t�K� ��[UD=��<�a�d��!/[9�|�<�jLz�r�x-X�3�'�n`��u����**����]�jA��!J��c��[Έ���;0����L��J������:�:>�2�Gΰt��ˍrR�JSQ�'���) �h5A�L�8�y5���]N���4nzٸ��Ί�A�4I���\7���mTt���ۇ�ݲ���t�mÔູ�ɸ{4����<N1��g��r����Kn]� ZxC��=����}z�X���2AM�-sk��nx��'�j޷Vi���awY�A����pb��Szu2t��ܫ��]�u��������)GGMKk�&moozP�+�\�#����I ��}CW�_�a�W��U�έU^����搣I��TE�����ߙ�ku��;k-����y���-`.�m����`��k���[]�ى<���\i�ҳW���Æ����£zP1h�HǬ�l�]�5Y���!�I���"v`�<C��ˑ�{f��PT�����������sOnV99��u�F46��s�s��s:�E`�[�2���ō�}`��__9��TJ��tTP�E#w��y�ن(o���^kc'��!`߳�ъ%�W�ӗG}�x��E��Z���
ه�r�>��a�_�j�a����nE�!���z��r{��}�g6.�
� �DN-��H��+)/�%TgI�WV׶o@A4�p�V�8����Sz��G;[ е5	�LV�K�+'�Ue�w�%��gA���#�\z{K��k>���s$�/�Νʇ�k��Ɔ��R�p�(.knS=S��*�Grd��I�Y�c��!a����{�!���6sHM�*O�s��s@����䶼�8����^�_��S��!##({/2��"!�F,AL�#zS姩
�DPc�%D(��fvf<ϣc��$`��&G��0VM�<�9p����s��%*l#'�(��=n[�Eult�\�>j���(A�d/�J��䀲~W�����K�4�.�b!BҵI�����O"/��M,RZJ~VC�3.-cM�{��%���9�%�.G�_@�K߸j��\�<�>�@l���^��0�o2ج��6T� �x���F�P̚��������L�f0�5��<�w����\i98�m��g�=�CU��V��Ф�XD6Hi�P�A��ɂ;s7���N�G��T�+LN�;���u���杞U��[T���dq��vxg�E��RW�u(+���a6ɲ;�4�� �Mݖ�*�^o��*x��|��u���F�5r΢���9E��rJAٕ��֧K@���WZ�_x�=<˟3�1(.L��]���fm"ʆ,*H�Y�G����t�'���ϔ�Z�iB�z���F]ˋ>��u�Ñw;}��*̅����Sm�;�Q�~�䓆��x��(�5��h,��&�`�T�JL����>��Cd��诧��=1�;4ڳ�:͛Hi�� C���(4/!X��j�禯f�%,���gv���̞ϊLU/2��ە������C�-�u�U��bR�W�y}�� �%�u����(����NgL�ks5ǣ��j#�43���{��ã��3�bA��])��-vͥ��yA���P�`�ʄ�D\�����$�rf��(8�$�{����K6���H�v�r��:�"5��1@SB�h|d5a�Ϟ��Z�q�+X������\�[u}}��_���p���S�C4~k��^Չ�!�{�F�nL+:�Ge�hG�����d��|ٙ�]��E�a��NM�g�_)Suov.�4�e&{Z��J�*��Juu��b�.hpq�a��`���(�O�a�`��~�V��4t8L��m���Y�<{Ռ]Iח���!xb[}�m��Ie�la�ͳ����"��.<�	�����ኮ�.�	�&G�BԢ�b?�ᾜً��r��"8p���9M��-��n����i�ج�@�q��	A��y~v��}Z�����6�Q�I�^'���z��N{��(�ev�q�g�G�q�+�C�ܶ624���@�6�����������H|���X��郗5����W�6�;ʩ��k$|64�-�޷�L{���#���L��}����k5��������9~�C�oh1�.�XN�n��������}��Ѳ���P,ш�L�B������xA�uX�X�]ܲX�3γ|�G�b�5ȯ_
�ݫ{hV*�{B�F�ە�}����3\k��G|*,��#�{�q6O;W[��z���=��Do�n��B���9���×%z=Jv1v:wl��M�D�8̇d>@�F'�Zkpm���y�pa����2 ����B�z[�B��������k� "0��[L�H����Vhg��!r �L�AO��f�
�q
sUGx�6@B�B-���36�찤X1G%����̉��1��� (�d�P��,8�ʷ^�5���'��U�r"�N��p�l$��\��!�!+�
ٗwAl}�<{Ӓ�'��h�5I�,]a4g������zT��d��E�Q�ȕ��N�cCpH�}Wu���-�+MAo��܌���T�o���rѠ@nn��Of�b�WS��F��M|�Lw���')`+ƒ `N�մ��s�X��ƻm��B��
����\�9�69  �`|҇�>"��t��s{�R�Z�%���YFn����3� �;�Kp�]�����F[���5Ϊ�z�	ͩ�"������r�M	CA��mNZ����tlIP�`&��AϻaA���N=�8���s��IA�T�$b�1�9�vC���j�� d���u[�v��#Q��y7��=;��iHrOzU�]�5�~�w����}��I"�BK%�(����x�&�(
�a��\�W���`A��6�(u�j�����f���u#������t'ۖ{�� G�uVd�f�]�r~R0��p����7J�b CD/_����Tc	��əW�;е����v�;��96\& &�;L"xc>�D�TovU���p�s��>��5���kۉ{i�b ��O�d�x�li>�����z�����UvZ�h���u\��`��;��&)��S���ˀlBL��V:��1}{�ے쥳�&:��خs�>r���+����b�/���u�A�h��� |V�͖��s�*��jDV��,�g����vx�^>��H�SA�Y�E��9N�F�#W��)^��R�ɕ������ͥe��y9<QT6���qk�N��s�N��$��?��O����[]\�,��c�)� ��R��]w+t�p��g�|9�畭/}��uv�%stlD�R��f������y8	c&�M���\�I7������7���<�����x�M/-�ev[z<�]Cv�A��{v�'`��k\�:'�o<v�sq��s��ԓX��E�oAǷVݎ���V\n�I��;:�^l�p���l���[�Op���^C\d[�ۮخ��n^�/��F������P��<C�;�bx(w�=�B�X@��F ���#k�����bn��� �s��,u�"���I��X�2��T���t+�Z`y�S�#�	�X�
#1
	��@�w�Q�n<�)5�הo됏_}|��>R��{����Z���+9��G�Ja�b�'��BF���Ę��0�0���=��'�1���ʨ�H�#E��23s�e��t\���} c��\q��-òhXV�l��ˆ�Ȑ�����0:h�����1H�w�F�=�}��iYR�l�5�J+�����gTXB>ǇՌyy��w�鳣c�A��(&�����R�����S-hҔ�Ԝ���������rWD}h���5(�'H�j�+iA�@B	Bj��� �ޞ��@��
��m��{z�N�=ɔ$� *��-+5{.��LT�}��/���_nR��e���T-�B4v�����l�&1𪺹>)c(Q�~�=ْ�+���7�{�J�B���!�nb��k�O��`�2����ņ�oM���'n�x�60ד� �aG�w�R1mr��3�q���)���4a�U;�3{X[�.�9�9��u��z�H�P�^$l�ud���\>G���H�:f������S��w�s#͗�x�ΚdrQ�+f�����'�hרz\6i.��P��/~��h V^�V8וk�c9���ѷḯD��������Oz��Cd�Wz1���$�F�L������x��o���V2�P�,�	�Q�M��ջ^ A�+��a�m���x8I��3
��PY���+��E��@)�lQ<}*���@����p\���i�m!nxܠ[���c\�^���h�� �G3�g��m��"�ԋI%r�Da=�^����7�x��Q�+��(L�ۻH�<	-,�w�{�Iy���v�=�2V����P�aA�}(",�?$�Y�L ���,����Tە[w���:/&gh �_��@�!��?����KվҨK|�bZ�*��(���0�D���{�d?tt�iBL��]}�ƣ��9�M<ܺ�v!����q�'ݨ�>yeЋ~��`�� ����Tk��4~�8a#���g ���(��zlU�Z�D�;��e�M;���Q�wt8M��N� C��3C��U��]j�u�J#���dx��b���n`Pv�l0 ���ټ��Q�Þ�y�W��b>����J�L[�s�����r6l��7r ����p����r���h����C���K�#����j~�ƩŔi�y:Nk5-��{�A����I�_e֙�Ǉ;9o(�#�e+6M�v�zO1�����O�9Ã��h��Q���^kL�Mb�Q63s+�ڊ�?O1�rk	d�l.��{��>nv������[kai�Y��Cm�J)�W�����u���z}��c
Ϡb;�(%�JO]w\@���Ì�;����{�+Y��к�j?�f��wkʛL�4A�o��.�/��F�%�T����=}�h�����	������"��J�0Ia����g?a�nn&����#0���}6�<���"	�ٺ�4U�����jOtf�y*�p ���Jzvy�S��<�w����ǷyK���gd^����	�SP�#���A�os.���7/M�
'M����u_��ҳ)ǆ�K���L4�<�F��(;fߑ�a:�T"��ώ�{��ua[��D�vwҢyuUE��p1и��jm�	�,��3S�:�dY�N���Z<L�7=]�1�/�˸t
*潹�
����#�g*�#���vt'D�{5�m��0��zΊ�^[[��Re8L������l;�)AB}�w^�6ߵ�<�_�r�9Y�������}��Iؿc/;p�v�x�*�	J�k����)��OOR�eW�����aP���g���q�M�(p����7)YLf��$uI�c!���(���]�GA�.Y��jc��μ�7�prq����������fIŅ�_	F7*a����{�:w-e'+�'N��+�6&�pLq?o�3�G'J�35�z�}�~�\�M6��.'�TneVĂ!rX�5��D�髧�`\�]0~���;K���Q^�j�O�Z݅+�v�y|�u�0������|���쳙��	!��Dа�!��j�ß�uK���_�9Z9i>�9��ܬ�+�'gN,w^`)��kՖe����z=��nZ�"0h��w����9��L�3s6;��v���ַ�fT�%��(��첪�K�[_#<��ok���d�Rw�Y���Ӄݟ �N����g�I�d�n����R%� �!è�x�F�a��gr���OL�wn�~��lc�<uP�
��Lo���ߝ�o�s ���SY<�w&�r�t�LU�3 �bb�O�,���IN(6 )�{�nvz摯D��6To^e�7"�^J�e��1���hv��r��٩m]B�~v�|]�D��=��2i���h#����b
�u�F_���sh��t�,��ɩ�˫�]��KN� ��t�|Y���E6T �`�K���n2^R8	��7m���ɖ�/6'�4M����__���ڴp��?,;������)\� E��������8N�w���c#�w7m��+3j��f�-�:�\9f��3�<Z�gnNW�9q�]��NN���-;��Ai���C!Ǧ|1�&9ր}��KF�n=q����Dn�U�c�]��F�
 @��6���g;�� �Xa&t
��Q9Ȭ�f�i�n��dT�(�A�|�x�)�v�t)(��/W�[�Ni��ha~h�F�/ufc���6�^0�9Ɍ0"zӵ.hT!�W�N�e�;��H��L�M���� q��]f�ن�>#���q�]�����^g�}��y�oG� ��˝8�⯻yYY�
y��P�0�3{\/Nհ9��U��ɠQ[�.�q���Ú�̺$}k7zե>H�@SD�#pƒxN��>]n���D���+
d狓I츤npD8�zx�y*�օ�+0v��n6�\���\j��11u�f;]a��GM��78������q�@�s��vۛnӧ�8Z�K�lr�pp��l��q����GF�G����p=��Z�q�x�N�Q�OF�#w\��15g���ۅx����A�n��������I����k j�rP8����s�2==棄RW��ʺ~z���y� 2��85*`��L�u��{Л�<i��+�HyB&�יt-ܬ��w��9r=����똑� ��h�X���k5QK��e�7t�/�YSםrF�z8Qj�K��t����yý�+ߵ�L�ȫG�r;�;�Kh�@��H��O��6uh��y��n˲�\0��dg�ªG&�Ru��:�����|��r�b �4ȉ��I����b�\��*D��߰�׸)�ѣ���@7��`{ќ�qޝ���xq<��_�Z&��[q7,'u��n�n���^������m\�Pm5��sD��J�|��ڷ��Ks�G"F@C�C���Ψgܔ
�	JE��v\�dϼ���$�p�Æ� �|�1`��rsn����ؒ��
6��H`�^��پ7�@J$� n��ΌK���tAȨ���>�N����g���_@:���=�*��t`+���
�A�����[��?Z��ܥS�1��0DG��흳�i�P�1��{��f.�v��w�� �{ӗ��h�1J��A���V�ƽ��$����Z>9�)�uP�38�qP
�o�lG��VId��XhBE@�Ny9|k<&aOA`D���S��b�h��АR�)��b�ó6,��/�]fF��6����
m=���"S-���28�������}\q���K$�z��T�f����ewl��}Y)ⳛ�q����e��ŀ��[��l���K&)mP�x�N�/�5�Jc8m�
���]ű�+;��p��	��9���<5V���Y:�IWE��7GU�r��0�t�Z��;xͣ��vw��5�El�4,Z"��Xr9f��O�c�Ld�
���z@},{�-�jcd��0'bU�` 6�E2�&`OZ;\����.ͮ�̛���tV��ŗ���
,�і��q�{o]�ܥ�Ql�TWs1�#-�$��|��V�Xd����]��Kd�-��k�u�]]E�:�_=�Z7�&j[@e��g+�^��ͧw��$D�$^��N���Qy�������׻��d�W��{�b����z�U֚P��݈��!J��]Wؖ��]0+2�P�r��N��I%�z�V�KY�oy�ŭ�&�j��C�����%�k�����a[�Gj���w;�����"��B���ezr��+�p���d�b����i�dv�9�?��: +}�K!������U��Ѧ���l7k_c6�ݝqm��/����������CE[��u?�ׇ�dmu�e�"|Wrt�Y��8�]��-\���@�vb���n�]���;��x�u��� ��w�Y��!��ssU�
M�4�Y�3�M*�_�o�{��-����7(ԫǘʠ�AwF��%��';��m�tљ���N�P*�Sfv

��r����8J���nl�U*�W	q�+��0��Z��&�����bϏ�aO��f9�8�:Nʼ���4�ι�wn<C�msyך���W3tU�.+s�+��ɞ�6nz}p�.60[�{�5]q��!wc�s 6خ�\�vy@(�Gv��nk�<WE=�j�v^�؛4�\upg���F�EU�N���p;��}u<�9麳�����ͻqk����7#�V��hܤ\�ꄻ�6ۇX��O�xp�ժ�n0/^{/N��RH"�Ѱn��w�������nydTkt����q��^���r�f��ZP7=Mv�	�q����NC���d^؞�J�m�<��E�ۍ�@xa�h�9"݋�	N�b����4�{x��7s7��1aa{]u>�8�x��wcb��t]�4b
����7K�Wq�{�]c;ɍųsƳ� I��\�
g,ҿ�_ �ogvI������������YWr�-�vrh{Cˍ��u�۳H+rMԕ��"NW���=n�Y� �m!n�BN}��\zgU��n�땬�]mmz�ϫ�^ng���|�t������m���x윱D�NSu'v�e(�q玞B���I���7��O1��r�����YM:�v9��p��ѽ�=&;N�XRW{H���^����z+��W�X��s���P�=I����,q]v��/Zn䋔�X+�l�[B�jҝ�S��z���](x���c��h��Hx�T��B7Y-��0�8��bqCܼ�{jX+m�4�i<�#wgs�%[M���e'#�b�q�x���@j��A���n�nͺ3�:��q`��'�����g�b�k�';����M�vG���cxCϠi��-w�9�;�'6�^x��8L�Q���<v����;n�u��%G�l]�<�ҏ�A��}�8��8��P='<.��s��s����k9���X8|g<wW�|��O��"��'ߑ5=��~��8�@�#�/_vWƖ�o#ɤ�	�[P���?��"��zn�ɥؖ����(^h>���%8L6�pK0 �F��rOYFrg���3YN�`9H�=~���^�o���a����X3nzN�(�OG��YS^٨�X��S����yӒꝭF��ML�;��j�5��!��Ul{5p)'4�mD�ނ^%�2�r�A�ēK�T�ك��d!��Z,�Hb��'s�/GR�A_v��9te�uW�ץ�2z5����X�P�hjJiqT��ξ�^���6�4��YV]��4!ܘ�YM�U�����Ɇ�ǀٟu7����e@,��M/������L��Wϳ+ �}'ޘ��fEvt��!���]�Y�>C�w�8a� d5d�F:r��Q���5�N�����Fv�a�9d��h@�WB���{.;�3�Nb5]g�w=$9mS��
l�ȩQ1Ýʳ3L�%3�X��v{)��-�c�)a�! ���	�bU���qrx�n{���x�����o��ͮ����؂�͒%>Χ�Tt����w<�~؟|W��B̝.�1<�۰Pjr�9�v���<%��m�	������^Ǎ��ӏ0���ʻY��>>.
Sb�N�	���_p)� J���pc�Q�j��i�$����8(�NL��eB�y�N��8�yk�g���w��ܹ�ە��Z���?��r��e�u^5DT����-{��NbN$`��D��l��ZN�]0 ���z2�&�� �ۓ�u*�䔯�YYf\+o+k���Y|ڠ&��*j����1Q��,��p�	Uǵ(�љ���q��ٌS ��H���?~��{��5�ȅ��!=�H�ަ��Lkx߸&�O���)���e,>Zá�Ը��vUU��<�G�)�)��]�&{���d��kA�����2��o�}��a�;{�u��s!���P|������������	��cz���w{��r���=���ݔ���B���tQm$C�ÂS9�-Lǂsj�D��4 ��ͪ/��Z��M�{�郴���Ŵ�c��]4ɇ�N�9�����SU�N���7EO%raYɪٹ��R���L����-�;;W�;�aP�n�K����ηm��-y���0��۾��(o����(/TK�f踡W��M��4J����{.�f�C	���aP;�!L��D�Eok�L�PaT{�
�@(Ģ |��U,�+��~s����A/%Yj�/��aܽ@n.�wF�p8!���ǂ��	��<ɒ�X+G��[6��i�rQhN�	gnGda�*'i:#?A��2����&�N��S��;UFֽ�ۚcۺA=� ���2+T=C(Rx�~Rsfڿx��q�H�L�]�-����:헀��`�a��:6�k24�lyb҆?�fD%Grɦ{5r�u�Ӥ��*�vT����0RE��L�1��H��o*�/��۷����fuȄIE��dp2�Rl��;z�B`8���shnl�Ǧv]=m�]Z�7�wr���L� ���I��¤�܂�z;�އ���2I8�_?D��{(����Z.�Į�L�j��Ȩ�l�j3J{]ڭ�T�g^�������-�!�o���s>��JD�P��� �Z9�bs7.��M�� E}$8�b{�y4�/;�Xv9e!��1�y�z�HP��35�ڔ�@ ÍkS��X��S"S���J���rTs�߃�L �@c�׼(���v�'.y�1Y��,�fd�N���
�wH<>/7��k+ډ0�&3����#餟��񛪴�$�N6�n�|���0�S��\ma�P��d)���y� �!�8d�S���K��!�J��!{׽�f�̹ #:�b�����V��4Q��.;�[&��\�a�5���͵���Wn��I���v���(⁯f�tM�F�}�q����ٞ�Μ@�TtmEe�yЫ��w٨A��N!A�'����!��jN���:���p�-CI�^���̤l�f��b��� 7�M������X��#�Ė���k'}1IQS�t�IS}|{���>��f�0R��t��� H:,!�T�g)�U�� �␇pR�ȻB���H�2�Ta�:m,<�txC7��]�Dp�9���r�����R̷Q�ƊY�{�&�)��R+u��潱uw�UuJW���`q��s#�(�*o}�H�ln�� �S��K�E��X>�ɨo)Ȏ9�|h�~1*�w"(}��uw�q�����?{{+i�b��}}�4��\�^0�[��EF(w㗯�����}ءÍ�]o(�JCg[W�ۖ'�|<�a�gm�����nZ�r�l@�ˍ��<oh��q���8���/iN�9!�u���p�Xu�rzv��=i	�6��m�!�h9�\K�H��cr]�.n̮v��J�9Raz��;�']�\b�cvHG�����q.7T��*��a��[����Q����8�ډܽ��WݼȦn�z������F�_��w�	^P��ӽX��_*RĮM�vETh��p��i�J6����1�z��͍�E�m����L�B����,�HW_���>"s��|��&5kg[���  Ӯܱ6w��u^鉤����y4��;~�,LϪ\�(�ݚ�ٯ<)hF��n��U#�:9"SD� \_��"DPwW����yڰ\��W0A�����=�eA����	2�� ត �x�\sv.S� �ۭ�G7c�)�}���;��1�>�Y��m��1���{�T���Q$��L���2,����Qu��3�oTlѨ�g!�ea��*�`��xȨNt��!a��
���˹�#T+=�.]ADSҥ5�c�Iܵ�=�"����{w�]�;�H�Gѱ�LO��UD�+B#V�	+�חcH�9�`�B쓠D��%��9�>�5�d�Gn���h�:}�_��G��j�����v{=�F~��r��NVzz�$��ÐE�h�}�,J$�_�go�7��p`���`��Z=0P���1�O�'O��&qə����w������{V��*����k"�|w?5�yi��bO@�UwQG�Rq�&	��BGM{�\���l/��p�(hTѳ��>����==X����Q!���B4$H~�貨,.���WT�c��xL��]������a��0��8ڝE����c5{�G�e��ә�w��O5�(5�o_Y�<2}w�z�K4���g[�i�YbfwA�%cr�����>#�}�"��9*W���.F�g�í�=�0� �M�ؼ�0��?e�LXڭ|�-��v���D}���ᯘ]���ѐ�uŨ��P$�kYh2�ժ�^B:?{�mfk]s.�c��j�%|E�
�w5��9��UJ�T��ta�HH&���o�:`J��G^��?�����3�E (�$�W@|K����7uϺ6��w��-�g�BS�ے6���|�}���2��^3��k���Α��>�P{PR�X�U����m?F�	�X��ܕ���� �i��=��G����QY&�ݶ�rp�c��>�k���(�Φ>�n�3]�Z��:QC�^kҺR�f�IZ�Z������0[ׯʝ�i͕�P��WE�#���%2ʂ���a `U��2��59Y?1KaB9�vg���.����dCGx�+�W�{��[�h�7�̝Z�Gr�t�����3|M�n��ziO��xh��C��pG�[�>����Sb7��rM0h8NM|<.7J͍��'#�:����	�:�>��5m����1�.��x2_��cG���j�g]]oy�yI���w��ݬxyA��e�G+�*�are�)��_6T�X\�T�s�}U1�2&5ų&h�\7�[������p�>t+���e���F�}WW��G��u�]곫���R���k!�$\R$��<��%�:(CӰ=�?8Y�r�1w����D�Env�w�����f�1A�j�0�vnR�i5Q�i��u��`���͖�Ú͐�d�H.����̑���q]�;�mnH�h|��M��M���FT�������v]u���)r`Q5G ����t����8"��6�2og����E�Ӽ��ʯ�-�|���V����Q�Q~��*��� z
`$�|l��h�*rb�oՕ��Gu��8��t�`^��^���;��y_�7�r�������X��ק�=�/nos��_�T{�E��֍ַ��+���@�P�Ի�o��'�<��v�e�	ȳ�g�:�;�M|�����/g��oN\���k�f��z�V)��h	&Q
9��s���Ѡ��8h�O�
�"77}�:�����x-�r޷uFR�o�x�@ Ы��=�>r���q$L�ܻ����`�v<�#������嗔"�8-�-��<��U"�X����5L
1�5oq&c7��f{7��<[ś��Jx��]����8Ƈ�@�H���	!@(E�ѽ��=�fg:�7�nq̙G����^�P�����z�㸙�jT���{��29e�^�[�N�l��S�<=�y�&��3{5�� sRvH�����5h�0�yƮ�㉨9g7���/�����M�օ��sI�]��[Z'd�	�h����ݏ&��ǜ4�4�`Cc�.��*�yFk��=>K�YZqU���	F�j��u�)�h	їo#'Z�����.=j��efm6/J�SR�͏�����
����j˂�1\�[� ��~�eGʾC�DO�jvm��d8;h.����\i,�#��~��uI�,�9Y�5|����=~��^����d��,��]�"�tޛ��y����+������	ݳ�zr�ʺ�Pyu�~��܇h�u�w5�����d��M�������M����jg�!���y8z	��Rp�E�\`1LTZ��]�.3���=�ZL
�1��ꓭv﫳�����U0�iJ<�w�T7��wk�e�\�]1��c�G|Kݭ���ksaMG�2ā�O��y֨�]A��,�9�����{�����=�`b_՛�}���ƀ��	(F��	���n���Á���H��P���6!CC���'��Mmh�w�??��_L���:ﻻuX�o=UI�U/�d�u��.�j.�h �U�u뚪�q0nj�wǴ��$�,[1�=�L=��#y�J3�]�U����!�1{��U㞹�4�M��T�wnޫ̗}��?^�O�螩˩��G�Bp�reJ��'2�VY�S`K�ݣ�,=��z��1W�P?5��M�PG4n&���>�u��� s����4�]e�h��!��	���Q�x�@e��wgvaz�
�1���5�[�c����+tȱ���^�9�"B�������a ��P޼n<�!�Ѻ��ӱEf/�"k��R��yq��%�����=�W��4�4s��� �J�&eQ��M�IRh�Ϯ�qL �tsY�<�/j(pJg/���\�&��vc���z�{pe1���Zx0��۝���I��B�v����>q��]plA�^Ssv�\�k��� 5�͸8Y���:���(����:rf��ϧ�lě`�Ivn:�P3^�s��^h`qo1�y��kDlEy���-��]��I5 $�D��#���b�f���c+2a�Ftǔ^�}�����:H�>��3Ϋ����	'1�p�F�xV,�5.��D�c�.��'Mb���D*U��b��ۏb<k)D�z|�ڵܕ��`.�9C��8�)nc�/ѹ�u�[\�D���A:I��\.�!t�9�{:�yx�y1�n%������>��C�xu�n;l�q��P���Oc���Fn�ܷ`҆��" ��ٛ�W+�gv��S�bZ���l��Ȏ'��-g�َ����݋f����\�辙�LvwrH�<
L�&㮬�jTO4T�9��bN�1j�f$�zg{%:�'��32�-%x<<���n�O�¡G�5k.�s��T��ɕs(��3J;���Gf�����`�E�X��+B�zw"�}��X����H�G�g\�Vx���F����Ý7@@�S6�lQ����]�F��nqj��d�br%}�5���AK�M��n1_�)Phݝ]��u$��e�����z� �u�>ގ:�=p	�O	@E�ʣ^^�C�8��S��{��:<�<�]WK�Ǹ�s� 1� X`��F;)���ȱF�o֫j}� �O5[T��oJ�t{)+�
�\�n7Ҳw��i��&� 7]����&q��^NI�����U���zr�RD�g<:�>w�HO)�l�)�J �J:k[�T�,WRbo�O��]-P7���`�Z�oБ�T�/b��"ެ�Et������5������g�����y�t;X:������qr*�:S�f ��]�ǯN�4����N�m��J�;�|��A���|�,T��խ�����FV^b�=�{�l�`�0w��6��&�3ʎ'=��[W��p��}F�j|�O��Ȓ禴��vN��l�{��Ms�IWCb=�ۥx�j�$E��y��.�4��Nl6�p�;�s����1�L����3�r��bbo���D�������P�^��<�L�	w���\+ɘ��<=�ɦ
L��P諎��$Jh�J,�d19ꐼ�H��ݧ���������4��ّ��Fk7t��מnt�7ѩe/��>�ִA�6�>컨��΀�A:dX{n��5���{q��N9 ��f��Kp�|���������6x�K�;t����w����J����V��	9�cW��z�qq��n�\�<��[�#zLNQw�!ܰd���ۍz���{�ۈ1����������n���nu�nnge�ݼ�ݷ(����hA�nV���P�h�Vv���7�zW�
�mH�ٕ̇��ݑZ�� �U��.��9-�������W }d���I�k����^�;of˹B̡����[�M*�{��_M��wF�^ѮP��(UB|Ȟ���w5Z�B�x>p�P�$��N�2Ni��N�Z�4��\
4��/3'�J���H���'F�N��ͦ��Y>S5oө<W׾tj���p�;]M���.-�Bp�,4�[����Qk�.�{v>�^�Xi?����zp���m�li,Z����m��Wl�']�&U9���˹��YO�^r�2s`��B��-�];��x f;�%2B*k�glR𷵷���z�{> MWU��f���ޝ�ۓ��x�D��'�<��0.�U�+�L\	\���j�:qg��fI�o �Æ�d��F�����p�f���S�vux�A/0慈�|�2��9]��ۑז0�P�`������ ��nj��4Y]�R�Z�;S���(��0�7
ሧwuW�j6ct^�9O�E
]� O����77Mt�㷛���(��#�2�mzzA���7N�������/����q`��7wL�����E�R}5�(j�{X�U�ũ�)���jfK�F˔;om�n�'^���Ӏ����VP�:>J�vG���B��ч~�s�8��b�`��ỷ�۳wr6&������]:(��j\X56���L,��A� ����z�#��k3o-TE4l��P��2=���آ-Qy�i��e�6�	9���w����J���BJD���i��)����#n>�v���?`����u�������:ޞ�x�炋Ý6�Ǭ�]en*ǘiP٪U� ��1�\������7��T��Ն���>{��n�6y;i����n@�JN�r�jj�mS�5>Cُ8��ƅ0�b��\1���6K�z�x;�.��)�q�t�g��\��p���@��%�L�\�qQ 5�F.#�9��}Җj�n�J�ȾEs�t�[�"'Tr�̾�C�x�\�t�3�ۻ�4,�4�d
9��M�>�tz��X`h�,*�S`�7��ݺ\%L;������S�5�RM=�gky����B�*`�F�c��\hiX�Y\�&m<5�,�h���a �i��uktW�����$NLB����dj^����x��x�����zcrgPʑ�V���i��[�,	�y�,�,!7�\�06Sú&�)�T�`(^\N�}���]�l�9�]�2�����,2K�m�3iԞ�iom^�����zr7���ac\�I�ޝ�G�)9���
ڽ���I���WQt��lQ��o���6�~�t��(0٧���Ժ�S�����n�y�C �:����ה{.��oxzI,u
��������D�����7�n���l(�֔�=Η"圴mIF���45T��g�Ѐ�Ք�u���#���F_m����ꛌ���};8��f'����2����d��F���U�h���P�ħڑ���fU���ۧ5����>p�0�"�I�]�2\�_־�u:OFfmMzZG�8I��?}�oЂp��/q��R���gI���ۣg#`�j�%�o}��^�I;	�i�������+8��;�n��z�.3��юx&�mGT�ٕ�_A_ *��N5lH���=���٘�@�^�*ۓ$D�Uh���L�p���a"�6Qu#G\��uq)��+7%��PH���$�Ts��\WXW�6������@%2 N!Ap�,qٝ�b��-��˔A�D'��D�\�磞½^9�F�1P�v�ח�n�H�O�')�l���A�AJl\�IX�	�s5�kf_�SS�N�D��跮�`B������^?v����	3��9:ϯ������[�^Ґq�ջ�9��1���.a�I6[�`i���u����\�V�����|���]:�f	6=���yIǒ�79K�2���=���~�t��X�1�= ��>���\A1�d6����_�]@�S�L*Bw���}ύx蔇��4��ÁL�C�TaU�>�@U��o S.�}J&Z��(h�-fw<���@�W����m,����0�P�@�4��;��\F{���<��8��ҝ7'�ۃ�`�I�.ֳq�D��͌iw"sf5.��Z2�Q�ݑ��h.ێh�pE�ٸZ��d1�l6�r�e6�MB=b�G<L��3�	q��v'G8���dyWiv��I�xf�\i�,V݃��ʖ<�ݹ�Phz�I��`ރF�Gs��)�z*�n�	y�;2WaU'Q�h��Oä~��Go�껹�W�n��^+{0���cu+���Q=��t��Zrr��Ŧ
`�JL#�0/�U����V��{�[�X$�j��c��'!��7�ke" V�S��Xw|'��Է7lP�ߗ^��r��+����A�m;�^�w�s��~��qGd��tpr}Ln��P�d�*?��%k��{(zܴs4�w[n��}��5����\��zs5Վf͸�"h�Y��]a=&@�����Oo�����e�Or�9H���]���=λ~��	�TqpR0�*��W�Ў{=ZOl!ar�g���tQRj��i���-X�����ȧ2y���>5���>PN��Mu���a�eH����F__��`�PjL�97��9�Ι��nUp9���;7ѱgx��%^�����A$0�g�ӓ�r��ǾkE���fxSre]�Tr�Q{~[����j��j�w�}�6A�4H�/����˚�4�Ht�� �ެ���=�љkuj�+�~��f���
)�<���9�+���.�4įaUݔ�tt$�PJ��h
Ya��s#ȡ�f�v�*���yr�S�\��(�O�5_nZ��X�3�N����^�%D�x��l�DH��OUX���X�˓�Wl��N
��|k�1f�l1�6��	�V�v\�nT#0�{M#cvi�����9{n�@�YSg�?i�Ur��׻He��4�(4�t���
�ҫ2�f.�mq}6���Մ$@`�&v��;�m<�`N��:С�e�v�h��3�%�D@К0���w��� +�+������������")ȹ�a�y!����NF肣�/3Mx�;͐�EAM��\0X�r���]ݾ�y0���;>�-���i�4.�NB��w��mj�� _y�������B��޹�om��Q�r �h-Fj�z����bl_��{���d���U��T�n^,B�"�4H�*@�T���Y�h^|V�'�&ayh��`��R{]�Y�C޿b�;4�q��*}1՞��a�J &:���A���϶��(M"�A�|3�oZ�,�Og�ꞶP\��;U;>���#(���1'F.�;�H
�53d���%��!�p�ݾ"����'`�p�FH��{l���z^�O��o/,N��S73�]n�b��^>��N2�ܚ��LOa+��h�W�����U쬁��F��:י��=p����N�"�s�fn<�slI�a�MG5�g���{6�c �
M��A�O:�\��)r�3(��u��U�UVx�ہ�<9�T�����{*ߠUU� ��zݠx�R�$ᦔ�M�>���5ll�{k^��:��z���&�S�i�8�g6�q�J�V�ۛ�606.-�ʅfN���v=�d'�#�ge�v��U`�LUe����sLE�Ѥ�(��V�F�e
"��]׿%y�F6b�������H��9?g�s��e� `g�&�P��`�-���%1�
39�CD�_�`@� B0ݑ�X�KB��U�T�� F�U~�|B�w�I�C�q����zפ�z�n�g�WO.9.����uoz�q�
 �jg/�z<w�����z;��] �	�"]���>K�沧.�(�ԇ�Z�WiIY�\e�c%�3�v���=����,_�u���D����]K���TDq��[��ïY?�6�h���h�tuO��3|(��F�ם]�?klԝ�i������.7ȐP���^����V̢P�T�!��;�Z�_Y�[����T����X9 w x'
	 �/���@�m�C���U�fV�X8v4	a �a��l�h��ݷ<у%/�;ќ�D��Dt&���׌{�3�7Լ2qz�.�"�*���F�8?�٧1�>�=p��)!{��&���)n��_z�shQ<��:AS,�i����+��[t�޳6H�|SF���N�.�i���a��C옦��ʕ/�������P򳇮��W3s����W~�J5�-&����>�M�s6�+����0c�kb!9�ܵur�>6��ֲ\ɽ���YC�9�N "���c��^/�5]U3��J����X#�y�r_;u.���
�LȨ龹�J��.-^���<F��0�y3��PLX�J����F<�$�h�LM��ޛA+�O�,�K�Z��K�J`�,�����vňz��;�^+6>����7+�����񼸚��+ҳ��^r��A�[�i6�t�~���5�i,��N)6fm��k7̅�	�,����XV:�zm���3����ŝ[���kjN���V����k���}���4=��.��"�i�|D�vUzT�J:�6j��tO/�=����r	�a�	��P�c*��le�t���3������P��`�A��`A����Tt���Ԑ�ƹ]G��=�t5�X�s����78#������]S��ӪS.M�l�Q��;��`ћ��%i�VB��OlMX�$�~Xs�3Q�X�}�u�*�����[�(�GJ�S�w=m �^ۙ���S�;�7��d$/��sƵ�;�44L�O}��Y���Q����ۻT�b�;f0�^�v����4�Hp�{z*��.�S�z������;�k�z4m7	�h��W��&V�n�,]b�oe=�q�}W�Ԅ������|����x:�s��I����;&��3Fm^��f�Ҏ轭J�/�[�f��
L{ ��>U��#�[S8�tY�m��٢M�H%=W��8{	�4��k�t�P�v�H�)g��m��_1���R)��m�K���<�my����SssnK���Ŝ�(����B��9ܧ+tz�ɮ�rnq�c�v�Ǌmg	qCV���՝�挘�+�����������=��"R����1Ɍ�y`�招`�*ְn��[5&�����l�PR,��2�d�����~�����uv A�Effua��;ܴ���6�e�Q�|��Ŵ�h���>쌞�.4U�;�M=�{��<%��7���.�<Mg�ѳHa�yE��8�GdGv�¡�_L��:�2v�;%k�H��ʙ��<Q�N�e���eK.����Sg�S���Q��F�_?qr�=`�6Wv��v���t絕M<�sv2�7���HD��0��ff�N�g���t����x^^���FxU u:"w�_���,e���6/��~�F7@ѥ�L��"&+��x�W�c�=�Ћ:�yj�X�T�'Oڥ�XKLo��xm'~�������P�5�u�T�oa�ӆ�"��p7��>�4d���{��������Y����D���+��,%'�|�8��W�D�9�'§�9�L_j�-f��N���e/Nj�8����P-B&��n0���/t�L�7��x�X/����q�է���(��T� )�7^��6��j�u���qtr2�Z�b�\�g��a#�!�"���$\6�#�D.պz��Eo�c �i���򯈜'5H̺�e�(���s�w���J}Z�e�]z��F�����Z;OK��`��E�s�����n4�I2,,J*­�fj|8<.���j�vH���]/*��x͚q���vW��a$�]�^8Zx�*F�ɭ#"��Ò�I9<j$tb�m|P`@p`���\]!��'��a��⠴���~p
h8 'y� '�ګb�`�qԺ�Z�2	�Q2oi�af�=ū�h�u��^�S�p�
7�;Xa�D�!��o윷ƭ��k����X@���ȡ��U��cs�ٝ.�\�w(`�:�Nϼ�6"3v)�֧}��ϓ����	�O\mGn4a�`�A�<o7���[�o���y�?/�v�9������/Q��g�d{����Tس�]��F�5�x˘��l�13�5v�� ����C�z��ӂ�k�V���;[[�R��֦�\FڱP�ؓ�3.�A�ie}�+����˚v}�!h��v�����E�`������Y\blh˕9����&! �r����+7{ӗ�t�X6��@�霩�[�a���ܕ|=�/ݦ�[��«�mݔb!M���˝���e4�0J`�9iZ�6�f���ґ|mZ�QYɎ7m�7ԍ��,$6����W�L.�4;����B! �l�PHD��ݳ�|�W��1Ȱt���.�`���[�dF���ٔ�V�Z����̋j��`�,��a�BU� �T�֐�������}[��p,q[Φ]ӺS�&*����������r��O��w �i *W���vZb�Nf�Rv�ڤ#�w�����Iа��"ǳe�n�2�������}�{;}_=�35�խv����x�v�tO��`��m:�y`����7���!,�c�g|����Lb�®��;{5�}��5��s/�qdt�K�Le�7�Fh�s:�T�����mu�nfR+�M�wqM�.&:Haf����Wi�O�`^t�9 ;;/o��ÕBɐ��8ٷ�6�p��>�֩�Ǒʜ�O�۱�Ċ��yתi�鬄 �Z?t%� ����SsM���ۘx����ꮖ|�c����yT��Wz߳:���g�Ԍ,D�7wM�S�%�[3�_bИ-����^���C(�ZL�W��t�#{{���'�2�E����틱pI+O��&��B���������p3<��ƛ�s�8���yڨ?�����Sk��Q�.�����.��EQ��Oe���הGa5��IU���dtO��ݙ��pď&`� *C�gft�	V������v�a@�G$����)��ۗ�h�R/��KDg]��|g9eJ�e{7�ݛ1�cTa߂p�&CN)�͘�|r�ʦg�5;z�,�*G�����yv�f�쬺[I��ð��<�����~ɑ/3@?����MW���/�>8m�+%�ɇ
�p�?�|;y�#U��+؛� �wX)��c�)f!���a��\��q˙}�Wy��Mә�r��04l�!?�(Nh����p�w��n���]��t�����P�*�N���;mm[����p�zh��9yy"T�{�˫��R��4�&}v�ݘ�o}����o}ϕ���\��k8O-Tw�����b	�ἰt����ǇV��O�;���{��˯��k��^F�)����ᬈ\�?�$�Iс��8@�k�EN���w�^��FAz0�'|S�u��i�i��)��(Wvw	�9��X紭u Rs�� ������_��/� |0:��g���cND9����5�KAt��}��{F"�eN��Z�o3QI�P8a�v�{�l����ٺR�ďm��;)��0E���ܥl��F����+]�:�xGx�u�s�1�NȒ�vq7���P0d��$zqP���+e��!�#�8����-P�kg�i�b��-}>51ҊkU�BA�����^�qS��7�^�3=�t��2wFWL_x�ZC��(-���"��,�Д��ǶbN��O�^[�ݷdL�qPq����L�U�Tn���r��qL�m���4����U����,�x��ǜ���O���Y�.�sl�t��G2+ Ѧ��6���\�'>��e�v,�P�3ix�0�gA��e
	5W��^̀�����L+��;{3��������u}0�n�x8�q��ֶ�����g�a�n_\���;�,]q�\\��A���on|�]I��]��ָvu�h��n秷>�ktq�W�z벯h�*�d9q���*q��AgT�Av^���֤U��V���z\u�>�S����1�	u�u\Am?}�ػ�T+~H�����(i�Pv�7ÌFn�[��W��ƞ��1�d5�ߦ��9F��&�s�r�D��~�y;�z7��K�8nD�y�o�I�T"h�e���{v{��!�[PS,�Bk��T��{������޵1�"�H ���p�I� B�ӹ:*�V֎rݝ��;�V�)��3����;}��y���T��9x�LN�\�B����kn<��yJ���I��V���r�H^�{��e4�},����2�����x�v]�%#M
�!F������]t;��r}x]_zn ;��n}�p}C0��=]�1Osł��!3��8 y��x�h�Ȳ��{}Ӑ�0z��0�������6b��'<���Z�۫l�_V���:o��B�s�Sk�pyf���=���p�hM���]:��7\�gٹ>9||en� vc���ٺ�Vh�^��2�v�ٓ~R{�I����t���c���o!']���t�] �_$�E1�ɘH��7�GE�}������IHo{�+�RO�K#b����h���Ue����6� ��Y��9v�w�pdNn �w��кST:��ج���e+�{L%s��̫
&wW�-�L�����t �����Y3&r��j{�>�9� l��{��;r�C괟dV�v�
���8-H�ֆ�:�j����U�:IOd�˫�jvnA̬�Zn5O�R+֪wsT$/C�YK�"fp�zgR�B��(��:���@o.��ݫ��kulx#�Nw��hoVf�H��k�Y�+%w=��KćJO� Q�S1�NyZe�%(ڛs��x�;�M<��v�c4f�{�Z�wE��1<�\r����g^+��j���<�F���Oy���p���&��B��l���M"�&w��AL��l
�Ol�r�s����u�Eq��8\��;h�n�o<�f68�v�t�y��1��UHB��vkj�^S64[�Gs�5�?lr�R+.J��i��ϩ҆R"��fHwMĵ����&�J��Y��-�h�/�a�m1ٚ���X䗊�r��O��rl:/6�:�ܮ���N�{�@`<���fQ��Zo��^��[��1�=K�A��Zk*e�vf4.vʚc�OM@���hLg��7����veva��t�#ӳ���8�5�A������h%�/^Vq����]���-V��>n��[�U���oL����O�������s��@��kfc��cX$�Y����n��(6B��ق�$J��'�iH�)�������w<ƪ����1��@n����v`82dմ���I2�(��*WZ�UU�,/8&����L;v����r�ٝ���2��)��\q8�7��N8�yC����.rn��f»;]�7\�m�����n2�oӻ�~=�����ɹ�qP63'��O�'��#��kgvƅt��^vxܣ��7<������Li���A�.�p6&a�O���������<n��q,	�E.�]ss���@n��].fv�R����pۮ.ͬXU
t$��!7�xCq�6Q8�\l<��;����]�� �xZ9� ǔ�s�n��b�ޏ&թ9��D�{��+מU�m.0qt�=�۞��kɋ�tۃ���wse��q�Si7<�⌘��l�;�D1�{�{q���˸�e^��&�Jc����c�~����=�1�u9磞{'F<����uc٩����uz�q'���n��YQ�m���b�ф�O�d+��%nQ4�v�L907gy{P�046�ݱH��Ɠs�3)g�Iv�jt����r�7[�z������Ǌ:\A�'P���;��61;t�2��ˈݮt<\Ŏ��,��h�̓r���$�q��>����)�r�m�}�M9��\�pI��tMx�4��;�I8���GvD�¦{&;��M��wts��8uvC�繺a9��96��.lb�&w'�����D9�&C���=v�p�l�f,���ː�ŷ]ԜHE�F�7;��&��N�۪�T�^[/8�')ʜ�úk���ljNy3Ɨ����Y���]f�s��oyͪ/.@� �{\�{�v~;�>���g����6w9�林gb�@#��n��t(�.#Q��\n6�V�p��3���;h�!X�<rvq��L���{7�h�{6�O����O|�y
�۶�Gn���Ŏ�"�yy�l/h��s���pq�9ݞv�A���'b��Gɇ[��=��,f���=����W�n3��y� ȳ�ٚ�oc�����_����B�ey%Vп&�o.R���ukl���t=��ݚ��wj�v��d�l�i���#8��`�2�+0Y 	�#�񎙐9��#���V'��##V78c���.����N�{���=��T8J�[:�����_�Ns�X~�^�	����+�]~���;���Ft�%\l��	8P�Y�|`��>ٲ�=S��Om1v���޼Q{\�qH�$[`��ޚ6c�j���fjf6v��7ƅM5��q4GoM̹9��F$������]0�r��2�+ʒр.W4�V(�g"Jgg<ӵEw]�5�zd��=\��	uUn�3��]�l�}���n߫,�@(*�%b�D�m#�5~�{2E��		�{���yN���}��P2���\�d͊u.ϻ�\��w:�J�  g֮S��~~�j]׈{��邙tSf�Q�>~�ߝ��s���7>\��w+1g{o)��'����=�O��RTO�%9{�<˚���K�>�8���*z�@R.
!"؀.�V�C�qv3u��^�K�5ӎ���7�K��0
τ�[3�:^���t�<u$�s�cQ����������s=��{z}(��}��[3�]'!T�^�h�����|3�޳���̻92���n�`�E_�a}��ó:��\��ݕ�v�^���nΦ���^��p�d*�$�]fc(��e{��{��q��t	���hڨV_�K�	����s^��2)�����6��
�F��#0��)�{~tM$
V!�ٺ�^�l�YC��|'�xj���h0���`�5g'���8��	�d�l��Q��ow=_q�A���|�*�X�ZB*����f��h��(��@[&5��j��'[ٰy�-p�76$nr�g���I/&e�]�ZQ�N�p֑�a֋�~�Ⲡ���i�S�V���=z�WORU�� T<΄`S~x&��y����#@RAQQJM߮_�q�)f��ιUT�;��m�r�*3�_e���u]�i������V���e�u�ljی��d^�^�g��e�pTC��jdt��;��)`�
f���;`ޑR������j���*�巾�',Æ�h��p��|��}��j#c&y�'� 6� Â�_�pId�� ߌ�����/�7�۷At��.����b�	������|=�N���_p��ϗq���?*E�E�j��wU��y#R�_(o�A�z}��������L��q�5����᛽�L�$*�\�VqT�k�W
�Tދ�^��r�����5������J�6��(b�^ԯ��^��vTذ�@wr����:J#�����zC�n�Cյ��\��;�8���)��!�9���<�Et���N�9C?z��w��"[wh��;=�Jlq���Ξ�?p����V%�o�:���]�r�3���p���-�Қ7?
أ�2/!�Ka��ｏ�f�7{ݗ�2��x�fI닮�'=o�'%u���o�+���C�W�cwF�)��.p���%,�F�m=������j�>��ܵ���<���J+��OڥH�*�+r�����kF����c�P!�=��a�%Y��9����|��%��!A0��JL�ި��L�2�����*z$((�Y���5pu��h���A�\/!��0�0�8hi�aX���Un�=����MGW��ƅ4�G=@���蓷]82���0VŻsb�+{$P���WW��ݔ��H���tђ�Ւ:�^����`M*�6>=��n��^�8n�����v��N�<�=gN�(:�[5O�n�+A��Z�gv�o{��B-�$�:������-��z��'�xn9�)&sFv���<�-�1<"x�%^O�=sQs%E��3��ܞ^��>꜌�0������b���]��:��A����&ț�ɐ��vkr�6���;[�7�S��Y�s/��k��דǘS$�bВ�R_A����+8<Kf��r�뭝�,L���Nm,��c�t��qz���Zb�鼪��9��n���32N������ռ�V7&�(V}Aceh�=
<�`���^�Z�Ezl����n�[��:� *�#�ם��`�@p"��sاH[cз<��n����..�G�����d�Cv���Z;pB�&ٸ����6����r����OV������۱&�n�:q�]�F��sۏt��,*.,�tq�ZDb4ku,�@�Ğ�,�z`��ՉQ�C�gWQܫ��A��b�v&���0M����j��OE��ᣉ����6��Ǫ�f�A�Z��\ь s%���S�9����l� Y�EfL�?���ExD��vT�uO:�tvjЀa�8(P����Z˸��E�rw������f�oͪ����-j�cy�mu�{;�=&G�8@�L0�"�H8���x���px��su:�����C^̚c;��A5���#/ݻN�ߋ2o2��jm������l��V	v�`�ʪ��I�&6S�=��bi��������NL�磹�)VX[u�w����5}1�#IV���*�U���`�Pd��6����k�����D��[��9Ս���T�f���\�Ъt�t�: p��A�X���:W�<��V/����Cw<H?�I�T� �u9���x�s;^X����8�U��݂���&K��5�������J�no���{v��W��a�l��N�܏f��d�0�"����/)`��#^�2�������\
���ff��\pӠ���/'���XA�#�"��VVY��e����:E̕���u�9������gĸ+��F*%B�T��d���xw|鋨�t�	���U��Lg���N�@:�,�lL7̵o��ï�(ͱ�[�|������&�Q0	ɍ۷g�-��ۘ��<�6��k9�98��Q͝���L3=g���-�˅?dD��I��-�7{{.�[�>����&w��l(h��h���A/�'[!��'�շ�u�~c���7��46ҿ����ˬ��D5��C����Q��}�o�ða7hn��ޟ=���9�7�q$��f�'M!�v���.��3n^�υf���{�bN�L����}�C�ٽ��<1��Ʈ���X+��Tэ����#��{>�>�A	W9Tg&^�ڍ,��l2Z���9�ݹS��؁5~��W��4�y_vEn�2���Yꎩk]�
�ƪ(��5��1#[���Z�36�������7|���H�ɼ�8
T�����f�n�ڗÜ5Y)	[Ԥ�~��F�D�yU��/=�^��kݞ��[�%T|.�����t;Ǒ:[e�aAAš�DnhJܯk�ЮG����U�(�c(� ��IH]�9�u���mOj'���'�zold�u/QpDge����5����ܰQ
,o�����tc�z��T����rI,O@�C:�h���!Ug:��
c2Y�J��A�;�lQ҇7,QU�b�rq�	1�Wt��IL�Tz.(d�o3��h�g�`O ���	p��cيUeu{r��� ��MjX�m�`���
��P���"g��#q�6%5y���2r��
��*ӛ�1A��w�H�D&*$vr�#�M_��cᑲ�W�"Q���$* �0�w�F&����l�zSFy��JoKD�YݮR��^�P�+��W)M�]���Ɍy�q�n��!�F}� ��smߋ�v�>�>��^vj_=e�������� ��X��*��<S�Et�s3�v�)�3k��r	�
(p���{Nz�!�9`	����>���鍯щ�΂���s�ME��2�+�0�O�xT�og[^�i��/]n�m#yFɭ=/=*��� O�T�H�}J�{6L� ͽ�{V�'n��
hMF
e�ɄC57^�wg�� ƹ��</>�������`���ߏē�ݷ�r��x�� �WcuHO��#Mi���vx���l���r��,��NQ�o�]�*͍:( �r8�h%�����OzeNhaτ�G>q�{��j�Pl�\܌�<W]��J�����e@�-��W���1�Q@��~;�s����E�E�f5c¦��;�{�Zjeg��K@�Q���LbL�W��|�Dn����7��"w~Q��/��L�/i43%+S��uCy���,��8n$����;r��mnt{�8��������Z�#�F�3F_�l�f��z�����(l(0�p��^-5�h=��ڨ3a�/��8�{���c��{ՖO�K�0��+g����<r�$y���VSIұ�hW���;� �)&!"�2���{i�1���E�~�s��\�wI]�4�����B�e�2��y��;QBV�K޲�U�~mL�T�
�V���Ks#@���Ap�|��6=��]�Gd�8v ��~/?�a7O�uJjٌ���ُ	�M�8�Og�m�$Ri&J �ؼ�t������n�J}�LH���ю�:��>�+��	�wP�C�<���Y�7����+�I�TRV��T��
?-�f�"�a�?�+�����kc�2��2sє=�ȴ���=C�m��t��x���w��2�mT���G8&!�Y'�s�nŸ�W�	n`��d}�}OJz��$WB�hz�__7�������;��#�O:E���͇Z3�NK�ú��(�O�����n�Mh�F���=fw+�H݈�&��f��/���C-��
��hѴ3���ʞ�������5�do.B���a��w�y�hF��	÷��"�镱�ݦؖt���y�c�.!��W�;���z��k��3��Y��yhz��(n�B/]��.�Z�7Y�y|���`3�[o)m��'t,����4Z����NE�Ƕ���8���?\q��q��h����y�pF���7�l�Q��I��ϔ[��.Z�t�㴝��B�(7
�I-�}W<�3�
A���&��[�j�#�;�Ö9�O�{��I������}���=�W�6u�7����p��`6�����_�hvm���fl�Ʈ�@B�&�u��q%�$u��8ߘ�΢b��]ꋱmd���`�NϝVJ#��WK�����2��@��G�TfN\����v9)U��z���`1
�Hi9���z^��|�<W��v|z�ź���u��7���ݯ+�x~��Qw�Y�}qX�eɔ�����ɝs�e��j6<���K}��M
I��mQ���e�ٶ�2~o��ڝ�O���.���dw�|��m�ڙ���s�dU�F�T0oyd��67�ƒO'6"E�r�	I���``���|=	��q��<�k'$��]VʚTE���Y���OA��r(�bPtd���<mM.蛈���HE�`��h�ZwU�O�q_B:R�?b�w�.ܝ�H�s����ti`����l7�탋�fv��]F�DF��t湺0Z�21�tw��b�FrM�XInY&ߡR��ȴ-�]�����Z��b�����ߡ�Pf�sM��\�v9�8 Tv���d`����d���+/�p��p�<P�/�͒��0����=�<����9Ȇ	`�8Z��h�y���{8���b�͟b�==�`����x1�>�9]�7y�$&�4��zyG�tSV֒��1����_�I|�!7���W6��<A�a�:�)�2u�ۃ� �`k��޹2a{r�[���jN�y����yp�B�����Yy6@���6M��϶��"y�t\�A%�o���w���4��5/�ݪ�&�|�Xp&�ssڅ@أCA���Vɝ��L��{5MNj���w��hB`i�^�a��嬚�E�[�ysN/s���R	��c����p4{r�SՄ�=+v�#N�G����Щ��Q'��:_w�D_|=ѩ�%��Q�Md1���`<7&�F=����	z��ő|\ϲ�����
�+����	ܖaC��x����y�t�b��l�ɻr���1�F��yXϽ�Y��}�-WL�
�il����F2��HN����������k�N����Ɯ�31˙�zcU�U��y��`�Ht�$�Tl��c�*�e*�)ˆ�9���f;�������هm�\Qؙ�I�=/v�C��:G6tp�E��I���j5��Q�B�/c��S��WG�>�<c[���˳$����ƺ�}�A`~�@�A2�{���y�)���s��U/+{jS�ېЬz�`��(W&�w^��S:Ю��M��Lz/hg�þ͙��`yJ-�I�%
�Goy�Ҹ����%#�>�"��,��L���k��)�"C����4�jo8Y�u8E�]��&�_�VPG\=~��N��,����hJ�]q��^��b��g��ab��;��H�3_��h^7��S���q٫��qX�~�;��o������ $�Zt��l���KB7����A$'
�����X��L�l�՚cm��3��toO� {d�L�ˀ�� �.οO��uCБ2g��럖=0�b�{s�5�}=����BIp�K�����nOpʇCߝ[��(�����ug�2Ag���t�*�v�1o�yt��u�����^��6=W�#[�����;o���{��e�D�%�3恴��w��P�p#�>�3���CdC����+
p�$�)˶h��ʆ4�\�uα���[S����ۤwv^�Q�w�`�
���;�.�j���o<�ݼ��0��W>푣nc��O�����b�t醃�( �������fg�q�� �m���.1\%�?�=+Q��{��8�"mWt�{ǰ��z��WB�i6�O���c�0lt����0���+�=��5r!�ua��	�79ITи}'%3w�/%���Q���6�s��c1��O�f�;�T3p R
���n�m�I*L�s-��b�{u�y�ų����u��8�匈q�����.J�7��_4�Ø���Հ��Y�9w �P���V���k�c�n�I�vU�Ҿ:�Ir8����3��U������u{ʳy"���k����/x��b�o'p�y�A����Y(�]�o����X XJ�"�;?s*�\De�=�e���E���c-�T4�Xai\Ž� c��>�4��dE���сVm�����s�8��Tä9NwKK�t�g,]�͵�_�o4�s�ٕ� ����Jf:_�tv�Ø�q�ms9\yd�vnkx�\����ج�U�T�*�n�od��5�u�������_P���=P[�o#eu�3u_�*mj�z�g �`���Z��q_V�>�R�g��r�}�,�]Jȶ*�p���u�>�Vl�r��ƴ;H�;�]'��P�;�6'#�H8$�Nh�{�# �[��`v+h亹�[�Йd�a,p�)*�M!s�9�׽a���ȑ1IyϮ��+sC{�13�M��1Z�a�{G$���ܩ�+��_�eF���w͙u6@5�A��.�u���5�j�m^�s�7�����|����޹�#��a ��Rn��jړ �U=94;���į�	���ƶ��[ݟt5{���Z7�f��˞������/05��6�j��1�{�Q<�����Y91��#x[��k��� ،����� ��:��Z�c�ڀP`7ޟp�"t�܃7 x̓*����S����.���xe�4,��{��:��e�����P�t��`��L}=ɧ��^H�["�d=Ͻ����^`T2fn[���vT.}5L`yIz
(A뮲��gg�?XW�D��������	$߲d������0$�u0Z���d��F�WvUI��*x�$������<�\d�]=�����n2+�@g�]����80X@�ڂ"�9}��Mv�PLa�aA��{�������E���V�4��,�S�sl����%"�m��!�,����+�𜥸���ǺwȈ�6~hY�x��ۓ�cW]���!�Sˮ��!3��3�*נ r4$�!�
�k���p��2��{���z�IjB�]Z΅~�G����\�@B��w^�f�*U�=�Njw�]}�^�8�r��%��z���S�Ē��SL���\�^����L.�b >�Me"�:[�i�j]��-M�=�`�ĺEe�bi�!����Q���+��U����gHZ#*;;]	z^�Q0-v%vn%t���ؕ�C�tG6��[/���П�龑�ϔV;+x�b��P�ۺ�ϥ�ǂ^5��s��&�f z�ٳ��p�\=���H���[WR�Q|�iX��Аu�FLs�عwm�:�g���G`�0=GN7�*�O]���b���n;E&n�;\��S�"�.�*�@(+��kD` -ì�=�,�Yg�&#�,��Ӆ\�n1úpa��8H��q�����LIn5:��QV+Q!u��,O������J)y�L��-!�G��7��7�ZG�|3���S���ڷc�; uK�l��y!��mQN�#����cӺ�O����y`6ջ���М8a�A�MhC�5NͿB�JB�b�P ��!��[�͑k��������;�@�]ut��6��<܅�z������0<@�|�~�^M<4��z�V����:�xH��{э��p��Ӽ�u��l��
" ����0�V\¢����Y���ߥ<9�Eϼ6�F��̓Q���B��Jo�&r��3Bt}���k��z�-@����}($����z�yw۾�Z���P9��epȿ<�(�5�T�(�[:��d#8����F�A�3��)�X+wh��ɤ#v�¤�u��.l��g�N^��Ŝ�ʹ�qܻ+Q^�}'O��{�b�d���yń�򚼻^:I�������^[����L�K�n� >��$�F�B*�io%45���[ ��q�w��c�	�r�va�}���^����r�S�U�/�^��=8�'��8J"@.��r�7;si�X��t�/�v���K�����"���j�ÆI2K��[�842F�PĤ��t7��^~�ޅ������?A��������b`_��bƉ�c�p�{q�ɼйv��
��w�2`�R��Z8��Kc��e�h,��39��yX��XAe什���SI�:i�y6I��7H� }�+���'�9�P���yY��t�^���SK1��ʗwQc0���|�{-@�5���a���߁�j��������z���ܮ)�����o=S��лJ�Z
��s8̿VRV��S�V5���4�r���4f�=J�kׁX�/����𻚵ƶ׸�Y��y��~�:W"���I��S�9u9Uu����� ��*�H�b��&���V���B��Ϧշ�V$�b��3Md��t=����!���}ӟy<��zL#�z���A�ϻ�)��e&�m�.���?�+r,�O�-S��멖C�=��#Î[�\��g����>EV�ҥ1��U鬹y��@�a�<	����/Z���`C�� *�	ԥ�������{{r#v����^�-�?J�Q)Rj�$tm�����3Qm�;b�Z�`�p�0� !t�n֜�U�״_=u����	����(%[�h��;[�L7Z������ZSE'Ǳ�j'o�	�3�댈�b����F��'��T/Jr�(�y��!G>۷��gAD-�I��a:��mqݛp�ų��ޟp��8z�rX}�dEoOV�Nk��6�_�ӟ	�6�����U�Xt ��Vȅq�I�~&�a��1zrx���d+�Ս��*���H
ܵ���B�3s0i;�-���4��eU����4R1E�u=�m{��h��L�gh֚V���B��,X�T��c׾�n����yOy	�_>���`��
��E�5g���T��^b:�|U&BF�ٹ�OA�QUإW���}Q9���V/m��5�]v]�qd�	�;��!����+�}�R�{�55��(�_��:,Tgz����wIi4[FlY�X��&w��<��_NpȞJ򽟏��y�u�0E��(v���w�ގ�5n�a�qn����$	�e��
/�~�m���TW*����s�f�eă^�d��^f�wB���E�(�ɾ뱙�����ф�
�9#��n��`����p�������V�䯋�vl\�8?fs!��ェx�����sɲs����2�a$4$� @�@b�����J����W'8lp�%wZɴ�
���w��zrv��2�7�i m"�um�ԟs,jC9r�@�S)�3##�
�@<9�q��>��;�(eK���R���e1�4R$�Y{�s�H�i�#=�H�X�}��ˮ��>�P�]}x�)���=r�� N���F�\�Ď���}�B~V<�=��Cg��B�ߑ�HF�� .ʳ&�Q�^�ۖ'GnV�xi�Q��Q�'}762�!�v�7h@��F�]�:;�6٤y�e�rr�9��ƍ��!�6�T��R�z�h��jݵo}�4�D8L��,2��(��,��n���k$�d)p�U�{!��8�wt�nL�t;��B�\���pr���7{�[$1؏#���^�Z�����������<�^��z$� ��l��ʇ��
뭫˦��=^��a2���19�]m\��6v�ͯt��n��~<dC>k��=8��A�T�s�{"�<�
�4�:�N�ᙵoro]e��sMd���5�F�n�R�vb�f�QKݝ^�\�U��Y���j�E�K?Nt����~��m��ΆU���Wx:U����5��U�w�գ�r�q�Tڋ����k+����6�n�Hu���vI� �P�*%���-ʺ�����)��M �j�y3��Η��ݻOn\!�c��^M�Uu����x5�'<��АՋmxwd��nO��ui:���ۋxL�y���r�qv�P�q|;���gԥ�[�o��|:�{r����tZ�ewOkq(���{b�u����sCV�Mլɤ��lzݲ-r�j÷]`��LZ^x,Fc��\��7r��4�	3�� �mnwS��%츤Ys�j��,ZUt�Y�p�p���Tg���j�K׳�V��Vm߿Y�I�[�G�~��7
�~u=�|w�ӳG����q���ʕ�n �Ap�'�.�����V��++] ^瀕����]$80a�)�3���eu���XK��&�Vg̀;����خ��7��Ѻ���Ċ���}8:��s�s���]^��v�r�����(j8�WWNi�I���b
��jkK�_���2Rt���
�Dg��)�a�m��k8v���"�e�f��߂p
!�Amn�O[y�x7)���|�_���������`��h}�E���NJ�?G�9*�fm�oa/�|�W��$�����T@��\�\����<��|���\:��2j�(�{�]�5:{s(�Z%N�ުع��gL�R	�M+Β�>#*�c_b�|������EH��l����=S[��Rhv���r�J�2fUۀ�n�@��b������M�F���վ�j��E7�ū�Ք���U����;�	��B�ǵ|0��S�z<�z�վZS�M�V���y��<6���y���.��sѤ�1�E�Ќ�S��(�v#�rļkrmד&�
�I�a���2 ��y�l���"��Z[��[�_��������>�sI�I�]'D�	�̘oX������z��o�U�ĉ\�{�R-�FmO��ΥO� ��85��0�HU�o˯34��_��n��Upڀ`쫗���s���=�}|Щٍ/�U!~�k��jK���������A�+��a�ǯzz�>��S���I�T��Z���G��'Z�M��m\Q�kd���xɯ�2��2l�)ED�4R���Ƿ��7*E��î0-�����{˲�J��m/3�e�w�5�׀�S�xw��1\2X7��}�ަ�-�S �k9K�ïrbm�=�:P~1�xߜ�츴��Ct�Y�ظ���� �����v� � _� Y���:�nA��ݓ6ۺy�/kث|��|H�p���>��7R�{�]��` �h����V�"��C����i�ݗx@�.�ѣ�#����hn��w!��F�gn��c��^X��77YZP���8 ����^��N׽Ҥ���2?:�k�:Ʀ����M7�ه�w�<�����;f��S�<.¢�F���%��h��nfvjJ���f����1�K����du��کB{؍���z�JeI�\尽��%
\�1ASi�Vc�q�sϑ#j�nu�G�F�^I�wM�+L��~���l{��G�hA�v�ͻufw���w�hC��D���e�B�??z@�םM�����Vy���h�֜�5��N��q����<;����4��'���Y��81��p ,u��u��w�:�Zף�2a�wx��������%e�ű��m�v[����N;d���m�qrP`�	�&޽�Ҁk�*^aGh�/ʼ�)�\;Z����각ݓ1��̘	��	CN^��9��a��щ�@e���}c�4�ו[�^=����]�'�1O��H�z�U徙�]�+�C��M&��r��i��������$V�*�%�-�;Ε��Q{N.����8T|]rԤ�,qȖ�U��Ǎ�bˆ��9�ñ�̎���M��
je���Jn,��O�iܹ䧯Byᬀz��	�v�@�_�ٽ�<�i�iS(���fL>n�r��;<����w��/Jm��HV��p�����r؜n�7vݚoW����a��[b��b6���\�GOh�C�0o�������#	�M^��m��b|9��T�Mt*�j�����z�RT��6@AB�$f��w7=�W[�
~5"�>Vo|�n����8W=�ve��X�8��m���)�]p�@0C�:�>�P3�w+ï��\��7g&��go�j�Lr�������L��C�)�Bi���Voxe�߉�qU�.�����aچ��/=~��Ѣ,��\���S�o����CLӢ�l���5�|�<�^���mfv���xp]����ʰH0���שQ}�/ݮ���G���+Z:�kEm$;╒ ����0�.ϩ��n�?<T=��� ��~�!c���zQz������
>_�s��ƽ�6ڼ��CH(�" >�\h���0����]���¬�Ű3n�p��n�DM%�@�kt�J�jG�2�XK�Rs����㎷nyq�[p��r�Dv3玕w�7k���ɑ9x�<\�ݙ�Z]ɓ�=7�G�w�^���v�%�ҐnƗ�p���<��<k��0뷑'��vY���<m����kl+����e48y:N	qg�[>�<=��1���V3b�#!�NTv������Ƿc�X����:�q�D��q����a�+��^}���?g<ܬ*����]�wI��a|K���o�0��c��)�z�a �Z}��O^V�r0��3m{f
WeL�e���s�k��)<NNV�X� ��RH�@���/!�ك(b��F�Ň��*�a4j�s�q�ֶ�:�+V�<O�%.3��:m��ӌ�1Z�3i�uqn�^j�%�V�)�ݨ@ljP�4�z��pf�����*^d��,�å�Wy�H;<�O�w����������as�W�%{ٳҽ��2b�rXR�{|��]�'Ċ^��"�!.cE�	͍EoC��}4�7Y�f޲�2����t��y��{dO/�i���Y*�1x�~����f��&�t�tUX����Y�K��3�^�󲶅h2��C��¹�?_��X�?4�=�������c����Ra�D��FN� �*egs�p�M �fm{z��<�|9��g	��7 �I]_Pנk��;Z�����T��31ncu����*�^���� ���`�2˾�P+T���q���x��h�K&N�x�ە�&S.ֱɈ��㛯3q.L�W��.�$�V�/x�\�w�U�����6�zP2l˚e:����U�xN���r\���oLt���GI�&Pbv[�t��is�c�H۲g�nf�\"���gƝ�\���|���څ.��qX��YSK��B_k㮦Ю�*m� �,�pXۗ}��w��&��o��\Լ$�[�{m�O3�U�K����;���GߊVz�#8�S�wB�iI�����h���fR��|p6z�鹘=�r�f��}$:Ȟ@6w�:H�/o��=�}�&��X��h�&��Wnv�[��wl�������n���.�xAL��`�lr��q̙�"�Q[�h�<N��Y�q�Sn�)(l76up��X�U���hҏz�nƔ�)��h�n��}E�v��:ۖ�7;VYT?6�3w-eÎq�����G^� TY]���Ŷ��C*�^Ĩk��Wlɷڝ�X��_0��v񱛂t���Q���OGT|�cv��7�ntݨ�VnQ�af �x���g��7��8L���Kq�j�Iv�����2l��ʊQnfK�[HsI wIŕ�)����tv�ا[���t�E�wPU`WY���h ��(%���-�Fv���ogZ/w&�=��@���V��-�4���c6a*f�zic�є�&Nd�Bv�S�n�K�G�aےN.�^��Z&�1������hBA�'�T�*�X!N8[�U��v��4��R>��[���:ځ9�����q���]vLt�/E&��C�;<��=&a�y丨�"c�k�Z�]��}N��DlQ���c��ܚK�oQ@�	]G\u�3g�ŕ�v�V4��8\�b6�c�&Wru=r���u��ˋ�0�����%����%�NP�����V��q�����s�%�6ci0�up�6�d�jh�h9�˺���(��WkG1�T��,�܈��-�q��J!�n�<hڹ��rc����&���v됻$�wY^�1��vwW�Z:)wR����6�8n�o�3��]Ʉ���@N$c�qۮ���/&n��מ97(tn�]���5=+��8���¼Y�]��]�����C�qu��S�y$�j��\�$V_*���E�W[:�����+���l1���b���E3�H3/kguۮ�d�xWn�W9���y0�t��x��,E�s璃]�����q�l�u�N�9��uָ}B�u�����T�]�TsFm��ے��4�j��y�ɲ���w�<�����[��	���������^�N7�����Ÿ�2�.S^%<�;�!�\�aS�v��i�<xŗ�cN�ϰT C���9��u�&�pp���x�
����h� 0ITs�/7�Y1��챱���!mԫ��rt�z�;�:��v�<�ov]Ǡ��;�����rc�nm�w]/]���>�Ak�^T�NM���2�x<v�\�<�s;iݟ=�Ü��k<\�Ǜ�%×&�ۑ��� P\���î�8��-��h-�)����9Ǖ^�N\s�	�|]���cn����Fy�t.�rOnz��ݡa��.�Z��m����\��1r#qK<�(Y��/	���gnW�z�e^r짶ͳ�������:󝛢�bB.xh��7>9���1<� .Z�t)���7��*�k���W�^ǳz'�m���u: �`��y��{�t�|#��n��2CD� I\cq���.A�X"Q�\���3�\�H�@�Ff�M�ԙ~�{^{PMt.�<
��ح{9���]��0.�K� �.�Uw�鞩3{ۦ��}9�^WֶҒc��d��x+~Y]^Ż7	�=�G6�)�c.YȂaC)��{�2i]���6��ȼcl]��H�죛��+s37S�Z�=�U�z>%5/f孬��@�-�M�=�o֘y�1Ǽ^?_��[=P��HQn{2P�콸�#��eG*e����uyo?M�
&YTb�:�#W�-�וL}Z'<���r��:��=�,���7���Ÿj�{}��ֽci�����OW�*TU&�XS��R�m�<3|ؾ�r��~�t ��&z
���Z�<A[l���b8޹NXr�3��x�������f�:k$�.��(�*�����-�=u����J����/['l�O*��H���#�Aӂ��>��j���U�ek��F{\�Ō�����-
�Ѯ� �6K�]�U̶�������y�Wg�՞��w>�&8<�9N������,���g�`��z��y7�,4,b 	�fOj��"���B��f�S<���Nl�z�Z�uFS�`+�n����V�u�2�6��t�tF�Ɍg�s79�	�}�-�5�}v��r��J���W�P^ 4{&�y�-N�ϽB-4�.랑vL�n߭�k�`0C�o��y��#jǧ���^]5����}�8\=~Z�� �3k��r&��HT3C+���bga�|�ϏA�M*tT��ˣ��g�����kEub�n@��#��M���Xн���o��ܩ�|�IH��c��׃=u����ۂ����s�p�7d\Il�m�O�{rȘ��Wy�@o��O�J��7�,�I#1�G���*à�6&�.��(��j��Ɣ�I2Rt�nD^h�r�IYB����	
Mfy�h+;7d�C�m\4���دd�ϛ�Ҹi)��%u�jVC撹�� �+������5���6:Q���Ź4x{��-�[�F��l7�K�Ay!Hh�ez�*�تg\�Ta����~I@�Jsv9"����3�/�F�N�.R�i��w7}�b>~O�2�&=�Y��w�o��� ��6��[��8��V���	֘|�����r��{1;iV:S����Q䒨|�`殗u�1��e{�y�u�xX3k��D���m����I3���wJ����:�S����7?��^�L�2rh^�{��ۈ#�k�h�F�2���D �	��
��� *�=[;�{��ۛ�x��Nw&�IO�i�-+��+�f�@B0j�j�jz.�׏3b��myL��m�<��9��R���������L��v�B��J�I�Z�,���I�s;��or��'��"�7ȼ.E��t�=�w�a�F��a�})��Mq;���rA$�@H8q;�8��x� ����W8�Ј��'��,j�9�*f����p����u
:����3WPǳk�1�t�풆��F�@�앱z����*Ɯ�%��ﯠ��c�8M�����nz�i��5Ó��a4��)ԥǻHs��=n�N<���'��fλ4ļpW�ybJ���E<���3��k�গ��]�u�\�v����9=(�����Ƥ�aR՜�{�N���7m�i@��Ƣݱv�����)�y�hm��7Z���rܯ+��x�a������W+�ֶsu
�[�N��?i*	��C�0�:�g�����}�S�P����Qv�^Ҽ�&��j	
� �z�����?*_���\��q���.~
c��
ѻ���n{W�g����;呸$;�f݌�����E߽e�RI	��ú�Mx���#�˽�T4`��!.�n9n7�K���>�v�0@,:tA�F�i&t�j���A�*w>ҽӬ���x|U�6EX�/,�+3�*�:"��� ^�ز��Y�7�k}�g+�ZG��*wuMڽ<�i����[��hr[�XLt�f�x�^�p�l
T�(�320^�K����|�{��\��v�Ş�ޓ=�9_OH�bɴ��������Q���IP)�ۥB�=���ެ���^'X��Q���bfɀd�g�w����և�/a���]���y�3�Me���	���#K:���k$�e�	�X�I�*ϲu*�ߖ%�;����Ȯ�J��#2+���z��e%���<��/�]�?���ӄ�V2��8D�]G�:���n�%B���צ���8����Z��}Yا�>�p j&��6��3�ka��N�[~���i'5�M�~v�n����y6RrY����,�ԡ����E��n ��-�n�x�g�Ҩ1y�J0ͱ�t��޲��u�W�
aY}"̼�c2�iEr'��V��8=�w�>������_�&��/
�X<��-JrP!���>��Πl�V�I:����C���Cjr��nɢ+��ۼ�<M��&h��[|7˦���&�o�j�Hk*�w���(W�J�J_�O�okFo�^�M�噝���ԡ�Y�p�b��|�-�g�Iλ�a�fV��=�o~���yP�6�t�ej �yu��ɮDܯ`2���Nϰ"M�`���~W��z����4� ��F�6�7tlc:[�XԷ��zg���������E�Pb��I�~8���oA���_��}&�9N��y�&���;sǚ����L��*�T�THD�Yj�7~��k���}�x{3�c�eY�=x���;��5�.N�	�:l�w����ko���1�RH�ol�]�_t�;]�.�����(�W�ZHIե�zsPD��ە�u�	b��P��rE:�H����R@�)���K4v9�F�xt�I-n�m����L�k�k�rv�vWQ��>hi��C���N�}߮�ٰ�$hT��4��ݎ� J?`�˯^�N����V��#�<J�^5�7�+�N�oY�5���=��L����!�A��N�
�n��܁���1�m{��J�O�?�c��>��NPs:y��z&i���d/��p�a���E$؀m�c����b�.����]p�yk�����w�H�n�6���@e��������2��#��T����[��A��g��
�����0ضQٗ4�e5-U1`[�]P�t��c�6ع�Y��Vnw�n�Ă`}�{)�Ä��{���7'f���v���u�ޙաz�����y�w���.d���6��ƕ4�����z�>Bwf�3Y�L���sУ����$����������񛾘����민����"l�F�J���%��g#�3��Ϡ-�:ڊ�ɲ�!���yZ�c�1��Ǵ;�陡��u����\�)����/���`f��^J7��,�Ҋ�K������L��L��9C^���s�Ҽ�{X��Y��ɯ*&��(���>WK��o��:JΊ����N��j����d甧���$kw<T7��xK�㧙L|�
m�����݉W�b»����u�y�~�z/o�3����:o�`�"���P�����`{����P�i�B@�{;���u�7��z�����V�s� H;]�=З����])�F�C�g�����<�B��F��6ve�ҏ�����a1�J���]����̎R��F�JZ�=�3y��N�2�"+o'�L��<�=�T�f?6����P�WE����>�yU��ɗ�0N��U�(]������ o&�	�>�
dƉ��0wgm�Uu�4C^Kf@�c���/,�������ԛ{˜K���͆�h�QG�j��2}LN��������+Ќ�� ��X�p2Ʃ��_u+�����&1F�YGF�x�f_b�7�I�(��f]^�Y�yQV[u�;�pփTM �0
�eq�E��%Oh箯W�Ύ�q���۠��96��$�� �cg-�v�%�h���>��6����I����и��y�!�9�oqɘ9��[:�;Ν�*ܻK��5"s.Q�g.����=y���@n��zx�{)&�u��G�A�ݬ�f�.�86�^y�W�d�c�I8e�vv�H�.9w�����t�&ڢU�D ) 2� ���]� m�ɋö�=�����!������D�%+$�I��n���#s�m.��PXXU�9=׾��O΍�rd~מ{�ן�R�=��M^:O/b��C�*��N�i�e����.�͍h�G���ƴzϸ��56�]�h )�g���M���t�
he��pV
n:�%8�sj�$N��+{���X�<��w���{3� =�%__:΀�R{�ڹ]hQ�����Zu�-fĘݯ~1ﳽ��lW�M����{9J��d]�;н��p����}D.� �E�DH`���nZ��s�;��ۅ�>4:yF�Y|QS����p��ͫ�0?^�[�1�{O�)���v�Vש��(���o�q�%�u0��eؑ����6	�������]��������ewx,�Fp��`��A6�7o6�{��yE���l/-��2���kf�=�} �y�|�ȶ�WvR4P�W^R�����V��2Vv��Y�O^�X����`e���-�/!�:A��̻��x#��i9��sm�̗eqE���l�:缜f�uu&
MI'���0VQ��n�離AY�zWm�ϙ��YyE����s⫺����4��G��ݗ�ⱂ, ٹq9$�����$��dãy���'|ʜ��֦��|#�~�z���ٶ3���Mm,ݱ/�����L��x�P�9�:�X����%�}��PC�r���oF�	��ŢgG�]l��?���<���L+<��7ۖ��^�O9�͎�2��}Kى��#����.:��z��[�жT�QT��	+p�7�`�6.������zOo��.{�:@��+1K�{�Ю��䏓��-ƻ����l�H6�F`�wΕ��h��s�hl�>�7��L�w����j5��7�e-������A��e�Y���K����ם=F�@����Q���.��k¸�����U�����������v�;���:��-�^׬Qs׮(
�D��@�Ѥ��5ڷ����f�2K��/��WY���F��o09��P�!���XP+�e�2J�!R�bCn�t�%GjХ�v�a�m�� �Ӹ;�rmmeZE�q�����-��v��[Ñ�j�(�OF
���&{}�4,�ͷM]���w]I��J>N̐��컬7w|5W��� ��&��iԸ�Bd4�
B0�3����L=5��=�l�g7�z��{҇玕�i<>�Դ�N�d�`�a�J��"��@�U7H�c����M�]R��G���>Hg(=5.ĮdT�s0��z���H`w�Bʱ��P��L����F�3޷�~f��t˥NLuv)�h]y�}��Y^C�[���{K�!�'�]S(�3C���WuR6�Z À������ܘ��gg�iLn�<����.�M�a��9,ٸz���y9ѫj�Y�_ąY��&�)Pn։�<�?JY��w��Ix@*��Q���ݾ�]�W�Pn���e��nۤ�u�c��'��(N�ҽ˛_�B���^�o�ѷ�s�嗮���e���@{䁢L�1x��w��������{���ww{�����w�����{��������{�{��������������������w�������{�������{���{���������q�w{����w����{������w���{�������{������������w��=���w{������������ww{�����{���������ww���{�������{������{�����w{��W�U_U}��s�e5�uD�peam� ?�s�m���� 1���(� �            (  �                               @                  <@  ,`��� @#귰�� =4M h`v��(�;44 �  P@v 4 `.���� @�  :
 ;a��� 4���:   ��@N�
��@{�x �l(4=�ʽi.�8lۭ�f��%(���pw9��(���6�6��]tt�R�ݭ�p�ё[��6m��  0   eu������,˭��۶�d���u��b��S����M���	�lҝ�[m8US{'{p����b6Q����iJ�t� $�ÎKd�(     jѻ3�v�K���v��ivʃ[��.܆�v݌���:î��F��n�ڲ�6��N��wwU�N�u;���Ғ��핡��iZn�&�  �   1����S�ƍbGm
��b�֎�n���4]wls �s�WRJ�(5]���v``��֝�0�`�"  � � v�=���C��0``퓀a��T��M �iGCZ�8飱��sp:�M4$�SL�( ��  0   6ݸh 1�(h-�5��]����( 3��kAN�l+��Wpq�6�j4f��  �    wkT���ݣvp`��tkM0	���N���.����Zh5��@ P     �S�
 �`�$
h5����h ���]��C  �`���   0    l
�t��0 ]��� ���� �P )ѠA�  (@� ���Bb�J 4    ��@��S@5=L� !��di���CS&�!�hh�=���T�%T�# � ��~�&���4h���h I�H�     �y�W�s���ߦm�w暻�ۺxk�3mf��Z�O2�����=�;�����H@ ���<`P�7%BE
����O�u?yT���y��Z�@q�9M0@O�mj*�ʄ̩ݕM����$��B�j5$�$!�ԓBV��$��� V�	1 *I&!%d���2L@H1$12�@�B��T���T�I+$*5�
�!� �A@&$d$Ԓ�$5$�$&���� I�H�@&!	RH �	V�E�P��%F�i%f(1��BJ�*I!1
�	R�$+Y$
��T+B�B�T� @�
Œ@��@1���$���� Ą$�²HLHJ��c! J�bL` ���+
�Ą*���%a
�Y!�&!�J�˖�kR�I�
!\m����m���-E	�Y
�P��I%bE�*ZaR��V�Dk��c�ԒI��H� ���R ,j��IY*I+*BJ��	Y!X�K��������C�g�s�J��(�F�����Cv��a�56��
�+��G��*��J��[�b��۬j���;��x/�u��eWiʎ�pO9���kv��l�wz�U�d�g�՛7�ه���4��ZxP]1|ԩ[|V�˥�,�e��.��s�t�B��af�f�p4s�r9��bn>��O&vj}�B��*T�h?
#�~A���f��UZ�)x+4:�+s(=�Gc%���}/,����`��fT��sh�ڇl�2�I�E�+.����ɚ��j�6�U��Qѫ%jBU��5�3v���٢h*��jw	�B���r�V��{��""3�����-���2����X��7Z$�cV�Wv��]c�@��)�4��A`�
���׺`W��]���J�����d������X�vop��%GLm��n�j-#WOq$,_�-c��WuR\��m՟��j�wN�0̇N��IO�f�$
��{
ʘ*�)Ql��{T�J�Y�շ�yys)VE�^�i��z�݈�h�,�!Y����[��֩YE��9��!�si.2ƈ;��=r��@��Դ"��-Ţ��@8vj��M�M�}�,ᗧ+l��b��f��l2k6Q�J݋��]+����.�S�˱��ko��pmkѝS�Ssm=�vL�p�6��a�e;�AcL�Q�4�i�ML����3"��udx�Nz�\���!���*�='U-�5B�|�^�0t9W,�ՙ�Nڨ�-8��m�8U�U)Szt�xꄆ%�X�F��_LP�*1QS͸䴛&�R�B��]�R ����mP�ܭ���sqlx������Y�k-�%7�R�%�"�WW�^�͘��m%�Yt�]���o4e�����ec�g�˷�E�����J�wL^4��;x�3n7�;�$�R^[8��uf��[�0ѥU���rc.a�v�^ͬz�$��"ĺr'���Xt`���&ˬ�C��+
��;�)@�[��k&i�
+���fI�uq-��L3��,B�ڢ�7��`�o��fV�g0A�3h��`Ѓ�<H��nf�����I�-.����땖��"��v�<U�n^�����2b���M˽b���i�.6��b�w�T@��{�"M��5�#$6
�Q
;�����GB�:tR6��hZ�� ��C��;�����#w�SH�t��Ke�*�"�P+�놣�eU��Y��e�8�m����������Ā�#d9�ԕz�*���Дcx�7�Sh��q�SR�͜Ȥ�Q��&��.Ky���&����/i齻R�*}6�җDB�Л[U�0�╎f@�	�+�4�J�FrQi��&*�����H�nm��>�f�78}V���
0PgL�p���p�$��m���Y�<�vZwr��o]�ԡ7~�q���J�5O(��ɚ%�Zڬ��skk�{�I������Z6Ui#�+hR���0`�A|�0s�������,FQ,�T:�f�J
�!���ܦn��нb^�y�ta��]�n	{���d6������#T@틤h�w�`�0���2�%m�K�H7���3o7Uv�e
��dR�&������p�=��I��$�6���rUa��b3X�A�u�.�Gj*&�cQ�gn�ed�kr���/Mύ�Q����#-��]+�aDMڣgF���8fb6/ɵ�`j�9n�U���h��n�KZ��)�O4�XE�Ȕ#ֽ���nĨv_Ɲ�.�9��x`E8x`�GE472�F����2���A��@�Z�Ul���k�w���-l��(`�I��DZ��Ɵ�eM�n�ѳ7/�����;�͟�Ƴ)�Dm#	Grݱk�2�B�_֪����R]c۽3B	K��UZU��#6��B-�T-m��w2�9��U��US�X����$�S�m�w	EaN�\+��ۉ��f�k	����bs��)�W�7�u��d�3�It�6..���u�YJf���cV����X�&�݃����f,�X�9����ӛU�Y-��+f����j�����9}���Ҿ��4����KtC�5Q���Z�6R/RM�۪Y�E�m��_oX�A���i �A��}��S�O��!�}vn�3{n�X�y�1<���ܝ��
��u�{��=Ֆ8j�5ۗ��)�'��^�k�x]���.�L�Fa�@�4��X{�T�vƾ�φ�Υ�\*��r����&��s���[9c�}�?d��R:�(�Yv�����)M�ڹ!W�|7|�"�v\�XN=�+߬���V����.�f��Ĥ��S	k��F��!��ˣuX)��kl�ܰ�M/M��u� 3iZs%w�J�gsJ"u�`�5�K��?���Je�I������<��W��S�Rj�6�`��VK�P�ok�k{����6��;y���C�����:S+̦���n��*a��?+Q��m�RIY|�y�D;+�ٍd�h��pl�m��dK��Tp�W����م[[{^$+t�U���2rQ�"
�Y����<��W1�p�c&8%*�w��P]��ʃ�1ͱ�!Ō�Z�͎,*��
B��%�/0�NT;�ii�9�ы0��d:l�&�ܲ�]�^itlZ�h�W4�{ZN�L��E[EP���7A��yT.��Xfm��k~��mc�Y�Wڡ�ɘ�Xu����K[S)n�e�
�Y�{��%�a��W�C�Ī�hOv�)N<a��:���r3��ܝ)nRe�2���ƶ����Z?Y�v�}J���(i7���ViZ�uKʾ�a��W3��PT�Yܮ�Q�X�}i�9^hB��k���@]IU\�c���PyW���j�ڭ7�$Iecɹ�V�6FwDi۱���t�u���̪�Ҽ����|-9��;���Y#l�0����H)��_C�l�5>���_UԟQT�;n��h|Hd��%p��~��B�HX�.�� "G�.�{3�v��5�b�+Զ����tn�����TR�YP=_Qq2'�]|&�)�ThNb�__eú%}ݛ�l@�ޮ���9���Ԏ��:Щd�B�n��[�O-�eguX������Ȯ���5�1F�Ì薭�ƏD�X�,r�q-��W�Wݽ���eE��k�yU�C{'#[��O�̣�[�e���W:���y�J�XJ��y�$-db�cXY�u8���G�FJ�K �^��Ȯ�0(��j��F�ݼ�Բ�A���"�������7>��ׄ��P9�X�����3�Lõ��ӵYY�z4���W`R6���P'0����b�η���8b
����+^����da�x֡J��������9�H�ۗ�Ř���^��� �VwUb)���+HB�%@�j�F�Z�e)RT��AH,R*��dR
AH),DQE�E

Ak
ŁR (��H�$RAAa(dR�J�ʬ���Z ��ł��ȡD+ԢV�+��	D� *�� ŊE �11IK)b�A�("(���¡P�,QR
 ��PF1��dE`� �AEDP�Ŋ(�1DEAb��R*V,@R
AH)�"��$�Y-�A,X�dQ�1�#"�U��RVK*�eAEUF �DDPX*F,PZ0*-bJ�X�����B�Z��X)+*AH,U�
�@D�hQ��� ���RUX�)YAV*�kAQ+
 �,X���Ōb�[a�XJ�UUV��BP� Eaa-��P��
�[B�#A�`Ȁ4iU()Y	D�"b�����P�l�[�
 ���d�E��E���VZAe��Q"�K(��U��E�AHVi
�"�V�UQam �(�*AH)
�R
Ab%��-!l	Y!�,��R
AH) ��$����R
AH) � ���R
AH)c
�RTiH)+*AH) ���X��� ��JH,�+"U,�����*AH) ��$��0�Y*A�k-JD��-KA-�@�l+J�)mm#h�*J%aP�(�� ���V����H(�+P�Qb�Vȵ�����RQPB( $����롆}���R��͠��j�i���T ��*�Lͱ�"r��޻zM��kն�m�LVkKR�uf,h*�CMZ
�ͬ�Y��ѰK��zS��ҟd]m�d^�\wO�Ї��CʟAݭ�̊2�=����_lѵ�T���v�ŢXzuc90@˴hU�����:���0���(��[i��[���<��Ը���|�,d�w����h\�g���9G��D*�c�����s��vd�Z6��U�_e;a��J�	��w��ЕYʪ*1�w"l]Ҭ[gb�f��5uu�-��X��J��b���<�*�ՃG1�f�l�V��Kj�+VۄQN���xQ��묩��V��g/M�˭�f�ϖ���*�88���+7wp�,;PQe�0˻2�
�76�0�H-��U֐�Puan��X�miį1j��U��RWB�A�刭��V��#IhRf�lV����B��zqe�wW��֌ɭ�S�t�v�)±(�1ܸj�м�O�}Oq�ѧ���^AZ�ُ�9w��,G�k3%m|���;�a�H����wRu�0VU$T�[jұ,�!�����B���ɵA�wa<��eaN�h]���fё����T�$塹����ٵ0�:�5��&�eS��C20��n�K;jiUF��c���kت�w`ā�eV;n�5H��&�њln#uw2��a
S��Q�&��U�d��J��f��yˈ�?]B�=A�N��3R�T��Ν��ՙ�y��^��U�X�v2�3�[d"��Gl֗�� O�V"�w�j����{�k��͂�q��0��M~��Z����ܭ�x���f����e��#7!�F%F��̕r�K�y/m�.)w��
�9bf�c�h����Kȶ-�ɡ�4㒲�)�!#�Csv�����0l��ܪ��H�b�t�S6�Z~*P�ܖ� 76��;�(1��e�iX:�Y�:�G/
�����.|�!ZۛJ��ڦAZ�f*v��K�v���!�X��L��k8�V�𙪩7)�}�Ϧ�Y��+�wϳ���* ��/AI�ϕe����Ale!�Һ�[�w���R&� �.inom�m�c��U�6�c��HZҌ�hv�&�a�ΩEi�zD��++FA������=��q�[�c7~�C���D�Z�d�|��)fTVm����/3�oDe���Jۻ�WA%d]ӗ�k�6i˴֡�1Xy)�P��8ze�Z���χU?����uim;�o��n�X5j\���OGU�J��eܼ�;:��F�rjA<���Q�+�W1�]���W�R��w��I����T2�R�q�+j���s�/�ӕU�/��P�gCw&;��4�J������*�8r;,�w����&=�a�B��*X�V�ݽ��F��c3,j�Py��Mɕ��:�s���R���YHȝUmJwLW�Y��)'�S��Fe�����E�ec�7$�����6"�exZ�z�)u*��dۨ�j�:ch5�6Jj���}ݰ�X�oe�6:�a
�'�f�<&�]6�w[}4��s��32�r�Y������=rۧܩJ�SKq�S�r���b�}�z�CX��K��ќ������g8��_��l%�����DDcl�aW��)V��	�S*�j_n���ij��P*�]�-ʑ��������*�*T�j������Ui
:;v����p���r�KUT����v��Ӑ4��p�`*���[j0��KWUUUUR�R�UU@UU*�UJ��.��Ti�@l��%ZU��t���jj�UV�[6����4� p� s��d3�F�j���j�їbg8�F �NԶ�N.�B�.{���h �[K�e+j�3������+x���I�2I�5AQ��p'�`:^��Qʊ���v�7��y6t�{��u��&.`N�-��f`���Y6N��q��u�_Ysݙa����pu�S��#�����Nۭ��ohw)cs�s���@{Gm��;��T3��[�T��D����Ep�7\:����l���q��M�1��7��zq��Fy�S�g���۩���n4X㶻�uy��k��R]�aS��k���S��Q��۲pp�jrt�G`1�[��^�=��c�]��pd�u]v}Z���8��܃����j����r�D-�l�a��z�������t�m�ah�=�뇋]c�'e7;"Bb���Sm�wmsn#v�g��d�S��i��N���=����s���0Ec..�6�Wl\�y��[����u��͚1���>�D��v�i{!��S�b����һu��c���^y�7	��N*��W�b�<���*Dky���b^��g���l�����'[�=�����=l-�[���E�=�Ѩ���9H�u��9�y���ӹ���\�R��U����])z{#<{n�^6�9g�NX�Y7=���bf�D�9S�cM�w��ڧ�����sV�P���⻱�d���7I6�&���[RV�Lt���L�\�"�m�i,c��.�����kF�{4��F�ە�) S��tc[k�LZ����7lv�����8�sѩ�z���:�/�5�;�2t6�fz8�\vz]�;�q�w@@�k>���������a�6.�٠��\=]��L�����q���=��+�{o9��!��&��݂}�7:��=�� )����tѝ��=���n��d�p���=��h,h��='jG���h[��k�V{v��P�s�{!ݵ�� my�˹˭jR�����۶�d0�v�[\������7=ͽ#<���e=v�:�K�.�-�2���yH9�vV���ʦ���NKt��=�$�6��ۻjn�N���H��J��^��ϐ�ή�y��]��HhǢz0�ݻ#�����zpc�8nlcuݎ����Fd������Cؖ���9�5�W���E�ˑ��<��e���,�d���ίGvq;f��*=�:�U�vj^OCy\��θ�A���rx��T�9�f�m�=g����]�st�wkn�F`��ۥh��h�]��T��]-���p�����ıF۴Q���4�������q�q�!�UPU�A��n2k�Ns[�;	��G]fw$۱�ַi�5�{F݀���^d5�q�Ͱ�ۍ�7B���l���n0hD뭰�X;m��@���n�s�#su�떘��%q�jD����:�1����3���.��]nw!n�vE��tޓ������7{g�ip3�ЧNX�K]sэ۷m�հ�wc���;��K`���tu�8�k�M�n�x@�u0��t��)'�����neU�7�g�%؈^p-֞y+�^���Ń�-c���<C�m�Oi���iwn
�b��jy�s�r2�<�	nB�/h����	۶��+�E�k�g��;�Wn,�`�'��6�>�Y=��v-m���^ź�h��x;��-.��#�t�!�C��6�v��Ϝnwv���m��;i��v�M�6�n�lqΎ�c�|�ع�K�%�wC��ܕ�#%�AZ�v��j�tA��s�/\V��Gk�+ȼ�'����gv�N`O]m������W������v|���.�e��ml��pu�К!n�k���l�VT��6C���,������x�n���7>v��d���'��tqO@��%9O'���n\�npx����7ulsGX�v��ٴb��8�}�=!�q�{r��������V���[�Wg]R<#(t���m�y����֛b�e��.xn�N�cZt�&,p���a۬G\�Z ��p6�K��z�նGs�:�j7vN��Y�ӭ�PĜ�����qq�n�NE�u�krT���{��[w4󋎦�FVݷ������R����^�@�^����ɳ�9�m˒r�Y��]����q��;��{���o78�o+��F��I��C�֛c]�1۝[�l�ni;hϫV��q׎x��ck
m�n�h}�ݻ2m�r���E���h��9�]q�@��u��g����v��]��]e�Tq�cTg���x{(v��F���m���8�\�f���b�ۜY[����\n.�L�ݻ@�S��;..�8u�i!���Y�mn���3�{"v�]kp�$q��q��m�.m%������뮸"�E�0�cЅt�����O�e��Nɷ9�+uX�]g%���8�8�1�Q��_s�M��l&��}��wn_Wk@�5�u�k��њ;-��Q5̖�v�fmr�pZ`f�^�����S͎�3郗z�����:,q�/���Q �Xy��́;nD�ӎvN�]��m���y�ˁ�Ƒ{z�*�#,ۨQ8�u�5�Vn�6�E��W��C����C7d.[��v9ؔm=�X���V�.�v��N�5�O\Z�8K88�0��Gj���E��cp�vؽ1�pǭ�n8��F��ү6ƥ�CM�n�C�\�ϙ\j��G�]لŸ!ú��jR�qǎݘ�t�]��o'�n^v��[Wo`��ok�գv�ƽ�v�N�i�z�N�J]Į4�3kQ�F#�-��:�wr�bV�v�ʺ��{>yݶ�6��P��K�m�=�.�n�5��ݲ��R(=��u�ݩú�	��l��{Yպgz@��5*vѭ����/WE��t���m��:�ѵ��7U�T%�N{In��S���;�ݧ`���=�y�	uƎ�si�cch�Q7dh��ǳ��F�wc�`#l�c�ς{	�G����v��F�\�x��`���Uu����OPnV}��x����|c��\�ͥ�H�&����X�Y��'�;�nւ�'���=���;/toX�6%Ʈ��9NŽ��+��\�]���O<�˷o8#�7^���������UUU*�T�*j]R�dTRZ�������YZ���j���Z���V����
Y�[;*mH6����tUU	)(F�Z���N�+UJ��UWUUUUUUUUUUUUUUUUR�T�UUUUUUUUUJ:����UUJ9��T�UU]UU6��(��
��j�������Z�j55UUUUUUUUU*�R�+UJ�*�UT�/�UUUUUEJ�UUUUu*�UUU��[����Z��(�������yZ�mUTYZ��Uғ<	5UU[U�cv}[=��U�VғUM��HU'���������enWb�����UU�2j��-�Un�e$��(7j�*��s��f��aj�V���-R�UJ�S�E���[�t9g sK�z�:�+J�j�����W]lk��g�P�:��m%���x ��;U�)`��P+U���:�]��Bj������ꪪ.���UUUUUUUUUUUUUUUUT�UU-�"j�y���i�ሢ��SYFp%F�UUUUUU]UUE�USj����������ꪫT�WUUUѩ��UUUU�j����ꃊX*mU�����T�WUUU�USj�����MUuUU]UU6��(��T�WUUU�USj�����MUuUU]UU6��(��T�WUUU�USj�����MUuUU]UU6��(��T�WV����U�S�1;6�U�U�	��k��W�U�J�QUV��������YF��R�+UUՂ�0r�*�t�ͪ��4�i���������UEUj��ꪪ���mUTQW�z��j����ꪩ�'h�@9�CC k;��S�R2��!&M�[&Y�ꪶ���������-UUUUUU�U+m���D�N�v`��iM6�e�������Z�����(��1�qT�UUT�UUWUUJ��C����UT��R��9�j� ���	���!ԫ*�ێjF���U|����������U�4�UUT�*�Ίڠi
@Z�
Z�����0�J��J�MUN�*VV�S"�*�T��UJ�UUUUT�Ԫ�U\T�UW����%T&��#l�1jq�cF����j�������&������T�]s�*�HMU�P�9����5m�fBI=�Ɯ�m[h�G[fEF�ݢ��CvA�)tk�g�	e`��:�\6*��U;��bU�mlv���UUA�UuUUUUPUT�5lmF�T<V3�<Ln�k��Z���,M"��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_U_*��������������������j��M��(�TUUU�V�UUUUUUUUUUUUT�UUUUUUUUQ����T�U�UJ��UUUUUUPR�+T�KUT�R�N���Zv�;��k�򪔖�������j��j�Ij������"%�����Z�������������������|��~UUUUUUUUUUUUUUUUUUUUUUUUUUUUUT�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU[UUUUT��UUJ�UUUUUUUUUUUUUUUUUUT��UUUUUUUPUUUUT�UUU�UUUUUUUUUUUUUUUUUUUUo�>|�*�UU\��[UC���UUmSj�2T��TR�UUPUUUUUUUUUUR��UUUUR�UUUV�R�]��]��otP�*�@q��P���q��8b��ƪ����u�����;�����o�'��ד7o�n㦍��%U������c�b���5UUUUU֩vV��j�j�YZU����Z����&ӦB��F�֖�gt`�w7�`����u*�=r֪������GgjW����*���j��7d������UUUU�j����ꪫc]4njUmUV4�������V��k�kh��j������4�T�J�����F��-Sj�X�U�$S(�J�UT��R�ԭ��V��g��*eڴ�5հQT���LWJ-UUUUUUUUUUUUUUUUUUUUUUT�UUUT�EZ����L�UUR��Uz���U�Z�������������������ej�����jU����T(%VBj��U�����D�`���J�2���! ���$����@I"�E�!	 �	'��N���j��n�w5�wsW��Ӎ\c��-^�b���M��Rq@������h�H cUUUUJ�J�*�J�UUU U;��C��( �cg� ���?��o��⺎��L��$��YR�5T�lʻ��{/|�t����˞ם;o�9���ᒑ�����.
u�!��Q=m.Y(�fT�q�c��@��:�X0���{�u�jج�$K�R;Z�P��`�0B�U�~��>�í��/i���G��Y�BD�0j�kQ���`�\=��r�������Û4S�ҋ&RcR'%�(�5���G(�Z]�/WpZF�Ey��^�l
V�m��Up��#���DT8E{��W�����%�)�����ђ�wl��$�0H��AI������ĝs��_��1�rt�=:���Z������)>v$n���z��;��>�=StS��|�x㋩����ϟ��Q
��X�$e\��^hn�l?`o��#�[��$���*��궱~��{�@��ԭB��)*�� ��C�t%W�����R�yx6�EH��L�'�J��w�*�m����)1�)��(K�8�Q������oZj�`B.@�u��v�c�sv�r���&���PM��<�2J�_�8o�[�3��CS��&S�<+�I�Q�a�4���N�૆�h��Ua�C=7�h�W�_x�s_��l[��X7�f.����y�����άx�#u��XJ��<H�PKh��X:
0��Q!ӱ��8�N�x�(�Gs��L!�GZ�i}A��ol\j[&_�Ʋ��:�:��w]��`�+&m�1l�N�.ݫ�+V�����Nͷ]p��K����Άݨ��T�j�k�Ņ⋒*�ۭ;��	������=�g��Ms������I5'on�t�RS2Y5�ı��+��&��ɲ4����
aL0WN~��Y�:����'����}�k.�\�wBt&"�`�����ry�7�ܫ�b�1g�@��.'՗����p�:'֩�֩� �%�S��SJ���>{n�{�/ۏ�Ge�q��-�V��ϓka���;�t���}�z���z-D{[a%���-]��C(_�h-�p�х�����D�~�z�5���1���3��Dx�L�2��eU%��a�X�% ��RX"]�e�D�0!m#�����B�����f́Z6v1���(MZY'AD�P����n+�֏����_��$�]jt8�Vں�������)7� �q(��"NF�r�n�b�Z��栴�
�`�Fi�S7�'��Fҋ��IxW�t�q?j��Q�Ǹ%��U
+���(�I���[ �+���%#I�Lf������Ⱥ�*�g;=z�q�*[�e%.��U�Kt�WU�!�#ЀGL�A5=���_�t�]�t
�WٸN���e;˻�Kl����hE�����J	z�%-3���jj�\��͚C���-�dHB��XLF��2.+��[,�4��Q�9���w4���&*!��4E��P�D���!�G�^�4���Z���L�;�kE% ��n	&G��,��`��R�*!$*�rn��r������2�E�׆uku��w��U�(�jKE�YT����p��U�Չ�=y%��mu}���!9i�R�l����Ud�3�E�
�`��!��#C��Y#�/�!Jֶ�M؍;Β�\�8��R���:`��J�w�ja3)h�QO�5�b��ϫ�=պN���?r�H
�A�$�Ԯ-���u ձ���/+$�z��ݕ>���]�H)_!����}i핡�����L�5�[8vL���ؤ����ӂ��� �7R�.�iAq���n�S��ͦ�ъ��C�%w�W*��6]��j}�Ï�BY���l��H�'Y�f�-��*��j���\�����GN�K:�������$�P�[ �m�[�QX}�>	��IuD�f�y�rG�?T�=<�^,��������x��l�k�@x�)l-��u���� ��V
�$p�Ww&#b�;HǦs���%.)&FL��������i�n$�Ts�v������iPu�TK>�M�����d.���#�&bW��UA�\��qA� V�w{�j��9Qκ.�qjYOk����Z��;)�3x��8�ƺJ�8P�5�G�DT�,�Ğ�'h���iv�y�z��%i>�S�' ��}n"B���zf_<�Mkum��ߪ��k
���_Ĳ��q���ګ�M�]ˎ9$��������~j�����@L�4��)�U���f�f�z��h!$��K�!��Y.,-�z���ϢƇ%���I�kz2��΋Р0}K���ԓ�<4�ϣ���h�qq魥���:��Z0j��˫�:{+��U �|�~��&i=	m+�Z�r�E��Nw����S`�¶����5yT���m��Fob�𠒳@��H���F�W�i#����t�q�ۼd?�]�ۨ�fR3T�X����ˊ���\#`��Q�KC���Tf?��KW�
�oI�K����ߴ�Q�"�Z^`��/��w;F^M]v���+�u��h�-�������!�H`n�;��Ԧ�_a�:�Wփ9���:���9���֣7���F(+S�݊V0� rA�|naI��+��P����;�M��;g3\����(73v��A��|���+�NF����(��Ԝ5�|
l�
�pUe���c1��R�b��Ҷ�!���K>�T���L*Q���w��sϕՂ>=��ۜgko�'djU������������v��U6�������`�ہ	��vD^���O+UUUUU�[:*�
����)�_�o��δg�$��ݜ�Ҥқ_�D�	W���֤T9m$/��Ov:�g��#� �����|���^����:��)�{�i�����&0E"��2��:��PU�5��X��[&;*�$�G��vT�Wv�.�_Y	�Ē�h�aK_{��Kon
+ڂ���/Z�u�]Ǩ�4�O��i�_��0k,[%��1�V�~���a��|R�o��$5忎��w����T/��o�&��TD�i���\���h��G
�}Uԍ�m�5�̂�x~���7��c,��%�:�_d-C���KWm/m�W���1G���9ha���.���T���a�m��G
���L_�z��+�Tk}C���B�ډM�ٛ�������-�0Z���&ϹW.��"�!����{_b�O��"�>��� K]�$��[-�6����Ƣ*�\BݗAIuuvg`�Y�RTӺ����!:��V�YD�m-hW��j�5q���D*�H��Z])ǭ6ؗBl2���X�uYr�]�L�Q�`�TZD*���]�m�b���*�dgz�j'Z��m����h������������B��6�a9YlYܧ8�����>�����JL]��qЀt�m`���q�G'��;nKqn�ve5�ۑ�q��1f�r��ql�gGã=����{����8봀.���<8i�g3]!����6�JI\�j&��n	�u���G5�h�٭^zsp��|wΞ�?������ձ�B[{�2)`�-?U� (������eLn�ނAA�������^a�Sěa��䄂/{�{XR�	I I�Yڲ=�=I��-�a-�=�zme2��ݴ`&�皕��/y�JE�7�$��5���D�Q�$#���eZX���Oq�C�*.���^�d�Bsv�\Z4c�wk�W��yȏ�6.+�$�%�3Ї�+�h�|��T�T"1f�mˍ�Z�qQ[}�$wv��\+�/��tŉgB�hB�0��C��(�ѯ����l��p^x\�:V<>e�2��&���+!��8+j2q��Pɩ��|���]:"z@LH��%4�h說ک���o������n%{�D[ri�󦏈M'��n㔞�s�L�[-o��yGd#_](Q��|"=�� ��$ʱ�2K�ʢFԻ#.�V�B'����C�0��6�j�s����G��tx`j�s$_A$^���d�dp템=�V�>)a�7k��-<N�N��^2��ȍ��N=Ҵ�s��Sr��;5�o�*�$Q�n�[|H+�!�)M7c���]sJt�l�;�m�Z���ʍĞ�m00�Qk^�*�����6ηi�uս�*C
H�Z{������"�X�����s�,��֏1�����n��.�l��ms"�1�&i���')-����j��m�m�!�4=A�	˩��\�'�%kޙ2�3��h���(�J�965�����}bP5#�q��"�q���c����x�ed48Z9d�yH�0(a���q�ۄ�$Q�[mA��1�ޡ�a�)+m#�r�]2e/4/	�C����I#������L�T�����d8��/�ȕ,7�%E nݞ�8PLmu�-B=���e�ю,%�/���i�4^*�=��u�K�͍�1@[��6�L{eUj��]�&��[��0x��IK�":���E�x������+d���!�Y�)崆ECn������6���&�����>2I��X������X��[�M��Vo\�L��M�^m��NHbP$K�A'Ğ��s��&M�������� �ZL���Ӕs�'|����j�g�@�]��������7���;�����N�s���Z��}�����0����u�q�R�V�)����yv�lMsJuK�b�W.> �Ѵ����t���yRz���^�:�4nu�.Upi��1��a���rF�v��O����v�ϙ{��]���jͲaNP���4���J��J!*m�Inb$4�j�..I{���:	����i6���i��B��z�G�ܙS�p0ZB�m3��E��^�j������|�۾�3j{`�3��6{��T�u�L���S�))�B�4ku��m��Qƌ����zǔ�V�hjp_S�09��ͧ�u�k���ۤ.q�b�X��6���v�i&�nQ+ۿOP��![wƘ�`F�FV����LG�Ht�l�	�����c�`��ꝉ�rO�q�DB���}�** �i��X�6lӧ�iЮw|�9h<��|��sդ{i]����KˁE�R}���	(��8jBZ�٦i�匿)}
-#���SȾ;��Z���$M�422?Z��Wg{�5
G��"آϞ\w�{H�WN�<��R�=��K5ڋ�����l��|g�VR�ŜT��<^���mA�[rG$�I$J�u=%���Ƞ��uuuUU]z55Z�nm�U+B����p���
�����$�5J��UUU@HJ�
�8ôX������:j4���O�>�+ש��Y�h������g�q1`��e�I�/�&�h��/��o,=�T!;㬧Ff��22�pZD�ux?C���E��p(����(A�+G=~u�R�7a�#�~�mb��f��6V����U��=Ǚ���ɞMս��)�l��������(�%J��n!gOr�	�����Bq<�qZ�eb�$.�1�h�q��Xٕa����uv�h\R�c/'���*��TM��t햼8'�q��ci��ަ!)BZ��6Y����y�kn�0�ޱ��.c˫�D�Y�t!5�Զ����H^4�{���]�S��N���a�sd�$r��7����ͯ�����3�Q蕕S&�R��v���ds�����.�,��#�y�����1�����l�{=��wϹJO4�!��$n���yk,�#7�=�%>+q��z�L���rA�`P���rH�-�"P�$�?yWKڻ���Z	,B�y$P�#DcX2���_ۜ�XPf���9�w��>��7*�iҭ̦��)�
���J:���~1-U�n�F%�J�n��v"�Ѭ����N�Z���N��d�1N��,�U������W����$��e���UA9D�5�񂵽˷cnf�b^�5ą�s��8��r��ݔ����Ƈ\���mv$��v;85��]<��;X�;@/��۳��c�[���:`���<�5��G;Gr��*�;�χ�QR�������4O0��	�^�.lk��n��S��w%���lP�Z���{���� g}����M�fM0��
@�v�����4�U_N��aP=
�N���$��5(ڀ��p`��[�ʄ��ƭ	C��/Ή�ۭ���(�OI����G�'{/�}��J�i�ӵ�OV��B.����quh��}|��R�{�:�zl�m}�ж��0e?��He����{��WV��]P3����H��7��(�	7�J.�mB��j��p�k��U%�4b_3�W�}�a��5�қp(�A�z<��3�k��:��ƫ���W�̽�6�'{}�(:���MѺ�ҩfہE�x`{�m�ry
m{�0[�"N���|�'/��)R��e"zP,/gE���&v�?��rL���!�`��%��*���Ѵ����GW���VR�D��L>�
��1��5q�2uIK��b�i�����@�cVo
�[�R���a��m��	����[����E�ZdC҆�e�f����	?���
�Q��^��|��?o��[�k�oNȷ=�:�WS��
H��,�ZL=��7a2��{���/,�pS{"�÷��G
��]�۴�'}%C��yW��|ʠ�֯��[��N� �!��r[��ַ���K@�GYD��w�=�f�2	�V%ï�gE���VI���=H�/#NIpժ��^4��T|m����Ք�����`�Z�ȗc��h���:oWt��l��"_���=n�d��� TFj�!��|����ݴ1 ���g�t�y�!�F���g��)T�x�˶��:���$���v�r�ua�L��X��_�Jb��ӹ����͕��ľ���v���fi��,a��]�x�y9O���	���e,��y���v>�فU��C�O�DYIYh��@3�4ᙏ
�������K�}lC�-M�+/��^�#��܀I ��C���My����<��y����j�LAdm��D�Fi�F�h��0�:�{����h{ѐ�t���EԒ\�!md�s�}m��Т;3cO���>4�Z��g
�L!gR&��*о�j�r�x��6_�ď�ʓ�Z��gMr��/y
kHG� ��H$d��&��A"�3i�1dqo�8M/�"z�?_#��8n<v���Gui��^��gi�t(�êP�Q|�=>�gTb��=3FZtr�n��I),�4��9���i��t2eJP�0
A4)�+RFG/]c\�+*�N��F+hz�3��i���1j��j��E������S��:y��M�B\N7����i2fz۞�l'k����;sr]=m����ͨ.W�7d���;'^�]n˳���#b�шܼ��v�7N������pZ�pO"N��=���ې7�ly.�U�l<��A���:8������H�n��I�ۣ����ϝ��	�Wm�[��m��<����8�9(��]���@���q�z�<�o:Ź:1��]�v7<A����^��i���M�ʷ���4��`6�{u��ʼ;�4v���,�@h�1��'�s�n��rݰ;�X�Vwg������lk�m�2�Z���q��0�nt��%eèՊ�;��]@��Wu�;n��9��湳	`������JN���ks��k������]�G[	���1��w356˻�n���5�R���ssqֹ��=F㣉�X�0��%�v�V6Y{E��u�îu`�\��Ň��7�;l�i�����vãn��-��y����qV�mܯn׌��Q�2�ո�-y祲qu��[n��]�L��ɻk��z�km���n�����{�R��i��;��n��lL!p'���y�r`�*��5�]� ����",4:X=b p��d�|��'�:�!�16�IU�1�!���bbo�X]��un��������
t�<La�
��>y���ogY��Ч�<O6�)�M!��y��kM	��A�P0ɍ}	5������TƼ����C��߷��;��t��>VJ�O�Wv�QH[I�:��O���5�Rb'�{�=IR|�LWS�O��t����q�9i��C-��3i� M��v���1dE�t��~1�$�Y+5͞&�*����:�%���g$8���N��? VϹH,��}����2MB���������\��]|���y�$b�Sm�>a���'�����3���P#o_�P�H�0���"��I�֥dX��y�M�7��޿z컅��*��1�c
Ȫ(�j_|w̈ӯy���)�'�2����uUO+-κn?=��VVJ���c ��@��ʳP�����l5�Rb�5��;\�nq>�]f2Vw�����'��h��*v�S1]aF�\�B���O���t�o�~���aS�R
Fڬ<��~��O[�����/�t�4�z�0�ϜT�j����ɝ��{C���nZ<���aL��N���"�2��O���0Y<cl�������z��x���ya��;�i9��!�מb�a���50a�v�TRt�r�'�܋��y�O;�*C{��V�=��^����߳��<�)�u׆��һ7v���TY�O���6]����@�6Т>����ێv�xb����>�ܜzx���:f0�UE�v�sy��Y8��>OXb��1f��zq�5�Y�j)v�0�:O�W��߇G:'�I�5;�x�'�=�s����_S1�3�jx���:Q�N��N�x����߻�3>�-�ά钽����3�FӶN'��&��w��x�~VO/�s��IY|�΋���˝n���R������em+�z���u�C-���3y��ǧvϑJ����o���2сS�U�ϻ��<`�h.3�8eQf2{s$���!Xv�hbc�7���a�?~�����=��Ud��*FB{��\��4|�&��G���J*ݻ�&�v7R�gQ�5`�a�"[�N��f�g��r�{�G��â���Q	έ�DA�����'2�d�m_���x��>�]�oRj��gi/-V��bu�7�[ghb�o9MCm�!��
�Y���8���,�������'|�
��'��c��@��3�����<C7�՜a�q'�v��d�bc�1��Iۗ0:��/��o �ȵ��Cz�I߯�{�/��?�t7��fgl�ٻ���n�Oa�?!S�B�e
�Lg�1,>d����jN!��y��ҲVOD;u.Y3�Vq3|Ι�s���h�'��%�jN0��Ӊ*q>L`�~�����vv��3	�����3����{C��+��,5Wks$��Yg=��:CS�{���p��9P�Co�ۖ�Vj���jJ0�����:�^�\��'�`z�Ι�1 ��U���aߴ:��~Eg��������Y>�c1�:�!��}��{��Yr��IP���!�a�P������޳�����+�,Ym�c1���1�~ζv�s�c<���9��f�'J���q!��S��گVMI؂�����~�
�ώu�w���yg�!�H+�������I�ԟ���5���n=��=N����>˴P̡�P?sp�yd�y�}��~�|�5Y5&�C����:��
xr�'�����隚�)5�~��zNnr�0����˙�K���5X~O�gI�M`(��'�d���ȳ�Ϻގ��33���S�Adl�c�����|���\)�/���o/�q��mK��gK�t�er��߀阩>�?��O�Jk�8�����|^�2�uOY�!�>C��>��'��L*Zg�\f��t��&+B����L��:d��wN�kf2���|}���/�e����n���PM$xv�%�7��ԝ*cBs��d+>q%v�#ٯ��!������.)
�J�a�I�³��V�\�,���*ΐ+�Q`,��~�����y�Ooy��y���k5�[55��aӯ�̍�?�d�W2�����wl�C>��|��S���}�{IÍ����ۖ�mx�t׍d������L'�ğr�,����w�߹m��^���%�Wv��l]+��T�O����\o<�U�I�,��QT��p羾~}�����PR�T��i�霱��.�bd��Sp]���Sj�!*��ڪS��]>'������� ��MUUUUT�*��nF.�l�h�n� -�Vӭ�ۗ���N&?�ՓR|0�
�����g��\���$<j(T\LC��;�*{��ϛ��bT�У�@U��,��Y�s��8�m���z������x���~��}��:g�h圿���u�;�}�FM�~����e� +@x���#u~f�zf!�T+S�1
�{�jw�睭�]����+�LI� yj�Y1;e�'o�"��na8���P�{<�w�S{=dZ6�Vx�>�3�<�S�j
|�Qd:�T
�z����+:���A����j�L1'�J$��*,3=�]��}��a����7^��11#�o����r{����
��d�y�{;e^r�o0��q'�8�Ն*)�rʘ��m���t��I�
�'^�Ǯ��
��U
?C��A�?�mυ�4���)�0�;�^o}hVJ�YXw���~�'�YUĘÊ3�c=aU�t�ǜ��R��&2��?}��C3uÓ�O���t�0�5�ɨy�v�3z��~o�9�G�;�k��<@U����,
�������������;m͎u�X姁R�׬Yn��1�۹���|'L�����I�pX|�埞yd+:WRbn�5TU2���'|�3`bk>@���Y�����=S����׻=n�:�8�C@U��Y��)���e��s���( e�D@��8�`�ʕ ��?'k*击E'B�8_<��5���s0��S�<�jE��0�Y=o������g��u���w�����*LIؘ�f1��ڪ���I�����R��y�x��Hx����v�Xt����HVm�{���a��E!���,1=|dĩ�����h{���u�����La���*�<Maٔ�Ӭ��~�f1����w�m$ɁĂI�!rH�%��s��.�4��!�Ĩ|��$��<Ir�E8�����&<��5�C53�%TR���٨���11>癬>��/l�}f�+*=�hjs�:x�����c��y<_w
2�
�2v�T5��|�3�������������¦
���Ȫ,��+��|ɉ�<��;׼h�"��T��Ԙ���T�����ސkӐݳ�*�C��Ϩ��`��D�C���Kp�5ۍq�.�[�a��,��n[�u��<�s�qR�YJ�9�HIJ�q�y���v��wQmƶ<;69vx�V�c0�K��7q�Č������<;����cq�9�ue]p��q�f�a�>�x㊝^(���y��wWlz�a�jK�/���v<�^J| ���@Ϭ�%O�+'��׽��_ƞ����J���s�v���*O׼��l1��W��C7δ�u��Cz)���:�����1v���5<n�|����\���wz1���QI��\j����1aS�j^�c���!�0�%M�a�d��'��Xv5L������æt�m��~l�x�@Ă�����N����Nnr�GʲV<�u�����<�(T=ˬ5��dS�73��%{`g��<B�d�v������D}tB����=AGv���g�̶T��,醸��dJϺ���sN2�T�~��a�bN+)��Dj$���l�Ah�BILl�0c6��� .�=�w�&*,=��:��p׉18ϙ5�i���8�2Xk/:��{f<�0��\pa�
�ä�e*,���I�;:�;dS�t��听�d���Ϲz��u�������v�?,8=�q�ݏ�!Z�����q�R��1���C�u��ԇI����9CSF��,���Y~�:�w)�
�,�μh����$������~g��{��0�DE|���;E&e��g����`u�>�9���c=gOIS|��
�f*wKI���&"�TY�w�0�u�͇=����{sqz"3S�,�v�yOP���u�*,�R|�uNޙ�����ӫ�9��?M��c�]i�sI�w.g��ĝ�!��TY?!�Y��0��8���ͳ��=�t�SX�t��k8��'G,1�}�J�ss�L��
�Lg�$�0Y�+ ����}2���@59Ӌ�lDt�|0~�	'J!�#��Ng���U��x&�a+�Ԏ𺍯p�˾�m�q�
�g��nD���^~��z��D\Awt
%��8N����ǧ̻Hz��_���h�W.׾B�nvFկ]�ùޭ�G�����x;�ş6�7z��I#h"k���[�8b���S���J�Cf��~5iY�I ��-����s�O�o]���A����emJlvn�ھ
�;�i3��wʵ����h;��o�4�Ug��JQQ��Y9�+�u��2kGp���A�ר����V�����ՆTQ��T���Q�H�͝�FI�LBi�s�c��뗶���*۰�vl�|��	\��{&f#�M�[�U��J�v-�)�S�)Y��!)���j��lO���j����	.h��1�7�3"I	�M�xL<�Oi"ԋ-�I�}9�뻽�2D0��N�Sqqe����Ǟ}tMciƐ�H���1��IS=+	����P����΂��C���m����wz����䵗R(%x&[M�үU�G}}��?�{��뎃4�}���ض=��nH	{{g���S]�	�Q	G�?-%������N�/rK�c�m؍����1��5��|�rж��&TNHXj��Z��OS��-ytG kswJ<�J&���h��}~���m��j�����FMj!��el��5�O>YHz��N>d���z�i���&�
��=�XOL%���J#cf�N�\�����C=�wO���MΖ�˛F�K���*�"S�s�A2V�Ln|����2���L���O�m�6-�ݍ%�)�[����.޷#�7
t�U.Ԝ��C���[������U�}�����;�X-��ۖ��zڍ��~�5]�����'����6�,�p'x��?s�VJ��
�g+P��2��b0L�t���w+��2�n�5��M6<={��Mԫ��7��ݳ��y��v!_�aUG���I�y��U[K�fz�8�!�Flz\�����NvԶ��K�1J\|��T��S����F��~5[�]���Zd��&�SD{�L��g������Wz�P�6�)�*W�����+��[l�=�����շ��QdO�D���O(K)*�ECs;Mnn��ԗ0U �A�+�;I��F^�Wf�{�Q��ܘ��eSm��}���m"�X��vL�}<�W�"��72tS>�e����O��u\LG�%]/St48f箶�����"���6��G�=\9�-�ۓ�	mm�g|�ń�ҽ��F�K��
&�t^�I0��^���㰎G�Z�'��o6e~ke.������O��*��R�UR�p�&M.�ŗq��Q��N=�"���~S�/�uT	""���sK�IA�~����_�v羵nR	��ֻ3�.ٌ��r����dA:�w��]ՠ���y��Mg}�Sw�)��!$׏\��-��^a�\�.l9J�������]���ElI(�[� �{�
K9���+�F��<i	�M�d��w��R���ow\�Uy����[S�䷦'�N>�4�(̂	w�N���%v�������"�{^�(a�%êR�m�4�ɷ�>h�>����W���J���:�DN��.k�TRY�b��5�o����w©!�UiN�Hq���ITع��x�d!,�Y�Q_�ύ�U]HL�켑���V�tmZiU�Y�UUUUU��*UUUP�͡� =U�ɴ8�$�m������jB�TT~$8��ͺ�$i(�,v�u܉����$]7\�z/���X�'�s��;��kCn�E�u�;x.Vj�!�j����?K1�2:Ύ�����<A.�z�}RH��sqUv�mTDc�OQ�iU��]tH�a�8�
?M��Cސ�pI�c��.�%�g�	�몏�w[��?p�:�߽��U�Y[xp-r5�2��;��lw�/�y!֑�蹓k\�5Q�����^��c�km���������{�j�fj�H�t�O�7����J=��ACq��J�T�	-�޹z��]�$i���`Xw98���v���;Y�A��5�����A���Sj��@@�8���S�ku�əI���mӝP�ct����l�RuZ�C��^HY�E�9s<o�r��!��b�����$_��/�^]�}�m�7X��m 0���s�X<���|q$"�w���Z��+-�m�yK�P[�J�M�,���H{$���ꩃ3�wAm�`�%W���ʡy-�}�����R16�Hؕ9 )E �m��� ���+�_]P/}N��]1RH	���6��5c���i�6MI�N����"�Z<��Q�s^�T�Mc��.P�n�L�̹b�K���yO��U ��ȝðLt��m}[��~~ݩG�;F�e��s7�w��q�Z��oo+y��7%^�ܧ}��s�}��{���E,Y��>��"q��/YJ�(�]pP֝M�#�&�:�9ܦ0�K����`��ظ{�	Ǐ[�ӛ�`/]���4���̛k�.z/��^�Hz�7`�:�:��۩�l��U��3���v�u&ܸ8v��,�ڀ�"vR���]7�K��2`�g�5���qب"m�7��搪�{��11y���80Xzi|�N{1p,u�i+�e�[�ˡ4��Zُ��C�	�&�HZ���-�g>��Y�j�BUg�ߥ|�^��4/�xx�os��n��:%��j
A�i��?(M	���&��'�M-K3.�I+Im�d�Ǭ�t
���k۫Z�D��"$���z�@�^�n�f鶀No�\��As���n=A�ck��$IK印��AhJz��з�Pmֆ�{w{�7��W����݆�L&⎥~�Z�<��e� �!*i݋Ђ�؆@����U9ٔ�ױ��r%��^7��|߰IG鎂$�*x�ĸ���U%@����z�������{�٬� I�}�R�ff]��7���p�b(�Q�Z�J�U[U]qc�?����7�.�"_y���J�gZ�$�����km5b����4A|�6�l�͘tsk2(�Z��*3fEx%�>�K(e���'�m$�Ɛ�ͻ��sq��t�6P(V�j��o�Ji'�/f�f��}�_j�f|Fx$D8O��aָ���c����6nL�vD�ʱ��J-�H���g�ڂZ�"Xgnl�W�tL�{UF��yV9��v�3��j��Yǵ��QS)��{alU��]0�����hCW*"����]~�c���)�N��~�v�X�8yQx�N�S�p�t�^R]&�i��g��!F֮�l�����Z����4�M�DE���1ql4P#9iMt���࿸43�(RC�f�
�b;1=�w�t�2/�6��A�� ��{��j��*���U|xGh7�E���/�Α��0>��&�gs���I95�X��+��e����'�u*3��=�n'K�?���/�n�e���]�.M���0..:k]�-T���zGΤ�C32�h��Og�n5���ݗ������9�IoF����f|�ц��b��&���\C���O�9��6N*�AB�\̰�p�"&#�@�5T�p��Ș#bX��,�������,w�=�p�qlD�U#�H�*�ѵDW��?���i��].� L,/_V�h�D��+Ϣx�9s��ʹ	����v*8�����-�&EG�f�W����'.l�ϋq��I��$3�ó�N���(�hࠖ	���x"Ț�s"I꣙�vg�ѐ`�����I���R��i@�I�+Q;�F�p7I䚶k�K��wx��8�5��#���d-�A�n�l��3!rI�ʵ��ldw� ��-ٍd/�a���v�-]��h��l��xx6���)�u�[�2IJa��ٔ�۞�4}UZ�0T�$��.�����.�|� ��$]���l����C���&k�l�{��/v{�=�u���"R��Vr�9F�;&p�Y�څ��"�*ԙ<�4�UUt!eo�/��������+ɺ3������!;v�ݑ������7^xB1��s�`�5�΅��D7i|����Y�u�����´FT+�۹h�t�$Oե�7�#kA~���1;�?)��0:���kz�vN������2PI�ĉ!�>$S�_v`�J��'�Snw��^��ɦH�K��^�(����v��i;����¡uZ$eL������n�R\�F�K~�Z��<Hqo�F����[������:����roi��6�%n���ˬ<zظ���T����(4UK>J�Ǉ�&�nI���
Ŭ
�i��@�G�ץF�5ҥ��S�����YΞT�Q�V�ʆ�],�؅� V�̧���&D�e�mTEj�t2�������5���ɾ���*(ii$��1�\3�{Wg�[u΍��мdG�_'�]���~��UD����}��:��?/.�2����T�,aa�)�J�6���M4���M�	�:����Q�{3YL�E����i��v���o�a���
�Qq�2��ŧ��J�J�!|hHYA~?'i6�.���@R~��3��Y�������u����9Mm^$�o?-�I��N�iV��s/4�*=4U�E���܋�ҹ��SۮӋ��u}�,$�lC,��v8j���&q\�ں.��Z��N\H�ê�n{��ch*ѓI�;w�8�-Ѯ���mb��)R޷��ݾ�\�㻧γ���4�Or뾩�iuɵV#������J�XN/*W�_�fk�\���6�a�������k��G��w11HX�T�rN�1!�*��z�M��Nl,UO��ױ�^>��L�G��'�"͛���ܼ�C�Ot*�S�I	
JK�D*�k>�kxa�}d-lj��yL�.��Ś��yU-6:�U=������%���O,~$�e����>P��g��`�=;�MQ^����,�̣���v�Dz��֢�y<�^����hxK.��^�j�}9�w�V��L�w9�d�=kv����=5^0U{5��eש��.��|���n۷K��܂����q�M�r�D�Px<�x�y�z��=�[���
[~�f�齴$�fW�����ѕ�۝v2{�`��UUT�b�`��UUUUUJ�UV���U����h��ZE�ꪪ�U��U�j�ݸ���A��bY�@]t�EA��Yeq�:j��������!sUuU�U�UM����*��5U�UUuUTڪ����S(
�Gk�kP����/���j�����MU*��@�(U�Z��5�gp�	�PR�jj]����UT��e����VRe檪���%�v�SKT�^�)S��n]������
��I�軠*���������������������������Z�MUUT�*�UUJK�M���V���V�����������������Z�����_�*�RUUUHR��P��T*���������ƥ��j�������KJ�5v����UW�ףH|� +Z��V1�A��ԫUUUUV�J�T�R�UUUP�.�;ODM�5qD�[U]OlY����?���P�K�h�y�	k�������K��mp7���U��J/�+���.B4�T��+��V��[.��޶-��K��E!��P#i4ݼ�D�#�,gS�"Pm�~�������CgͲ�e����:�?�Z�	g�ADD�����ۃ0�		�U靧*�ɷ���"�BI*s9ԢqE��D��:[��d��[�M5V��}�qE#1�=	m®��ꛍ�X��&�(����]�&ig�Dͪ܊BH���Srjd��K���󔐪��^t4U--���5H�����D\�� |l��9=r�_UWf�̗��̬c�AJ���3U�$H-4�̭.gΖ��r���W����q�pD����i�\2X�Ǩ:����7��ۖ?�.����IRG�ڻ�*��I��0��-��._B��J޲�@�A"I(f^���μ��[O{y~��Tds������@��m.�H��h�M@	K��˺4!������\��-���+���q_����-��c|��34!.�b�ku4�T���d���Y��J���њ3B�{5@H�u�VWtc~s�kٓWJ,���昙��M/�U�TC������?Um~F��+~��N*c[o��JU�ru���Г�ܟL�7�!$���7:����u��!H�����]֛[��m뉘��[��၄���S��ӗQl�͂�i�ף�?��؟L���5z���U.o(�D܆[e����P��BB��ƪ�oM(~�[��ڗ����;r��@*����\��ٗ;�N������b�m�c���W����8͛\Q{q�}�w��h�:�K�W��k����ڞq�;�9�n�S����C����v�����s��=s�0-z����{\]$�.WRY�mqd�u}��?��{��mS��D0�W9T�w�s6I$�^��쪛�����2��g�Z�֘N�"3���<X�O� ~�eJ}cgUp`n�}!��>%[t��I���f��P���iϚ��=�B�Hp�Z�a��5�\��r�hm
m�6���5���l�I*���\�c���y��iˬo�T��-��*���*l������$��7�T?{,Y���^6O3jn�%�oOr{m�\s5<�[[h�Իڪ�m�K�UH�2vf�����x��u@�Hڕ�i#�$�m�,Ӫ�ތm����|z���1eyf��G���;M���Zi2��P*�
�u+l��L�"D��� ��?�OM�b�FRY�^���A���^M@}$�m��JN�s�5DiO�l:���D����=P#�6 Zn��-��be|�P=7���ׯi2#���ț�PQ��{KmmJ�;EY����=��d�H��:}o�K�Cm�․���9��E�|[t�}%�ޙ�u��G�>�����$���ʂ��'��e�>6��H*skl��[`���RPd7�00�׏����n�Q0��v��?Z[��g:�p�&��a`A*I3=)3QS�-vܴ�%�=5ɩ��	0�܃E}	g�D-�{����D�[n�}=EHFlϼ�a�'��p��M�$_JYwJA�(��VCBwT��"��4T9��ާ=���W�~"^+~�m�]���[�uTJ��[�UV��[�G�,k�+�Y�W�% E��uD�"Y�H�����u0���[rkp��!0�g:����!��O�m�QU���^/`+������Ւo�\�-���.)�<���L�@�$j��z�{.�/�ܿ1�\/��"�9�V�B��˻��a��RQ��~ �� >�����8�o�]@���ێ0���$����Wy�!�㇍"Kf�OdF�����]���T�qq"	����Wo>f�x�&����g�!UA���_�̿�FM��:�S�U�$���B�o���$eBS[�PW�[�5��]��E�r!8�fE0�B)$��v��@���m��?��^m�H�	�B�xC�iZ	��=r*p~V�7v�γT~/� irN�~��Ttm���[`u$�Ȇ0���9B��~aq�B�ȕ�	� ���Ve�*+�"�N�V@oy|�a RX麠�[��5������5�2(u	:�Aû	9+iO�󪺧�C�J��5l0�����h�Yc�4 �1>l�pa]Z϶oY����-�a�� ����)��h�-���t*����)$����[�j͐B[�wn+�0���y�aC_RA˦ꮜ��Ƒk�d��"���Pm)�w�fNl�m����n���˻�#|��5[��l@Fa�&��GqkH����BM&�+$��tܚBD�.DK$~?������[�@�	��k:�nfW��:��@_=H?�Y��3���Q^�Kâ�	ۈ��}���n�+-���x���C*�m�T^8���7��ə7��h@�P�y�!���!Z����)�G�{��S�$��^���N^J���6HD\cc��j�=�s{˴b�w3t.�	H��l�r����f�DF���C��{|�+�v��)0�*���}�s;��i@Xΰ��HN����)l�����}������W:�(DV����+��1��?�	iCDY���t��Ww������F�'�*mt/$ko�s�D�#9�nS�� iO�{wcj����3�j�*�7#�36E��a��䆭���*��gS�d��z��.����K�����4@V�嚄��L�;j��$�#%u�e��{ļ�I
[��-
��69��UK0`'����DkB�����B�^�)��H�		��'B�����Ԋ�D".�뺙� L�C��P}���ud�io�hb���{{,����b�Д�aE�ң��
��u�ÿ
�2��7��f�9����Z�Uiݘ��0*K��xP�=�\u#*#�D'	8"��[F�]G-�[�nl��|7���6�`�Yi}�Aw�K�	a���4_���ÊO�>;t�R2	���[����6�\���6	��,����"�]�����T�	e�J+��#��ĄF>����d�)i�z��{�Sq4�J0&��������ͥ	OuW�\�N*|%,�B>�Z�W����y��1�n����n�*���T%��Ҫ�y�~Ͳ9ʺ�=X�grȦ�^��T)\���ͫ�oYZ�Us@e�!A$a�H�Zx��Z�����UTQpY%^����`�L@��U��G��������@VU����j��h��ٛ�5Ɗ�ڍ��*BJ)����=�j��!�阛+��v�1��˚JG����e�!�9���my���3��r[c��ǻ�{w���B"\�UM��%%��qF����6�S񕀷��\eW�m��d?z@�	M��R����.��v����*�5���։����؞������U�����!���8�b���A�0���G9OweiUCk|��/�Ͷ2�U��AY!z=����&}2��:��Uj�)��I�9�ND�N����e�Y������p��H�Va�܌�����b���� ��[���b��wG,�ҋcR?p���59		���'tL2�"��Că+�y6/�*�vY��:�p\�g�]�ٹ�`i�[B1�؏�;me��V�����/E��;��F��n���[!gQ��~���P�
�i�B��(7%gv-p@�$�5�<g�/��0�v,x��S��q٣_���t�c�-�I':j˂Q=�YO~�������!OԳȢc�Um�Q��%�/
���f��4��=tgF�w���rò�
:�H�����*8RA�ؗ
.�%��t���G�ΎM(r�SD��x6A%�1j1�[f���CSӹ9U��	f�'��Wk�� pQ�a�1W=ȴf��8Ȍ���9��G6o��V+D���z�\�\���w5R��q/�䲮�!�p�l�����..�����*�Ovqe"3k8��HD6��)
Hw\�8ѐWmh���7���Kɬ�\?�l�
|B�=��x{7=��ڧ��:�щ����:��ٷi�'b�ٓ<�ۖ�A�e[�lr������+k��s��I����xS�׋a��pdHP���|\�8��]���
�nϟ�J����ޯ�'�-�\�"M�X�
���%~�w��a+��|ȁC�t�cQYr�7�8���u�L0���s��m�3�w'1=�q<���a�e����� ��p���B"���g>���O��ө��f�hJ����C�l0�M�r�=�Q@�-U�"�,�[���׮��b�XE$�n��u6$����*}�/���gm�:۱���+��������\n�w������8uh�����4!"1|�k�ڑ�>�?L�%���X��)�/�	@�T�$K���5N���Lz}��pZc$��b�2rJ��ݖ1��w#0y��%sm��������Ox=���Q-}�����Tb᭒b�U�����۽Dd���a6׼�&�:���ހ�[;s
U�����L�dJ����2�Ҋ��M)���F�$Hڐu�T���\� ���y�RԚ)�/��ťw~'.�$���"�d0�7�&�I��V��m��6���I�r�{p�+�#C	H���$� �{ŉN0N���K��Ms�����oj����o�|f�q��[�uU,�٭���6�Б���#*eP��IkyL�I��۸}(�v �Hr�����u�<O(ga�H���^��kL�Iyw�DR���������>�����^�OntU1UD��d��C/k��s���?u�V[��M�Y�����k��E˾�`�s\Q��h�x��{��kau�5�"pSe��_T�hw�r�Dog#�1�������Hsh�N����S@�< ���������;�mQ �$ؑ � �Uk��s��n�7���{WlϦTӁ@3�	?� ��n�}���3���;ڡ�J��e�I�;j���{��{�n�fvc�D��tl��[����Ah����]�P����s¤���G��ۧ~�WmV�ګ L�T���5�랦�P��~>$553�>Jɇ��/ÆUN_i�F�2Ꝉ3�F�SpɪI�:�P4�Qh�	��{�j�Ӓ6�)9bQ194�
��J=�R#���RE	���vf�\��M!U>":��Ѐ܆�̛4���!�����T�I@	�X�.*��ZNe�0�#h\UT}i�.S��8�W|��d�I�XB����:˄������lDk������#R��d���CCk�=:?V%�w*�N����mq���:�묕i����T���2�V�U�|x�%t	�M�H~���=\js F�U�U�+�$�n�b5������A	.��p�y��23N����������n�uT�3��?��e{7v�&�qx�4��o��[�JY
V�s<
S�����[�h^]�+h�d)��tp%�_�;���,S�A�Lt�t/��|ی)�E$'R*Dt�L�S�^�����|�ִN[I����'���c��Q�;�)��H��=�b�H^0�'PH����qf�x�,�9z����ud���[|�8�vpTZts�r���z��w�^�[�}N��Y[xyp,e5A�E�l����5��r�1��<_%���m�ʠ�����bÃ�N�).T_�G�3�n�}�����yA��Rԑ}�����̽4�[r�������*���c������-A�6�wsHu�?�C��

@F��'GD���Bi�$�:����Ϡ$e-����}tK�k� .H�߄	������jݧu:�V=a#�Y{�BЫ�y�S���α6Q���a#k�I�(�� ��d��}R��/Q�b3�#fzm�I��d�K��o3�y�%Č8
�%�T��	Hcb�tZ�6@�y��u]����0��ƒID�4�LFSa�R�P{:��B8C�Q
�ʮAy��_\WN1��VC�U];�y˾f��NT��BF��K�	e^Z��'4$��i���뽞���� ��	��v|/i��A�d�� �&8}^޶E�䊰T��wX��1^{����s.�Ϣ��9PC�۾�F����R2�6���l��A3a\lɞ��ͅ�Q��7xP$b�.Ș�7�!j�1x�쮇�'7%I=�{M	hc��p���k���x�UNqt�C�\A�0q&=�x!Y��ߗ�I��ӛ�rzuwG�C:���
��39T<�T(,[�oc�ӛ���4�5���7�H��%%*�UUt�-�s9�fh���ꪫ����MS��]	�m�Uk\�gR�UUUUl!Z*�Z�����Erh%�y3ӝ<�M0�rH�,�!���<����<j��e��s�T�Ӝk��0ص�l-b�s!���
�1ĵ��V[���ZbH�Z:ʁ�t5�e \Qzo<�����X�yV�S��.��/|A��#�=+�1/��#_XM�_n�|u�*�z����:��:��35C���WZ��m7����8�'���{/��_�],}�X4��dn���8��$�N0��Y��|��Y�?�EC�[�뽝|X��%�)/(���T�e#����߶���š���C�&0��"��'�P(n�-:��c�r@��=�q�ot\>bU�-���	�푅�r��p2����8o,��Zg#��QZl�Gj�4��`��2'�e��C�������RW,��� ��ρ�z�l�KK�HZ��cl{#�9�6������L��tp�� ��;�/eg�~5nC"�#$.�L����?7���֍un1��"�#@����!�Fg=Jy?�Iu;�ޕ�E���KJ	^ԧ�8�6�3���m3���AV��R5Aj)$��=�t�A�==��~�Sv�.�u;���U��WC�d���W]h��eO����-R���q�w��לּs2�S�YOkNc����7��@k��\�Z��=�QJn�U=k]��]�3�/���6�R���;s�g]C�sS��6�nց�7��t�˞�?���{+�d�庛�;�����Hm���G<<�.�	�D�e&��g� �r=l0�n�22t�[p��/�1G=<,_jl�:�^+�ףO,���Y&RI�&+P�B6HճFi�"[R ���
l�+�����{�#����Չ��k���7�D�KȜaT�x4>����H�2OR���kn�%�e��Z�[�f¬Ƥh�S@܎κR���:�)��U�Z�ǴG��"�1�	�E/�'�qV���	A�����8���/��g��@�#���<��<�댮%d��iD��/&c�eH�`��+���*���boL���ɚЂ�A:���Dٜl���fu,�n�k�'T; F���*EL6w�l}�͛�'��w�gkד~$��F���$��$�mȔ�J#���/^�܇���gL��@l�PS|N^�U-K��&u�X[�4	�
��-ɉ��;�=X��@ O{Z~�3�g�%#��]�A�v	i]��m��_f8�l���I|�.
M�����T�}���~�y{�R�X&��&$��	C��/6�R�r�%��6�&��z�
 ����P,?L�?T�bQ&QuS��h!��݂|	��R�r��NF>�x�ĕ$�]�IW�($L|%�>;nub�;Cz�P�eu�V����2�P&��ums�yMl��_P,�:P��G݀��Wo\�ݭ���1�-�Y�	�͉�=�ٶj�Ǯ.�ٝwo�,�UaX�5[���S�2�f��/"��/_�����D����Y&9�_Z��
���{�p���S�*^�qꨝ�U���U^���6���t<0/y�Q��NAwf���+1n�Q�D�������r$�1Y:}�؄�yݯ���G/ɵ��|���l��Y�8�(�T��8s�`���^����.�q�Կ7KOC��⇉NP��Tۡ��S����Br���n����C�n��53��̇*�
�Z`��63������YO=*Ueh=�*%=���|>����s{�gI��j�&�;Y�wdaW}a��5��r�tw���ޫ
zE��κ�_���Cr)Y�Jk*�û�-YL.[՘�˳�u�ʱsz���p� 뺤#P}7l����߫+��ҭ:�w6ĭ�)�*UP�M�u���8]�_�tt����b������F�T-3c3�S&�r��9����Ca�52��S%FB��5UT�\�l�N�6y!��\�f�`��4n4�p�d��\L��w���ܾQ�ձ�[�m�헀�\�b��W[[�3Xck�ۥ��8.��۶�ݵ���؅긜Y�ٜ�\�m��'/@b��;��&�q���X��،r�J�Y�n��qj�S�c
�<Rq��/�i�b�nױ��q�-�p���ݷjsm��:�%�!�ͫ�B�z��é��)�9�<g��m�:�2ն�:΀b}ۢ�O0u�v���ل�r��A�䞱/;�c��w%�=���S�n� �n��z�}Ru6�������"�E�P6!.��� l��уv�M��6ۇ��6�Q���vaw7Y<Hu��}��2<n
��/`;��s�wZolq�/4:����żf1�;buu�Vt��Ҍ[�p����)F��χ��Z�c]79���.�q�mۭbڽ�s��Zs�N��vYn�í���v�h��Ռv�۫�c5u��[���@O]��A��8�G�6̸����<��F7en�ŭ�xxLzC�f .�P��zl�m۝��]i��l6�%/B��N-x���vt��b��&�j��<F3ɺ.����6�5ڙQN���[k�;n8����od܇iE�A)��G���sbYC��t�Rzfd�5��H�I��	D��V�l�c	0�5�{��.CTZm&����*o>%���c���ΌD����������s�*Q��H1�"���M���pI�I�IbQ����Ln%&�̎�3>i��ߛ�I�H�d����Z+ћ������?"�rd�B�F�.f]�$�J1�mkt�Q(�=��;ݶ�XY-����<F���=X�2�$�oR�BX	$�Ჟ�ao)���|�*@`��$�����$�x^s��zhhJԣi��(�nF͂8Vu�T�*���?77��n�%�zv!D�P0��ޭ�㚱j/d�	DzF�@όA���
ä����6��?]�H�4�ց�\[�o ��_��[�˺�ҴĳA�o~��;	�N����b�<r��N/��%.�K����	U�J	jYG�nM��ܣ�dK/$C[��(#���͵q���Nt��B�~%k�'�jI[>�|�Fi]�UI��U��� �B��,���r��m��#7���-�"�%�i$A6<�!g)r�����b\s������R��j��,����B��$NO�tѰ�(�E�dNy�͓��r��n�v�>�r��B��+�"b
�rL�c�Q��dئ8�a�����'%Q䶵��"3}�
��*Ng��.X�5�&�sI�([��oD�4_cᓎ��X����ը���J�-�{�v�G ���TQ��O�6��Pa ��Y�D��?�g���^'�Ɣy}�[�U'�/�=EW�i��,h")%4��)\�zd�M-Joꭢ.�{=L�j=����u��絛��=�d����BaڮM��T����o����������n�_o�:��u$A1h��]UV�Zyv�l��t��5}�Z�R���=m�[!� ��i����J`�L������A&���mP븄=�MBKe.wIjyH�c���?���i���}�g}��kD�� m���� �J��1��e8��w�!�M}-_��|un��aosiْ{ҍr0��R��%�¶Q����j�1$>����H�+�q_�U^�T-�v�R"�^�KBfe�m�*j_m���չ���n���Oڪ�xq>d�&v	Q�YUx%�����F��^�d��֜,B2�7�i��"P��im�6�;��z��������[�i,-�~���YwAW�;���F|��Og[��Ffq��J�1oyS�}R�eP�A�c"�,�	27��qo�v��r�ی�~Zѻ������"U�4��İ�?p�+�ػ�������F�d��ٟ��r8*�̗A�W�ǒ:�!��~��`q���zRl��Jsfnmn�^~�*i��B������0���t�}�#;.����\�k�T3-eZ�{	���r$ؐ�M� T�Т�UWX��V�����W���(�&�:E�3S��&�-*�UUUQH*�UU*�UUUUT�T+��0V;U�*�UY������>W�>��k�Cpd���F �%���f����0�aKm���g���U���}��o���MD�����[U�΄'O�y&BN\ ���RA����#�T�#p%\�m� ��-��Y�҇�=���U^�K7M�R�g�-�(S�&@ ���Lĳ�-��&!gw�Uț*���TCq�r�����L���6��^ݾ5�m�A%��RUn?��{v���ƥa����HܷgO���1��3ue}�M�R�p�$�"�̞�wt�*�;PZ�O���>�m�a�U3iB���f�$aW�����ϟ>����0ӻt�ȸ�g5*&D�li�(�uJ�J��|���ҷW3,��LɔU��`L���˲�)o������z�$�UU~�ᖤ�����[���D���b[��*�v�/���30K������[!��k��?C�UVd���+�^�>����m�m����ׁ�l�	R
h�
$�&�U{q��Fc7X�a[�fo0���<؛��SWl�T�-Wx$���~�O��I2]�fe��J�-�o#v���Ъ5	A4�hHa%��*V��n�X�ȈJ>���7���z�Hw�7Y���,$�w�ً�C>�wO�|�%S$�L�p|.V�1��2y�)Տ�W�+��[�P�Yٳ'S��ʽU��]�9�x���A�"�e��I3���N���0t:	�S�q�=<�Z��YC��u&�ͥ�kvj!��ɇg���_�$^""cx2�(�n�C�����ػm9:��Vp�%�v��l�����5��
�ƻdC��� ~!��C�_�m�8�Hh�����[�SO�&?*��&�t�5ƙe&�'BMn�������!ՉF�%<��'�l=�R�����-�YW<hQ���D����"v�mK�(�����2D�X~/�$�z�[=	Ntvw����`�o[��ON��p�)4��p��w��ȓ��1VTe���̲ �Lk��~$h�[�~1�^���[탟U����=@v�[oۖbP�Q�d��8
�	#��}}.�lպ��q�	淩�����_<@�&8�_UK�Λw�N&��gWȑ	��mUJ��L�D?��&"0�?m���
��-|��(�k��Xks�O4�y|����$��
�~�޽�<�f�s�`A2��ûE7��	`!�*I�OV�ܻ�2
�xWK,��i�F�h�`f������oߥL��n�F�L^M���饕R�u�^���>��Ko��o�¸|�+����1��ҁy'uUUsn��E��/�zf�ɿ7a%u����'>I�бŶ~(-�.%�L��gK����$��6Z�uGsC��_�$'o=wuM�*F�:b����T���s�\��	�CR���Iݩ��hû"֒�,��榛�ܷr���0� VAw]�Խ�l�PԖ7���S��
�`ؑ˖��3�m��OoCJO�N1�g�7�]�o��A���;,���'PI�"�[?Vf]��G2�F��J��˴Is�wQ�7Nͮ��d�����ه�O�~`������Qp=7��7F" � E�$h���y!뼠(6Wv�wO��,�OoZ��IZL��5[�m���bSѯ����i��{|x�&ZL*�RD���o9����S�BJ(���W2JK�.Eż�Z���F��b�8���g�s^�寯��	8*�zլ5�:��UJiL����B����o/�2�<�H�|���2_JO��33����D����}_��v�V������\CmB��$"eS{iHib�^�j5:K��^,bt��yB� ��]nl�\Ta�����U�ܤ70��� ˦�](K߶�'Ơ��΀T����w[�Gh�F�O+b����Pw��B�b�+���~'��'�EuU�-���$l%\��J�`O���E��Y�T�A���U75��Q`��1r	ι�Nw^�/�`�)~/p��m�a'�Y;zڨ�U9P���!/��H�K�ż������z0��L}nn�NG���_x�U1]>�JM�v p�Lv���di�k���ܪU���4X��iW7�Ȝ�]�*V�LE�Fy��7b�w��1qu=�A���r0��������;�(7ޗe���9�n.ȅm�{�����l%�(�=���1�V��xIh/Mz�0����L��F9L�@qm|&�^����*���^����C��^*9)�|���,�ʌ3�	i-�%���Ew��uN�ݼ�f����\�#|:GF�q�1��K_*S�!�sײ�1��//�_���i��i�w��M��۫a���#�	����)%��f�MW�Ԧ��ƛ�d���!Cn2!*ID�L7�ypm�4�6C�����5�ڤA&�d�qg�2茓g��t�`v6N�p֋���x�uq,���?'^�[��$F]�M���?�T[i0��ݻ�T+�F+�B`���ԁ�VWn1w4�!�V�~��%��+������!�B�:M��D��BI��������J��`#�J}�א��b�� �{}v�*�	%۽*SDӲ�RI��G�%�PAV��ۺ6����䎅]�� p���~�w�Ɣ���MU���	@�� ��E��-z��ᝄ!�Dۣ��e�����v2IK2�U�h��5���i۪?���z��2�q��f0�2��Q�ڧ))$���$���ͮ��2]d��CD0��
'�!�a�5!|[��LO���3l� @�I�Z8��t�s�.��[y�]���x�7�6���I�E�I�.h[�ڔ��'��g%ќ��ߏ���
՛�q㜖�I&�2	i�˚�x/�?ʛ_Juu@�	ZF���j�OG�7Ĺx_� ��GCI!�$�x_�Z��|,��	����q*�/�h=K�l�'jg�-�̛��]|a:�J2Y���a��i(�p�$rTN��Z�N�÷M���.#[sUѩ����p�uc#[�l�UUUU�++@J�UV�*�o�I�cv�Q�;[:���p���[��ۭ��),'�m�{�-EBQ�!�A�L��쐟(Qf�A,��Hĥ�F��턬XsWdl;�$~$���>��'����
��>��ʉ)�j�]��0�4*��A�tT��$eg0�4�!�Ɩ�Y�T$I�P��j�	��?i�a��mD��m,;U��n묊{~��2)����K�_�Ò�!3�B����6���L¬������l�^L��2%�t�=m(\JU�NR�j���SA���w�o����J@��H��d�Q� ��H2]����?" Kz9�J9��y���pJ�>�h�����Re�)���u`[��z����=n*�7ta~Mr;˚f�N�rL�!�j�[k���R�y��m��41�	�E^U�N���~#�BM�O�O��U�j�H�R��~	5�lt����vn���z�&l�;:&P�^�oT�;��\�F�$l�$����Խͼ�����b�ў�'�8����9�S�di@���-����[1��i�!l�DʄT�h"�T���n�������&맢��>h"	l$� _.s�$ˀ��(��2�C;�wv�i)�u��ݫwIJ#��v�L�z/�!X�n��֐�qnS}�ir��VbC��HKp ���T�߮�ÇЩ�%�;��ԇ\缄��@����Z�.�->U]8jƝ�ȱ�;�R?CI������'�ŷ(��Fs�`�+��v��c��=��	�烋7kO'6��౷#�F��k��lݎ�cs��ے��+�M��3z,��ۢq�! u�vI��r�kk��U�.�iK�C�8���R��h,����uh�bzy+!�t��"�AF�F�Bw�.��w~�Oj�H�Fm���M��nv(0ˁ�W�V��)�c'�c��SM��y���/�	Ш�z��	��I�Pﲣ%"�{�Є J�O:3�e���'�����}Vɉ�1�5�`�+�I����e�$o���|���m�ުeY�@��&���r~ۢ(�i��O�P$��M�.c�.�Tc&���]�Bf��OȾ;��W�r�t��)-�2����D|��n�|�L�m��pP,@B���~w�ZWʳ���P�ՠ��	���(�+�.�d���cN�	!>��
�3�<!Bj4@���υQ���c٥��mG��if�����{���|�><q��[b���ձM:�7�l\�x���������I��ʛ5���͇$-_";A����?	�#�+7�����2~x0�ޟG��||E|��5݅]7���J~0|E!�z��;}�B��N��P�^1�bŠ��Dń{tc�u�!HH_?}��i����;���OL�lͶ�6+�3+��e�t��u��[v]l�q8��� ��AD�����J��J=�&!�8@�F��Xd�BEC	??-��m'Qj^'����n�e�	׶�:Rb7"�?����PF#�ʁV�A��z >�y��A�9��u�	�؞�K&��ᒁ[��"7~�\�I67�o�z�l��m��}�/����
.��*s��*���t;�Mշ<��$�f�.`��	��a�#�"	����z��FE��4�C���J$ۄr6�28W�@��#I�3#'���۵X	�p�kzn�AiC7o�C'漑sF������'q��{�!�%!U��VlX4��f�P� �[	����(��)�W �_�^��=�~��Km%��P�n�zҡ}���|�R�^f�"7�s��ښ-��E_�j������{P�p����pȣՈ�*��!T^�m��F�N/Y����h�b2���=<���p���j�L'i*[�=<�L�+�A<=��V!of�4k�a�!]7�D2�Ef���wՆ�����t�-��E)���%#r�q��!��W�v�u�Yλ���f`38cJ����r�f�p��M`3t���,(��R��Ku��_yu{���o��E�O�e�c��UI�`�M5	H#!����vWs��u�E*H"]p4��r�Q����\0У����2{�*g��">��o_��^�&P�=�w�2���*�Bh	��e�!u��6�v�}�-���D@Q(��s��F ���q�L@R���p!t�B����NABH���4%�C�_(��K��T�#Q��L��(���E�i�0����gNsԋ�*��Y�ws6��M~r6�%���f�Z0��M�)
@ǱhD=������c����D��cް�Q��p�H���ʩJNW�@%�9@���K4���'X��"���=�z�wďW�U^���Z�+��e& W?a��L0Yv�H��a�f�f�rQ�³�F�ݛV��.rW@����w�#�'	e���n�/A����
��`�B�֩�ss{�i�f�I@��r|ۄ��suDț�4�K��w7�Q���?(��$;�!��(�Â��[ԔLϗնTdJ�8h����Ɛ�߭��O�;5�Z����%(�ɠ�$:�.�BpO�YA ���Rr�qS���Bb��B��*L�'�G��Iy��r�������n3�+�������@}-�T��pR�c���vV���.Uo]���KC�V`��JI#�r���sz�dq�2���wdy&�Oj���(�,�ᔎ����G�jً���׶m�Ō�_�+V�t�Q^z�޲Y��7rO��:�Zѹ�ې���,8�aK9Q{u�%<�=�Gu*w��E��_wd���U�ݖ�N��D�[�h�4+��$��(>�yԏTN�̬�u��E�]VݡR�"��ls�Y�;E���Em[ 覍�K���;F���29V]m'���ev�L�O��喝{��Cj�{�^�)���M���+x����/sb-Q<�M"����1V0�"��V�iL�v���Ajֳ�s�����n�9ie`�U�-�A)x��&}[�wQ	n���k��<�����RLv�̪�/M^�:{���8Go43G�aj�}�#U��̱��]��Ē�ã���:s+&��$�I$����kd�i�����Rڪ�����X*��mT�UU*�UUUT�9j����R�dpZ9ڔ�Uk�;�j�yj�]m��(B�(	AҫMSUUUUUUK����������T�WTک�UUM���*��5U�UUuUTڮ��
ZV�eN uMUuUU]UU6���ڬv+UT)Ɔm�`j�M��,��U[T�r��T�����9�UU<�T�ԭ]�VT&��YSZ\dW��՞�lѶ
�B�C���x�����������������������������z*	����%��*�@�UJ��UUUTUUUUUUUUUUUUJ�UUUUUUUUK�UUUJ���jU��Z�7�e%�Ij��5�HEv�]UUuUv�ժj����D@�!UN4�ɽ�5���������&�U��V�*�[$��(���j�����˞?��� ��b�'�$9�7ZV�����TĘT�l�G��	�#��=0�{���ث�?E�]G�? �f��.P��Z���[[���4ȫ�I��c�9���w#�>+�g��(�A��Ud-�`bU�st"+6f�P�:��N"b�5L%{]����Y��>����kΣ��q����(	�AOY ���OL��BO�P}(v�ˈ�
�1-C��o)�)����բX<"[J1.u�J�۱�4�D'Ůr�=�Ͻ4�T�$a��<9�C%lq{��*!�%���i���uȼ�o4k�$�a���;��hr��3�F���D�ٽ6; �����%phi
����p.�e=��t �P���/n��M��J���m�k,%����KZ�SmX�)�}������>�<�^2�A�73�)x�R8��\[��eR�ld�G9b @�Lp*f��gn�`�\�PFb&˒�$�r$��g�d�ض���=!,9;�7�xDn��\ }��ƨF��!��v�'�dj���T0o�5�o�R�!ۇJo�&Y�')<ܨ�E6�Q[���ul���\��c�xc޹wj.�z��q{��t�v5a]�XM�KE�w8�r��⚟;Ҿᥗ����T�z)Z�g�:��r!�]�CX�gr��IQ��ci��a;r��݃s㳮i�Q�欻.Zݳ>��HC��=<`�sTlv\���ּ
۞n{e�X2R���c>����6������
��I`@�b26E�ds=��R>��Tz��9~��Q��WGW��QR_�6���χ��Py�H��&�.����$;�_�آ�b�Asg�E��4�zW��c��S���`H9�^(ȋ��)Á�<�Z+�ƅ����9�ϕ����r�rQ"=UGy�Ƨ`�3~�ro�I:�ۗJ��I�h/�����N>Ic�,B��Тk�0���W��r���g�.P(��dX��u��L%��K�Ĕv��/�}�L����c�+���ԫ��G*��Ѣ�0L�wr
�o�Iq���>̑�9��s$�T#D%H.6n:�&#aH�]"�x�ŕ�B���3��D�ݏ����3�"�nI�(dJG�'cG�����<����2�R���w
�7�.�q��j�\9��,{�����Z�b��i��6�Yw�.ٍ����g�=(?$0�����P��t��d�UU�0:
��$Ͻ�(��̤"�T�+up�(�[@�&�WL^� ��P\_����B���]8R�RO�}hLi�Rg�%г>7C*�W�U�q��A�w�s#5Y��������W~SfH���`����',��i��'e��wM�C��ǔe�e YGA��3�feλ7�HQ�ț�>^b�Pbݽi�H�#,z�UY횽��R���2�G��`�4m���Mz��[H��<������2��34��)��5�B0N��hu�]�-����K�a��7��V���7^��UW��Nu�s0�O[0���^R�����&߆�-���ԏQ���o�[�GG��t{�)@���u��&B'�(Lm_JR�ߣs���j����Q^�y�Ģ�aS��(%�p��P�"��>�?6��;i
�K�0C���R�3A�"=p�cX������ouv��}�l�Q��,�ٺ� ǈ��fþ�u~s�Q.�����E@��-�7�1r�ee�Eg���/>NxS�;�I��-�^&$��!C�nn!����@�7��/w�:��8U5'T�W@��O�mx_؏�݊�����@��,�&W�F�]gŧ�u%*6�DB�O!D��DL�{���m��r�
��fu�&ŎV��l�`�i���D���r9�n���{z�@�)j#szQl�QvOO~��]��� x��D�B��ر:j�H�n�������Ow^J�r�=.�x�v�+	y�-�z��6��o=l�����8��`Axr�ºxA8dI%-AvJO:���^l������te�+k�L�So�Nϴ)���8�s�zcp��,Xn������'98���ۣ1:)I!OlKu�,s��u�~�"��LT[=�Hx�w��t�DwM���8a���m��)�Q��b�B�_�EBI��ߖ�*7���a@�K�X��L��䏺�@��}J�Ohu�{;O��a�J�Ή-�A{eވ�����O���@��2��q��TC��zz9򉻸�h�r��7�����$D�(w��TR!j��jj5[�Qֆ��DȘ�?�f�뮧����1��m��~s�W��O�i�I�z�������>��{�[���]~P�_4�6�.s�}Vu�ߞ�nT}��}�0b�W���?s�XӢg��$1�'Z����q��ky�{o�D0S����U�&p���퉋ti6~0��#�ދ�ĠU���n����}6��g@��u�u/�m�}�0m���f0⑤�m�!���˄F.����m�uU�j��v��.R]���0��a�N$ �����e%�UU����U�Y���o�.eB�����%��B$_��� 7SH��VX��Ƿ��&U�*���f�uh��h�
�_֭p�����6��s�a���p�`��R�\���{/�x�߳�����g���ztW�<�h\�uY=Ui����$�I&�O}S�^w��!9¡�}�~�=�4��*�?M��QV7� u�����R�X:�������q�p��t���YIݱ
�"h�翉�w�>�M�)Ɗ��!�������o�.~m�Bq=?�� @���"?8���̄�df@1�9����/�nƟ���\��#�Kɉ(�bF���v^�#73iBZ`�<�D�����c�A�6<���.����,�W���V��V�(Ȗc����V���=m8���D�h#��j1J���q�V����}o����1���c5���&2M����}�!R܈Md�9�_�xè��#hA���gW���"To��]Z��xb��9^W�vB>M�
RN�)Ź�v�s��̊����7����t����jj�%�7���V�m;v��8����M��=�^�ۯ<܅�wl�D�\�N��Sb�ٞv��5g��	1��� ��8<��m�uқ��c�(�ja x+��ړ�7ny�.z7�7b8.B�-�J������b������ȶ�i�q�����rL�q��%$�0�5��zi�3�$�n��ڑQM��N�7�R�ʈ=�o�W{-j�7��`��(�?��D@�����\2��G}�9��g-X�~
�/^!o3v�U  1��5$C���^�;e��L�o㿟��{غ��Ӵ�ͳD���͈7��ԋ
^�/��i��oOA����pԘPXO�%	+�ȭ���-k�:�z�9�f+g�����B����I�q�7cT�C�	��S��T�ɱ����*&p�9V�������N��Q�>�o%^�u�K��҉�������9�����[e���$ђF��F����4)�K��9��7�/�yFR���t���)#^<�lh��=�ٰ�a^\�m�IEJ�|הS���,�����1,�guE���ر���[=3�A�3���D4"��YQU����V~�âokh[��t���	˓�˝{�E��2�sde��o����1��+��E|P�1���D�c�'øo�`���9
���3��ݷP]n��19�Ha����͗���5���L�S�N����/���7�]п�*bT-��8����j5/jd~u�%êt��Ö���ª��5K�e�y�V�d���$��J!:���ɎY_���8 �����pI�D߂�C��s/��P/jx?�Q�!���>�����n�6�S~Q�N�a�)h'w���ܦ����}�Cc�u2Q���S�ɇu�k�&���(�Dg�1�}�2=�&E��.�M��w�i����PwW���w�a�[hU}q��Y���Wx�6�(%�^?��eת�[��e���>R����A�Z��7j��..��Ҫǫ|��v�Ζ����� F��(�Mћ.���wn\ճAB�>̣��`.UfQ-=�syF��N;j"�X��6]F�3($𸒧����2�|���ױ���D��x�L��l# �%g�x{�}n/s�(��w��F|�T��̸pf�to�-�f����?du��=8��o]+�n��p�5�x#�c���l2B	�`�)�yv��5Z�[4�m��cP"m$�Cm�J,���7����G$#��e�̉������Xы�~5{�~�n�gxuR����c�hAXP�A�L<xrm�m�w��3gs��TLw�.�Ǡ�bƏw)th���>!m\5A��3��غ�Z���*k=;d?]�B��fl�P�#�J��+ͨ�uG���*�wJƎ4���p��}�h���B���I>�Q��sħ���Ir�f���d]2�W�r��GstOq`{l��u�����M1ח{X���K���hɂs+Y��غ;O��C��n �:ti=�N2�I%�U�{_&��]�o,P����u1~��e�J��4}�%�����$%����*�y9���]�Fm^�l$=�T����*��n�]��L���":N�{u��'�m��ͥ�D�|�1�ܒ6�nI|��h�ܳZ*�u�m0SU\i��ګf��S���n�,� 5UUUUn�@UJ�J�U�)-C��ݲe�mCZd-�m��a",��d,��1�6��xl@�}����#���zyG(|&$e�u�(罰P;�l���|�ި�m�IH%Wӂ�>�W�70tdׯ�|�P�Dh�7�?l�BA�@��6va)��	A؆!�B���2�c��|�"Ϭ�g���OV�]L�ggv�N��F+���f�K�H�A�95]��I�Ap���u޻�y�	$Q��Y��xtF�M(���ֶ��Ϗ�p��j��Ns�PA!�C���o]�aZ�@aՏ۞�n^#bG����P�`��{����eU
����<ӑ0�d���$��n�\��1��*�wo��rf*;l_��b^���G
V�tܯ��^]��#��S2j�͉�PtpFHO��(��d�X�Y���#����<�HP:ج]2�A�Gw|*e����;��9����H����ȣO�j��}�M���bj"j����$��p�{�y����)��K3m�G�I�پ��n�}�.\0e`Y��Uf^&��ắ����l}c��8���'fki�g�w睍&�uv-�4���V齶^-"���A���.۰X�K���wuM��`g�B;[��.�Xڔ�6ݼ�����P��j�]r���jn@p�N���v��������WQ��;]�ٴBI�Z��:�������' �)|�v4j��YB�읁����LȭK���M�b]1����Q��+j�v^|c{�Ti��;��L��x��s_�[*C��n��`nd!`ϝ&n涵�MA� �t�d�G	-n`�
	62��Q~���3�9�z��l\�� 誌�|�G۱�4�s⎿�����Y����D���J������e9�$*��{U�!����ۓʶ�L�Vǃ�py��Us���!̢��f=5C�И�\G����FD�b)f�R��!��y:�]��2Ǒ�\c�U�w�~��%�mn:�F��qу����p<<�ʛ�/�S7v[�rB�{�{+�r�L:���yksD�y��v`=�?+��ʮ����Р�58����*��0�JQ>$����3yer6l��_]O{�1����<_�t��{�R�?�;:��ę,))���k��mY�����������{�:{��4�䚻��w5�V��v�����!)�2��꼰��!���H7�����4���.��4�5ɽ���y���2Pˊ�/�iN�fWwMD��:-ҸR���8��uD����lĸ5]�M�C�N���1&nv�M��b�q7C��c7h��_n-X�̠�}��c���V)-=�u�}��]�*��^�x�\g.�9N����t����J�͠��
�l�t:]�q:z��O�uW>K�W"ܣ�>��ڥ��۽ʚ��Nν���V���ܔ�泓c��Y�F���g�����6�@�������ͽu7�_ܻ9[u�u6*T»R#Rt���hm����ǐ��z�]�y�=y[5���SZc�U�7���!ۘ�}�+U�<���ۤ�̳k����3k={j�y%L���k`7�i;?��>e�)����&�KUUJ��U�U��"ʮ�3�$k��I�9�P�c:d4n�<08��uŸ�rڷ�\t\q��ܵ��+��]�!�7j�솻Yq�reƮS����b=�y�k��n��\�d�����q���uk�"���\(^�T�ջt�dS�����쩆g�f�J�X8��8ʛr;�n0#�]Oi�\��7�=���
����J�`�mݷ3�y��Z����<q�*R��Ee�.��0��c�j���ŷ���v�vT�y�3�Դ�;�Ńq�[��^ؼ{֎��q� �9{ɳ[�+۷/�=��s��I�[���q��<��|�)��u�m6�`�w5��b��Uҷ\'���8÷mu��d��{'�ۭ�t��{c��N;�iO�]�7[�5���2��4���i�ƶ�u����M��*ވ8y�{v.(��ݟ���������i�[���6��S����8z�m�:���o�������q�	����nr�;��d��s֓ �.���\t�0X{k>���1�ܻ�88�Qў9�P�s��6�E�Rwc��X�7��"����<t\%��ݱ��������8���q�ݣv�n�s�+�uӽV�B�.92��n۠SwO���v���~���ł�O�;A�ǻ��
!�}������=e6��������ԉĠh[P"�G���1��e�+מ1e���qB���V����D�#e�n��>��ܗ��D�~�^f0d{������ȶ�%_Y��V
qЈΙD�=�wt@���f{�`��o�g6ਜ��?By��E���/z��ɵg��ޖ�Տ��@�
QH����4K�M�I�(�R+�o꥜4�7�.�+J���g7X��9��.f��q���D"����	"�GW_g�&��d��*��]T�����#�s��qw ���~[Ǻ@��ل��<|�'�*������1-Kj!EǨ{��]�"��Bj1�QDN9�l��6�&��ʞ[y��>,hFBx�]�Pp|Xi���l�ޡ��{0��ss�G�+���b���ۧ�ڳ�i1
P�	�FgJ:��^$�{ʩ'3��H����NT��t��Ʃb�Z���Ӷ�}.�t��5T�	}N�p*�ͩ���\��5W:%WRᬇ$m~K�����c��}ջ��=�tT�cG��_�&�~��ۃ`�tș�����G����ylBC�=a��'u��k輼H#"T�����R�g*�r?���pNW}
N���DU��^��[�,�5���j��<Σ�Cxh�cbZ!�����~���K�Zp�{����]�h���@y֪=a�l$w��Ge��[]�-V�B�F0N�M8j,'�z2x��"橆%�s��+�fU��{�]��Dz��C�s$����Q���_{�mG��^��l {�f��;\�!�\�W�1�UH�ࣅOp�����[8i�7l�q	_4�d�^�˧Q5��>C�F������#�{x���ʆh�X�{R����D��I$U]���1{��;(1\9��b�s�e��ۏ��U�m˻�VL�9��򞉗C��R֬��^��ް���Gߪ����t1Y/���v���{�{����5ރ����3���O��;u�+K��p�Q��I$�A]��\c-Ӯ:ꪫ����j��*��7l�!+R�4���A�Z������*!.j���VXj�,�[A�صK��YVک���HX���I<:t!�����ߣz4�d����hja�u�}�GG(P�ߠ���B�M�r���ݩ8�1w�f���1�\��Y4ahk��P	�b}��gU�O(����L �&�����xze��n�w�}�zE��9����N�劲��_�t*[��#}���<��]���:�%AJȏ/y���-�ف<ȁ�z`�w�'�E�%�)^�΄�H��Ү���������0y�{���\<Gu�]׳�Pv!R��k̹v{B?	�������Շ.Pi0v�v~<�v���'{gb�Ѕ8��#��х��f�y���$5�Bv���ͩ��q/������Ӄ-4[p#��I��	ȵ\�׮��d�ˤ3��W������C{�E=�O�U�K�A���nM" ����Fv��o�c�J&%#ʆ�B���u�]{���=A���5T�d�t�T��zfe-X�8F:��4ʷ�U��d�4&���Q�d�6iX�n,��u�L.�ۧav�@t��.�;m�8�f���nN%��F�q�n�
n�ƽo.��v,�k��x.&��a潸{�;����z�Ճ���M��W2FB�ݵ�"ݞ<�i=��N���l��e��ݧs����_������"/��1�~��t>V!YR֡��<g���7Y�_�+@HȤ�vD���W����u(���n�Z���q2�2DrT�y}�bl`���8��q��Y�H�z��5�ԑe��m��٣���*�T�=�I(�)!Bٹ��n �ʹ�m����;w�ND��3Z�dN�{ޥz�7*�'�UN�Tk:5}̤�(���U[�P��	D8��w~�{�P;!*ȉ~caTF�˧�ܣL	��7�W�'�ۖ���"��G��u,�(tm�.�_ϐ}�w�Id�˻���K�PR�gkre�W�׋�� �����owL�Y�9A�ׇN�G{��5���"����נW�qo��H�|8��K �舅8��F�����4v^2t��Φ�Ϊn�Lⵜ�m�	%�;K�(Q�3�/M�"zo4�����qW�������}}��GbGv;�a�\�x4L�wZV���A3�:�>�t "��.�Ayl����j��n�w6�ta��Fn�X\���V'�F	��}�?K����."`�F���ذzb뮱�뜌f����BeB�8�Y_u.�W�b3���m�AY�;4\�g���@�a����\?L�t/�a��v�����Z���;��-�xQt;�ϻ�\�x�1?w
�������WX�ECp���3U�0Ow��o�ϝ�ڧ2q�5UV��L������S�\S��9��ݐ�س�Tة�>�54D�e}6`L�g*�_�yA�4�9%M<S[�3hSh)���{8���]U�eP!fs&.���ǩ��?(�[\�Fw(�)�74s����7�ӷ�jc)��"�{(�v;���C��^Jӥ�9�q���;��#��!�vP�N�8��	J#��u[::��^�f��;�{�^�s�f���[�;�Ӂ{rAI8D�%�O>�ݴG��G�`��ݏQ4�����?����ՠ��W���+Ƥׯ��o��I���f(X�QWyUx��ڼ̜J
^ym}��9���W�D�]V��ca�w�\�:�읥��%$_���sһԢ(G�Vfz�^܈߱@ـ�׽
!����\a��������|G>��gk�[]8j)LBl�-p�g��ڹD�lnF�p�W���j��(/߻��y�"'H�� �Jy�اU���e������^���?h�����ҡ�!!��zQܭ�B�5����=s��7`j�L��ϐ]�~���O��5�W��G�n�d�^�������r�7��{I�%}S���]���Wh[����
LF��푈t�5ڭ��s�TEK�Y()�B8T|�/|	@����F�D6�����}be)E9B>�������	Wy�5��N�n���88Hw�z�^O���z35"8���U�V�THl�e`2c��4��W\Z��,w�yU�5����m�oe�s#`B����K�o3	Ex�b��we`Xz�}[Ym�	�E[�oUE[�A%E]w��/��2�7C8�gv����_����~�"�V��(�b���6⪻j�(��`.����%�����[��T8��6�KUUUUS� Lb�U����
�g��S��Ŷv먂u4ab$�l��7�6����n��~ �B�md��>�"�w��x{���PB"��o��g���r���v���V�*�4���}�������Ų�#l�ޜQ~}��[*� س���R��e����i�kbZ��G|k*��F�g��{��;�Y�5u�\���ru�x��uh8�͑� д:�l�^�o�R�EX?L����lzfT��Sf���N�'&E{�=��M���O���$�,A�K19!��O������C���u�K<���*窑�D������t���� ���`�py����N����X;���o���ɷ�Gw�du �������W��0Y�e@��݂&�ȏ�Lջk�?�e�z�f�L��:Nv檪ک�z�����C�S�*��RU\L(���%�#ְ���F�s��xc˵-|Q;e{Y�
c�������,O�+$m�$4�����+�˜ӯ�'ڲ^⟄�\���q�����6~,�,+�)Ɗ��5w*j�����[�i��I:M��9$a�#Z9�7	Xݦ���v�M�kw����ghڧn斓>����jƳ�{iIx�ۤ=�J���uy^�nQ�n��`��X�E	)��9�
�u�����f�04��4�;Xέۑg"
o-�'��&wz{}yΌeи�GK����y������L�aJ�h]�
-�I�:59ZW�y�}Y=�I�|�k5�^��������h�ʱ/C�_�_��H��G����	��M3.�}Z��	sæ+В(��L3$�΋��Ԣ��qu�=������B6'�h��Z�<:����ﻸ�ٺo\@{������E1U�e�"R��V��߲�}�p���[l5hdm����h����=���x���-��PQ�O�Ͼr�LW5�GXU�����>���0�zEj�YiXl�����ʗ=�D_��Z�;�h:���A�
��D����;N7�;cQ���3η�驥ĩ	]��E=���i���D(� q�Tw[̂el�؁�Ev�#n-W>������NBF1a����˨o$�\�01،�~���Ӫ��#�>��d�j�ݦ1�Ʊһ�M��N�����{�ʸ{��0ى-6�5\����pf,co�S�<:�N�#&����̯��������sD��Q) �bz�d��?����n�Z9;�ıJX���
Kr�}���WPϷ�Ѝ	��$N�)�5�o�r"��
>���oKL��~�5}�UP��\�1_@��z�q�P~}������LI^#�G�N��
�}��I��U
5����������vWLb�	Ԓ*!0�A(Ϝ�ݯ\��v��{V�"+�Q���p�/ϝ�"�7f�Xv$�S�V|�`9ph�$a�K���tQ!�Wt�[�E��Yѭ�/��T^�Es0w�o��:�$[����}�zc��)^�#���ji|o_�8��X]ڕ��m�y9�����a���K9�w���!�K��-|eZ0�|cH��V&륣l�Y	�`�&a���_��]��v���FK{c� �/�?E��~� �2�(/j���}Cup�	lQ������>U�A~�@�]�c�T+���%Z�h:��7���}��q��ҁ�Q&���B�;�C~�b��.�$Dk�Gp�	���}c��J���%�I6qO�C	5���;���Ԗ�c�A����#"7>4�Ip��9�5��9DͰ��i(�$'$�I$���&!-��~�a�Φ���i{��}*�~�'8��	��J�����F��i
??�9�!z�6;ާ�SӐ����?�ۤ&�N�{��dW��/�ӛC�{�Dd	Gu�ofgE*���B����|�EѺ�1ݘC5���S��.�oph���|3��ؔjm�F���z5�W�����o˝������[��A��&AbD�nR�˽�^�Ê��aQ^��ޫiw�� x�t��G�?5��j��lf�Y�p!,z���^�!�Q����|&��/Ӆ����w�P'D��:b�� �=+��HrXm>�A����,愲��ö��`�5�6�"��*$�j�櫬�3���&�ә��L�i7/tmV#�3B��(-�b�b��l���/T�"���#q�]̂�8�P�X����kt��x�hl�C�R�����lǈa�ֱ���Ǩ�n�}WWo��b��-!er��򴻮��r�f�hf�����VE�i����b�o=�j�[v���x��N��$[�)�Oxu�y���ҭ�Y#(��5;�k*f��ݕ3��M�F��Y\�ܡi�t��Z����pwMϺ�QM����:��Mm�ޕ7~��m���F�S��z=�u.\;f���F���II��Z� �欮�{Ԋ�D)y�FN�/��m�R��[/73�����v��u���U]_K�O��9��j-���N���SY��U�쬮ʛ[՛��AU�ڽ�Y�U1���p��:C3��֭fo.�*��/w(bG%�ξ���n�F��5���/�]uU%��L-�|2޶��5Z��o���o����U*�Ui�e�檶���	���������j�V�������V���e:��Ciݪ]���LjqGb�tQv����Rnˈ�&�gtJ�uUUUR�Ns�5WUUM���UTV)��5U�UUuUTڪ����SU]6���VyZU��IJ*��5U�Z�^��F\b��i	&ݚZ�	���R:Wbڸ��������L�dU�Z��&��/-K��I��k6���x�kQ����H�����`'l�5UUUUUUUUUUUUUUUUUUUUUUUUUUUQ]	A5UUUIQ5R��hP��j��j���N&�����V������UV����Z���j���V��	U����Z���ϟe��_>�ꕕ���Z�M
hYZ�:z궪��\IW�����K��+kW5l���Un�j�����jY%�j���ڥ%������A�qd���)D&ۇCm��;O�zZj�j��e���p�C�J��ip�����{_�h?]\0�/����Q�H��u�dh�u�7�5!z4��F�=��}w�]g.E�Q/���x7�z�YlΪ�s���FE�(WP���]{��Gn����K������*�vk�qؚ/7.	��0\7�Њ�̨�F]�m�v��t��EqF	�'D@�B��V����8�����4ߴ�3�a�2$@_{/F��U�N�,/xU\hh�N�D`��Wx��ggQ��>̰����A�qV�÷~e`^�k;��z��h���5������K/�ֱ,9�\�O�	;�qd�/h�;t��#[J�V�'C�g�U����u6�ܨ��
��a��x�����{慼ֿL��o_�@�zѕv�nF!���ݏWlT�Q�;E�)w\U�\����ܞB5�N�OA��Nǰw\�27����ϟ_�����%qN���#ˊ�p��%�O$P�{&��s�n�iܡ��=�[v��K�C=��v97t��7%��N: �
f.t�m�4���n����{�� :��p�y����x96�����I��̣�u�֡��y6CMؖ�C}��"{��}�3=�BO��a����͇P���UMy_pUp�M��=�wݛҸ*��P8.�3���ߞo@l!ft/\�ʭ�	�$�����I��c�a�j��I��O��A�a�X���RCϐpB�2DZ+�5.�Tļ�bC�##y�U�2%�ܷ9oyc��j���ȟ"
R�EBIl/woc�bX�t:�3b/i�����(�Ǯ�Dn�����	�Ĺ�Q�dl ���/��\��Y��S��,"[mB��@��"c0Un�k�m��g��_3|�ֻ-�7��0���a`�x�*�i�t�o�4a�Ex�W��'������f�4=�jD<:y8BN>���<�F*[���jB)���!�����zk�����ﻶb�����38��,]���i�B�˕�e��+%�������ݴ�%�3xJP�ݳϙ���{\���w�O����+z^�ǦD0r��>�=�,VDe�aqDn�V ��D��u���˂�<�ڊT}�߹w̳Cop���P��+�u���i��sи@c<�y��y��#e��^��zxr�e>�9tY�4�y]���Ʈ�%^K��Յ��Tf�I��!��gߎ�^��5g�湮�[⭶m!lә�r""�VV�G�����z�,��^�Lp����'78�-�M�
T&�H�(܅���UTvt�8�qϊ����V�3�X\u�l��1	��'�Sxg�T����L��W/sv��ᇳ�@�j�4g	�;���e��||�1�竹�5m�r0�!�p�9k�h�܄�@����__x?ʾ	˻�D~`w(s��)�a��.8��;�Fmq5�_!Aџ)��B�X��H��A˝.-�/�e��n��5	mk>[��E�m)��z�!�%��I倧������0�4��?�C_��CC��P��<�LX�E�'���BR|���|�+7w���ʀ.�}���<�w}�����T����A�v�xY0[%������{�X�ض�z�5�,�!@�z{�;]k�nS���X74����/�4�[����)P[�(�_l��K�sοf�k��_�3~=*w��4,����As;ӑS��%���r�FbqD688<��%q�Nn��v��Rhl�X����z����6⯘I��x��N�����$0�M�M�_7��e=�cD�&�,8�2XM�nZN.)��\X��7l��{��G��E
�1�VJ��u�6	j��YD��2�;d�%0��阅3,��m����ߎ���e��h�pna&�Nz�ZPkX����X�m`YZ���j��o�EHTl�j!U�8���5��œo����;q��1�L�{Ľ�ҺT��벻>���%��5�q���R�UUW��:��U�MUuUu�TQT�e�3���{EUt�]!�ƬCUUUUUp*�M@UT�T�U;f��4���j�ڪZwM��_?w�����'�|*U��+TQ��a{52B�]SCӰ�+}W�s|wg��[.���A*����Qd9��>����)R�t�Ξ���ٟ0�P�f�:����@����1DDq�,Ӵ���tr�6xY�^_e���,�/=�ݯ}�m���o�b�������3k��WW��d^f0ߌE���R`�>�A��r��B����T{\f�5�Nw4�h��8\1�!m^{�7���ގ��Qg���^P��t]���7/!nmuD;-�#
0d��p���.�`p����	9���K�5�rd`X3�eo[
�nE�����׭il�̙g����8j���Uq�f Q�H�\]�V�vj�$�}v������9t���*q$Q�?c���W�ߕ�c5��
÷<��ه�2br������Eț���v�x��z*ܠ�C���ȥ�#WV��AU����q�Q8[r����a5���`Q��n7��9�RZ��G��h�{]���t�Naڭ�cnsϝ)=f����lT'&�vɹ�����{<�bQ:��E�2��{N�m�+n}�z0�J�,-q�:��Z4��ڒ�G�Sb9��l�?����)&ځ�������~>ɕ�WA��,p.'ܦ�B���$r!�`ȳ�jW)�M�w#,\��˳V���h���y���`7��3���y����x�[r�-�;�Ǚ�Q�H�Xڵk.�䴑,3d���BE�q7=���fΨ�V�w���݁������t�����������f�Ʋ�)�|ڍ�c��X�Fg?-�dh����^۬�S�>�+©9�K�b�S�՝�MY�l&����\Y�9�����+�$l#��j�u.�٬ߟ���^�UҜ�j�_���joT��w J7����G�&P�z���l�P�i����Y˴�sYE��'+�3I�M=�
v"Y�=�Y1��vЅ�3o���J���M����W��Ř���ʫb6]�Βy�3���.@��z�&6�"�摽ʷKh�Uf�����suc%��4���O`վ
>�zz��/%���۽MҠ�)#�|���U�q�v��>,�-�{N�x�цjܚ��3�e����I�тwhD��M���rB�{�iݴ�(���СP�$�$���M����3\���OM�_bǰ�l�g{a��}!���kwh4��r3�!J��_Z$ʰaD��N5��٪���8.�go߳���o�����(:����C��m!X������x*���}F*��<��HZC���5.Ou �(
"#/��8b3
�����P�i=ܿ�>�iS$���f���~c���*���Rf�ڋ���2&�z|��¥��krDw&�=�<1��;�,$�6��Qo4W'6ˮCBܣ��Ib���2����O4���.��- ����gM��u��z0X�-Uj�&�����w������t08��p���c��g�cY�N�p-۸�VKi�=���AaKltp �����65>i$��;�c�Kh�&H}^��W���yp[[�6�F_�[��<Qw��˱����0D���N���/Y{*�dQ�) �H�	�27P�#F���w��]��9�dOx���1��f�H��IY���	��3[���́�6��m�����ZJH,6f�!��+XVh�-��%�c�-_��#��X�vƒ�irϜ�������������yΈϗ�14L���\}v�t�����}ٗ ε�qQ���(�*K̩e\M�X{3w6�W֪����I�X��O'-�ivyin,�cE�[��@z�Gh��Ѽ��tP��I�����M�#9<�`NR��p��}�E��90,�q�z�NT#ׅ@q��T�y��]�U�9il�\5����{��VTz��w �����"Ap}�������Y{�䋚��p�n��7{�5J@$�H�"mq��n���WQDQUV�]UU6���7+�̵�*���Y�.Z�����ڀ�j�U����P] ��

:�f�E��I��� �>ͣT���Rɳ�
!�v���N�bn�e�3�<*�G23��#����Aw��)~VN9��1A��47��_����� ����,3���~���;�>�-��,�g��
u¨�Wv+�="`��H$!\�{i~��n�ʉ4��gm���ޮRN$�y�`G�0{��U�r6�)�_������tr(�F0�i����E�^�8t�]�
�߷���1���cr7b$m���I�^�a
�8(�,JYit�fpˈ�)�J�J��'E�U��^�C]�6��u��L�'A��^�㔏o{�Q�E%-{�%���w��j&\���(7"$nH�I�%B��k+]�.�Gq��N3�4f\g����x������C�>�ddIӄ�D
�j���Q�ٻ�Ww�[y��e	�w6��<�vl����Og]�9�R�ѩ�N�{�FU���GUdq������Yy[cL���3�-*ˍ)A��p*�
�I��繵�n�Zǭy2^Mݛ�uY6*�&�we8�)�Ikvsc{u'm��^�V�ռ�����£��a��ۥ룴]�]]�
S��q��>]���ruσZ2kb�[�te�%ӄa�e���,<)����FvY��j��K�*���rH��^yφ�߮pI������1��<m��G�{�+���2ՔZ�{����_�%C(`�}��龄��79��n�n��-��a0LD��7\��j�v��a׿���&���o�*�}}��_F�X��=���:2����;"�4*���`�d��H͗[�YB���,���¥쬒i�ˑ�����J荈�E�#n�y`I��U<u�Ȱ�:�"��V�����n�5+�U������ M�٤G8'ۙ.n+��B������Pmi<�u];��-������&		�Z������H����o��ܿZ���U0�(�=�C����C1�T��,�_Hd��uJ�++�~
�;K��Ah�/��] }�(�ĉ���Q��ߝ�4kO�Y7H���췊+�;��WPp:�]�v��P[�\���`�w��Ըg(hK嶭T�D��o����k�otf��l�op{SQ����WU@��G��D��ɧ|A���ꃈ�(�ƍU)�vVUuh}Ѯ�[��TA��������Wu����9�Y�s/$�9dG�7�U����!RЪ����{�N*Ɨon�����۷�s�.%���8�����|��=�]��"�P�)m�]l�'���}[�jY�����쮢��!�6�D��9�V{�6�v���w��Ln���`NbGF��Z�_Q�}ws9�i��w{�(WQ��������Cj�j�awwH��:&�3�T�FSҪw�o���ݫ��]e��Er�sj�*��]��F�Sb��1"�wp�%uo-��tP�yg{&Z�\�L�F�7N�kJ4ʫ�Wb��n>A��8�8l]�T/QCD�B뷻�8Y�A`��L9�j��"onq�B�z�C��t|����{��+�2W^����o���iX&S���|�p�����h��b��'`%�U|�j�j����e�v${���糮�݆^c@f�<�W���B��aw��]v-ð(P��X}b1�[�z�	�,��x,h��t��qb�\n�;v���$�^�rn�/k�4ɻq粺�{kc;��X*�]�e�tWm�w;-�v�.Ћ�,��\Ū>XL���A��gf���;r�}�^:���whz�6�{����Ny9�Z�]�27>^���6��n�.y��0�H7���`n�]8��`���b<�;7���w���Oo���hZ��_'��|��;è�ф��[dv3b�v���1�����N���p/,pBI��:iz׷�W�����sҨ<����������1��;e�;ص��Ea2�]f�rt�H��\�0mY�l��gN�$|<.q�n\��v<�5���\^нsnQ�����[��ӗ!����0c�n9�sEOg8�\s��qx�;=x�"v�qm\�����>�� �u�a�܈vqj��L		s�h�JN�]�30:����n������3h�x�n\e˺��iH���-��vw�xi�n\h�]�s�bS0��ɡ��Ƭ��xW;qI;�;q�F�l���v��tm�n��;q��)u����]�b2�?���o����;��\�����x8�.I��[�uPSrF��������������N�1�@��ˀ�<\*	#-�҆��i�1�qF���<�zE�1�qϲ�wa<^6/�s-�!I��՜1�a��>���#K�[L1�&V��'n��B��{�@�߿>ܘ��7��IA����0�)L-v�װp�9�([%�d��/��#f5JH���w�_\h_z�~�q���~�r���+ާ�h�m���ӅG<�Dc�\ƁI`��^~$^N�0;~�h���-�\|����1�-g+�U���+[��� dJ�>F�T��A�z�l8e�a]�,an["�T��(�"�R����O��g���F���QɆ�!_:����œ��ݯM�&>9ǃw ����6-�z�s�v�ӑ�Îy��3*V��٘xG��B��Z��Ac=���7�V�ƉE�b��c���[/,�뛼�|�O�M⺛8fhN�&^�n�>���5��H0(]�.���!�Rm+E@��2vv�wk��T��k���D]���$ho�4��L��݉
d�)�����LA/H`]p#0�ۂ`sNYU���6�mo�>vx�!ox10�?\�M	ѽ�����o��+y}�@xy�.�<�=����t��ԁ!�T�qs�96*��V�^�A+���9��f�#�	l�ff��v�Y��%Lrcs���}U��B00d�q�{�����,�[3ϒ����d)I��4٭f1�i����s �AxS8I xn��F�|4V�wW�
����9��R�ݽ,�ۄ͵��������'��U��U�AAG���IHV��0i����ǒ<�p��Cs<��"'�̓(%I&x��d�߽��p1��DJ�_u��0�l���۰��ܐ���<��F��}B��'���.�eb���s�C1�	���X�s7���4���m��]��Iۦܒ6�Q��(@f�PU�m]W]UU6���/UO$��l�6��r�el��W�f�Z�����JU�Z�V����[��l�>E3�`,�$��M�4\��{�C:nq.�D}������>�^�*���Vѳ�c�����z�+kQ�Rh

~����lv%�_Y�q^mYOs�,3)�A���k���:5����xl[)�s�^�:����p6�ffK��ZO��p-�L��ç|N�����#kN��(c.ez����$�$��8{�o}�f7h4nl�s��Q��Y\H�b&���pD���T����i��u*s�]��4�Ye/�n,��H!k뻴�T��J�yx�p^=���&��=>�<��f��tc4j����=�>p��]I��{/s5,qT-h��%�-�T�R�,PBg�~��M��QO*�k�\c*�4���$^�����s�M�6GF�ڗ���L���݋s�/w��s�B�Mj���g49�0u�4��(�T+17/i4Ň�R�����lA�������f3mi��Ur�f)��kε�N�}�2��e�la���r]D�WP���v���8��r���ظ�\�������s�]n�۶�g���#]��=�d�1r<����7���0\���d=�;]u�K�r����7i���}	Y!����Y֯u�i�n�H�&j}N��z`{�Tq��G�ɝ�LHu$�_�K(G/׈I��mG�^�|Q~����&Eb�>W��O>N�j1�xt�$���DF����P�} '�-�	��RjFb�ʝ}��nBť�y�2��*�Q��m���oI�G��ӌ�T���UV�b5j�k:���O�;��K����T˽a'�F�W~�s+��	,o�Ht!��P�w��~�l}}�իi� �.](��6�rBSP�A�| ���e$.Ή}֗`E�Sw:7�!��b?�>Z}��%��Q�J�a��V��:���u)�I]14î�t��26�l��޿����J
����C&H˱C�ڨ[�'�Ω����,bI��6�9tg���d<m];UcM��&{�:h�M����nA��k���@���2U}0hC�h��O�kiT�m�����F�-0f��$��2�*DD�K��7h�d*��۾^�G4vd�u_N����{��������T�ww��1#J[�7��Wv[�Dd��2��E�7+rŮB��7k2j.�Z��h33d��sq$�����n��+M����m��;pDI��#q�	r6dI��ƳI��홙�i�[��L��h�,g+��o:�@�q&��ʶ�b�QK�"
nwc��EC��|��Z�i���}�GWv�y���n(�%o0x1w-�ie#%#���s`��_N�t2��]/i�:���l�rG�jN-���(f3���6�����౥���*>�f��f�sK.�gZ{v�zqB#2���O_wa�x1=���Ԓ���ɴ�����+>鹗�r����^�b��v�����TB!�0X꽤X���:t#��_H�F����ť*��E���2ꑅ���M��z�2ĲC�GN��u̨>~켫��c5ic�!"h#mF8�%%�7$k� ���v�Os=K�i;K�ڤ^g�z���G�;u�/�;��$$�D�*�U��B��]�|�=�B�[�;ֹ��.`�&jt�)�m�2T2e�{�&����"Z�<͚r��}�-/_�r����U�����m���Lrq�����N��cjt�[���6�3$�񁯷=x��簑�ۖ.wj����f�����7�y:��r���d�nx�z�:v�U�~����l��pf�ʬ�MQ(��^��B^X��kw_Aռ%�}t8Ք�o-h/w3�.c+�u�����C�����l]VwmWծ?��Z�a�|І�|����6"�w-�C�!Ux��Ή���FےI%O&hu�$R�U�ѩ����R�����|ɘ�v@j���mUUUUU\UUU*�P
�+U]LE��8.���]�����14 ��+�F�ڽ�Qb!0�wW���0��9�8����W��AB#c8;wj#m�lrN|;xN㚰[����̫w�w�>�v^���dq���_Jk�]¥��Kh���Y��ĕ����sh~��$�:�el�nU��2���׭�!)%L ��՚���i��ⅶ�����+���	筛tm��3)}�ЯMo�⃋������Q��xK̺��-�i������2 Z6*�oy0�X$PHs�ծ=Lꏇf��u�2DG}!�t��� �:D�����r��Խ�w�~(9{��-�1�j�P����f�^�Uމխ��w��Kķб�#������f��״��N�]A?!Г��9�q�AR$�35�}�,�Lo�e�U���v�����v�پ���E��ܽu}�K�o,����{(N��6�i�D���8Cr`Z)��m��C���f�r�]����c�����H+�V�ؑ�@`��[�q�v���ъ^���GooYӴhdga�7���.n�Z�Ғ���ɸ��5s�Ws��{.{��\k��7A�\�~5��Q�
����{���%㸸�9ŭ@��s5��}����/ϥ����9�e�sw_F;�鷊��J�R�}���ݢ�R�'��lp&�plc����2F���6ՔFC	�����E�����ϵ�����3�d����E��d<����YD]��;*�x��~m	��Bd5��F�i�缥ͱ��]���o}����Ở�
_50](�ǫ�A�~�Lځ5��I�R���sP̊�¼��-��`-��6�j��/~}��쉌�+J�K-*�ξ�SNnj�8G���C!��9�Y�^�P׿����M7�6��`߱��@�g$����|U��e덥�wҤ0=�ܬ�]�V���d� �+��V͑d���;d�~�X��k����o�p��nf�鴸ƨ�"�XZ�v�|�tn��T����#�c3��`��;���H���5'-�zq��K>�"@�l0R����wHa�vں�;X�!O��6�`=j	d�~�2�,�����j�:l����{����:��8��N�b7��\�رc8���=��<�ː}DЁ��j����xU�]1�3�`IO
��Ͳ2*�Y���$X"��f�B���f���{곻uQ��ݚ� '��J�J��_>+���׹ʸ!�6,��f]Ua�k)2_�H3��z���QP��ߠ�V0�>lA����&�k�)>S#�����;��N�1j,दsv5U�ɴ�s[�����z�O���ԟ�*C!>r��[i��wf!�&[���>��v������C�ʚ!����X�2-���-A%Y�8��dX1̇;�v˜4VU��W[ܒ=��v��+�"��Bڗ�O"�UQ�w���P�Eϱ8,Q1�^;�{�4#���b�q��9�×WY��Ƣ�^�`�� �{�@�vL�)�[�^T�-X�# ��Q@��T�D�-���r�7��y���+��z������]1���/��f��F$Ӎ*�~�w��6ۖ�Wf���_<v�"�T[]�ŗZz�mSڥ;]'csl'p,-�PEYd��0y���		\�`W�]lB��T����ם�B PRH�R�җuu�ɴM�4���r#$E�y�s�mw�<WWvn�s��Q�c�<=�=$p%����V.��'V�I��4*�AqϜsk�]�P��1g�ӛGұy��h��W�67¯)�-m<[J�X�v�IA��0���i��˙ܝk��g^Q]�w��i1���Q�Z����e��7���e�H�ч���6�٪���[�;�ɱź� �e`挦Vv�n���2ԗd�Z&���mt]C��!u}q�Ź\���gky���m.�f���"���f��WG%]��5]��M�z�e���mi�֢�*��8ƾ��9��G���V�]��k����U�rWmp�/r|M�V��%[5��K��\�[��ˁe��XH����fL�q���9t���tH�e�T�o6+r�VVe:�L\��r�,8���v�N�o*n�vP�ޫx�To+��8o�����B���(�e�L��ۼnpq��5�g�8�����؟O'?��R/kx�c3 8d}*�|�Ө/o�\%�r�W��l�X�#6˱jG}���}�5�c5���J^�����m�v/
Õ��F����;�u�B��\�mI	��^iֶ�ה�+(um��#Y��t�[���ӑ�ը䑥n6ꭥ�a�q�EU�UUUUUUU"��UUT�UUT��UQEUZE�ꪪ��NR�I8��Ȉ(VW�X� �M�WPqƸ��1J	�dډ�U�UUUUJ�,ԫUuUU]uWUUY�%UU�j����ꪩ�UQEUu[[2I1T�f��T����UEUj�.;"&x�4�UR�^{,6�;R��Z��SQej�j�v��K��R�j��UU`�@x���Rx*�ӛ�F�glT6��QX(�v$��UUUUUUUUUUUUUUUUUUUUUUUUUUUU:*	�����J�ҭK�˱-UUT�UUUUUUUUUUUUUUWʯ�UUUUUUUUUR�J�UUUUj���+UUUU����|�@UUUUl\d#
�t��WEU\�UR���*��[J��UQÞ;{U3ڲUUUUU[@HJ��UR���*�ٚꭣ��)HJ@�H��yo|��[1ĩ6<�*�R�nd��n�\�i�ϳ��2������6�b�(p��
h��|s���������d�f~���ëOr)A>��$xW��%R6̗�q�M��k��m�ҷs"7�V]��0��q���GwC���˻t^CM�)wb4��47~æ�D#$�Dp�+7Os[jV'vb�)� FV�?�<q|^��}}т��y��t��:���G81&�\H鴭$��`{��Q+�TN����y� ��-�smu�ܓ#J��(�W���'#/w��ݶ�A!n$�2C E!-�ܒI�I���]r#e8�Um|��J�P?���c_O%�۵7۶�0��V�Y�{[͙��m���u��e�����+A5[�Y]	O��׷S^�|�癇v.;q2�[шX���h�%�W��r4[����M!��qn����N�y���\���sSd�0
l�)�mnu��/���t"ܘM�ζ�ڜr�<�}���tȋ��2�K���<e����9�����k���>|�U�.��yxL�>l3��(�|�AQY�fe��uo �24��V�i<��ϲU���H�YB�θ����������nS>�a����nrE���B�qĘ�j��i��4Ӈ!uO�n8ȫ(�Xc�@���,�&{kZb;k��*��qh|�������gg���sܙ�-"Ǘ�vѭƽ���Q�5^�B]z7��hKɏ�rz�U8���n��]��^Ӳ�����h*�3[�Hd��AwJ]�W���� Bu���H��6KrH�H%w�=��wm�rt{D�t>�+�e�Ճ:b�|��_���H����B��t�2 X���^�T�W��[��|W{X���'�	*�y��ޓ�_6�	L5������v�i����zr���/w��Z��-�Tw���&���e�7�	�[����v�&���X�0݅E4IG3�";�Y����W�}&dULr��Ĵ�D�a����r2�,FG�YW�z�f���n\��HO]]T�0D%��mF�Yՠ�5w�]�Ǆ�2Fs�z�.�]��e�\QlD���x�Z(�8�3ʗ�y���X�e��>�+��x1oS��]�"��k���Ήț6N�wy�?x��[^�I����f��jm����U����x����U��듷�'uxk��>��4�<����m��jm-��ۙ�J�l����݄'W��J+R�N����לGQڛ�h�ݚ�) Q�񝭅�����J(���z�i���}�Ѣ\��!��/����ɺR{��N߫M�:3HZ���J���.�p-�wek"���߯|��=uVR�ٔq�/���b�M��e�_��o����f���vb<r���뼽xJ�G��Hi��t��}�����r�e��o\����N7ɓ�e]���S1�[kS��JA�MJ��n���}�1��c����kxS���v�8�v�|1��r��ͺ���e� %��I�#@�[��a�ۃO幗4�/w\�%�����f���c�}]�^�0ڗ��p����\���h>rL���7�|	Sn�=�mR
��Zp�z��gv��C���P(�1u�r.,�f� �e���Nl�NץZxT��U����c^|{�?M�Cy5*}~�>���v�([a�8��̭��rFi�N�s���Ǳ�"�q&Sp"Ufh~yR��{�^��ӝ������ӤK������#��g[��6�R��c���ϴ�e��:[4�z��|-���v��x�Dw3B\�3�x]�w~��n�JT�ݪ�:�˚$e��q�jZ�ֲ�5�3X.TZ�ݙJ�k��I$m�Q�ےIq�h%��J���uMڪ���m�ꠥ����)�S�P6ʉ\�g]p�UUUUAd�R�UUUP�I�yL���.�3��$�Jbk���Ʈuxa�*�g�zvx��T��A�?^��W�<
��`�!�b�e5 a�d�Q�{ۙ���,�����}3t��X�r���d�P6
4M9������%�[l7<���Zjz�i�6iz�Q)��Uk�ʾ=��)�1,���=�ޢP�1�	ra#��94�N���qk��vh��	n4�8������t��[���y�E��<���,��t�N����{�S��q�{��x^��o�持�@��!U���F�V�H����V��Edl��e�w�;������ގ3l��6%
�#�o5Y=����ޣ�4���WB�xN;�3�-���m�-��[V�}�z�e:�y����ۥ%Ȓ眙�z�F�k�-���{�#�<����o(�A������D��tX<���B�B4�o=X�W��´��c�Voi�k-���h�[�J�,Z^-cqU��g�q�����
	2���a��8��&��9��d���:9���w���N�uz�Ŝb��E�l�[[lyǴQ�ջC��Y��f��6!p�Ԇ��;/k�]]Q��b8!��G�����'lnܦ�`F�x:1�O����q�Z�|+����F3G�\��9Ehzv�G��E8zI�	°���wPoVjݻF`�D���8��A��7����� :A�u`�gzHO�JJ���~�G�FP�e�e�G9�u�Bf.�(�����P|�i��h&{k��̈�j.�6D_'�k5۩�%ʋ9vfSʨ�sq�˺�/)^q�����sG���\q�0h��{>��%k$B�a)ܦY�jIi�p�R����RB����b;��۾�2����;]�(ǔ�O8�,��Pu"�乤���F�D�N��dn=�>�H��n0��RiAl�#���^�D<��بǌ�߽(�M�riDYK{��r�A�v��T!�G��N��*��zL��a��*�����M�T���GcHe�Ļ޾�����ӽ�U����)�BOV��a�Մ�x粋r�����z�������]�ad��O��lK��HF�O:(��܇_JTZ���ZG\�]W�i��5�B(�:ym�ύ�r�t�.��U�T��s0�bJ�g0�����)�Rn��VǏ���TD>�so�b1!x��4D�ѩ*���Ӎ������d@�A�؈@\L��V�Gp7<{;���ѱ��n�)wh^�a�-vSYҵ�k-qӞ���y����v��nC��U����Qc�i4�r*�<T^�#Q�(��}�`��Xu\�T�G��e7v��R�w]M=�{�f�Z�[����������z��)��Ԑ,b0�9$�$c	C̬�.V	Q8r��YMDN��3����}��Mn�9nPt�egy�7�D�b�cΟ��Z����[Bv�ɛ4:�8�+ג�je�o��p��j�E�H�D��Ҙ���ܰ΢���H��N#ޜ�ϪT�p�%F����^�]""̐aY�ف��(�2u�ރj˯zCKŜ,��KN{w|�p�����fL���4�"��O9�o'�K�~E�Od�z�׳kg��0C%�Lz���Pm�yzy�*�*����=�����Tk O��d��M4�?(I�N��X�ˤq�2����Ա��c���{�kѰE�SL��d��^x�`bF����{I���c�j�H�Mp����0�@�=��z��[$OI������U{�A����^�x`%���Z��ʆ�^��1kn�h)I(ܡH�m�dq��Hf�AY�s���x��T��}�2�Oqj0{���wd3��!�����z��i��G夽���ϵeev]$z(�z���!�v�����v���-�\�Y�����]"{,�Ar{r{��R�
9sP<���(,�]�ɲb=fKmo���3U^M�������N��ߟ}�>��=ީ�'�i�[�<�^�h�o�H�����E���@`���m�q�.@�U�F��5��e�������G#�E�'w��\V�� �"���麮ڄ�5�i�����_�o4�HҰ��kF��f��d!/I�ƕb9Ɔ�W���1^N��]�:G�B���gL������D���:_Q�<ʼA]�g>"ʊ�z>�fw�绦���Ar����Wղ��YVs,�gT약Y��fm�~��T�UUU׃�ֺ-i�k��SU]U\JVQ�V��ح�U[,Z�糪����� *3U*�UUT�UDդ�Tک�%���)�[����݆�?t�u4�Y��0�ɺ��diz�m�l�G�u`�,j��+��e�Zz8J�m�M�UUK�)8T�3\ED4���n�)n��S���D׶�h�ԽIƬ/><s'���:��t��U�5�۔w�3��[q�!yJC�^�.�u�>lW�mo����P��MUV�7���(�
Շ&�;=i����!����<X>�;&�e�V��Y�#3Ƹsu�$%���'ȴ��	$j4��8�� c���ϟ����u�����N,:3����F���pm�9t�G�t�5��a^����޽�]j���M�(H��bE�u'wڏ��[�qS�|l�k�N�ll��S�2�������A���Pf���fH>�<E^��K-��1�fI$�$�$82%������}�X}��jΡ��쀬B���爌��؎��H��,miI��dx��8�ʹ�ъ���pb��zۜ�X�լ�
;*s�\ɻ*�����Y"X��n�6斓غ�GMZ5><�����&>�3J�";n+K��x���W	�=N�E�8�\v�M�F^�۱ǯ*�ݷF�걺�v7�1nQ�s������&:�,���gdۙ�>;;�74�q�V�Cǲ����Q�9�ڸ�to��w�<(޵��Z�M�˸n��Z�_
�C�_R)(�:n<��G㨃4�x�!f�/�JH��^�ve��>O2��R4�m�j��բluuҪO)h�`��p����d񮳈��U�)+V�v�r�>�NU^���oM+	-ff[ܺ(�h��h��K�gӾ^\G�.�e
�$n���]�l�L#��Q���������y+�l(���x�h�����c��X�v��os�Ă�%�V�-T�J�i��X�څ��c���m����,V��b^�6|E����i�:v���t��>�(R��w��)�F�i|�=�r�j�>i��	
5�"cQ�L��Fr�5":���V[�L�!��t�Q��ܐ�K�Ο^Ŷ����^y��L���-�@��]�t�hô����.7c�6ބ��^zK��4��	|��"���Z�?g�ߙ���q��s�ڻ�0Ρ��s^�}�D���FX�B�'��F�+ʢ�"ף���e0}���z_cU|�o�GR�A�����Z�nF��ϯu�UUx�,*&��5�̧d�a���7AG	���4�w�˝�rBج'!z�2WC��Y�#�$�T9}d��;a�}�+7�n�4QV��x�J�˘
N�ۅ�&����̂b��ټM�����ݡ��փ�pSz�fc�&^���>9��B��l�b���������L8��N�D�:n��ZWJ십��o:��$��s�۪�Gׇ9d�ܳ:��Nn�G��BWD1i�
�s���<��ܽ9�!�l��˺���Ϋ�8��cb����T%Xf1��&�C��;��N���{C�f�.�q8�|+�3����Ǟ����ܕ7%�-[�iR2��Tlt�u|y��j�n���S�����{7"���Yxin�Wv�j�zcc��'Ug3�ǝz���e	��v�慂��N��uz��]*�Q#=�����q����/6�J�(�&F�iE��1��q(u�ꭰ�i"&U���)P4\�ђv�۵�f짍`�lS�G4�W]*�l\u��/W�h�X�{I��Y���꧍�E��x�1S���F�����s��JΔ#�ͣŧ��=e6l�S���;.`��U��.��-�ss��n���#���7K�������Aȡfwۓ�+�6��].ά�v�f��얍ܷkX޻�N;�ݻܷWl(���`ϥ��y s�g/1�헎�=>��k[�6�ݚ��*���ہ��m��#��<̇cv�@=�j�L�]s��l�kv�{s��6$�Y�h��!��Q�Y��z�pٻJf��vM���9��X1;��to.f��G�6�N%��%G�mˣ�Cny;v��L��Q�.r�瓗H�krp=kv�Bx]�s�K�w,��h�Ԙ�����7
�H/C���%�8س�K�7��6�i�qq	�IA���Lm�;<�*�=�ap��x�������ɋE�gs�33ŷ��ù��;q�;���3�t��zյ�j4���kr���>1��뗃=/:$������Xwd�W�fك�풽5{q��.��ds[�2N�w�.ݻVg�Eʓ�ە�&�ۣ�]q���()һ�t�kxuf{6�o'*7�xs�k�i8XP��a�G���<���{4�5�wzZ7�D��(��̾���:y8@�8�H���s����-6�a ��F����ʘuv�����<���FB;SĽMċ��8U%`��0�C�=�N>�����5�Kq�N�I��o]��kq����]r2��tW>"\��k������C�紨�|��+�w�r׉��tuXPO>^�LͬDIV3�����ԉ"Biٷj .��`N����|�J=�H��E�{�L(��.$�wT�����%��^U�(A�%uM����$R��ԇٓ}v���#�4���}S�\v}w6Y�j����)�{����͎�ӰH��zE=�	���	�@�w&s�7R��!�=���Z���Fi�4�zO]f3���g�U�^�L�IR\��r�m�O����-��돏j=w���ɤ����0�q��y��ی�n���m�p�^\XK��k�Q�dy�&�,��[Fdx�/:�xJ�[/����e�u�ݫ[���BU���};��ljV���+����7F�(�~7�77�{�B�e�ā\��^B�Je^:H����2��;,����.^�,�[����^�����dFB�>��|hz�8o����d�&/+AB*�x�f�=��[�g���]Wb6���e�5h�a�w���]L�Ӌ��"N-��^��q�A�o�9��L?]��2�xr�(��yY�ڝ�����iX�	W�d���`�NA��d�&�tT�$�9Ǚm�7����z�0�5%��"`�J�\̞�ٞ�P��,�pƘN����������K�<x�-:�=X�Wb9hJ�y�c����r<i�lvy�;�.f�4���w�'tKhCw�A�>9O<׬o�E
[�л��#�qf�E��r�m�
d�dds7��JRy��e���A��B���gG:����粅�>��p�����d6ߍc"�[^�v�A(���$�r��Ы�>z!�U�]��Q~�ƒ���]�O��>����s<ь548����R�YW��F�z�x��[�����;�O6���Z����t2tq��j�ɻ[c���31P*���Y^��,�j��ꪛUWF�u*��kSr��wm�%Z۝���������
@I���������<4���'3m4�M���='h�~���}^�=ɜ�XM��A@�!�z�q'���GW�"��u����x�_EW"r�k����ix��L��	�����yq9��]TΗ���g3�$�J�T������t�3�.�4���wfj�[eA���/=���� ��r��^�`gJ�����N�Nb�95&~�����ŏt�e���-���~���>���1�6FN5ՙ��ʅx���W����4Lb b:#�mϱ���n.�b�Cj�\}�q��>�&��+�뻵%Q�g�8N*�zD���:҃�R�������ˬ����|ܑ�d�HkI�����fԖ8��@�K�j�æ��(Ek�����{����o^�U�8772�"d�7j��:�_z��<���P����l�[�J���0gz��հ4�J$�JFآd����V��[�U��mk_3K����($�BpB�H���aq��-XN��K�h����*}�؆�Ųw�,�Ln7�,-|g���N�����ΟfpP���2ܘ�}�J�Y؂Žj����o3^�wW�YhgɄJA��-��A�فMq\n��g����\�\��E����{v��������Rr���6���ѮeY�;�/σ�c�q5�Z��F���9u%�[cpl%��u���/g�awKw%�ֵ�`n�-�8��x1��1\s��ާpd3�{lz��?���3-�#�*��|��ܧ���'�;��}�~���+Չa�v�S�8x'pC��}*̢ ��f���]/I���xwr��-�9G-z��¬���0��)Wژ�$NC�qBb�ʛ�M��5�dVuz<���Ӆ�1�P0�6�AD����?��6�3���&��GQ	��ԥ��"��T�x�f
]�z�sb}�}�-4���TC�+x̒0�_%?{҄^\�AR�(w�'��B��ި�/�����^��s����&Z.l��+��������g}�&��y��vZ��!����TD��	��b�3�*g�O���DwM��3�h�ƠC}%S����!n���E��t��WԚ
_#EkC��Ԧ'��/]�z�t�h#I���A�9�n,#l�}�EJ����I��H5���2.�C��B�&�t�Wmr40����ޚ�u�\s�Jv=}�����U�`����xd�X[J�O;J��Ř\��������9;�#�-H�H"{������0�m�l�ϟ��?{i��¹w6��b�r�#k�$���S$�(R���U��Nؗo��/9�l�����&��Ol�U9˖��w{A\T)ȴ�㌞���ͩj�)4���#K�Vʤ���{T0�u՘�H-Q�8#�ټn��B�!R�U��� �<$q�S�~���w�m��8۟�-@��T�������Oݎ�N�~8W,�6��0gw��8pr��E��׭��MTQ뼱̵�N���G��U�dH�m�b��c�x0���QRk�hg����8t􈡼��H��*��hU���^�گ��0,b�nZ:�Ma*���A�Sh��ㄑ��n��,~�Κ��U8���>�9��z�{�U2Rdiio7+�o�m���r��,���xSAz�ܨ�ӊ��/;ㄙ��"�l�d0�4�J(���Of���?z�����R}/���w![���á�Z`��1FdyG�8�8TɽK�?U�Yb�֮��u�]'�/�y*���I��3n�!#pf��#��b���	Э��1
�<GyWeo���H]��M��4k�1��Ѣ
��R��������t���0s+`��$���|F�o�@��
n��P�B��`�2����8笪�q��Bԇ_�8U����w�q���,��tW$���ȇ�`%�K���'B�w���;uF��*ȓx��q��{2��pU;,��dT�?F9B���쁩:���΢rF�NƠk�b�u�^�!�#�S����O�`���eI��1
T��d/���V{��{�[�%�E-4<̮�A�r�[2��|E�5�d�#ң��X
l#��Y������F{�z��F�'M���wv�H�N4$F�y����[B���	9XK���zM���,�yUDy�ǁd>��K���/>+��Bz:%�x�ԁ�w�b�&�D��@��	/���Ҷ�8�uC�ؗ;2�:E�8Q�XVu�C�n8�n��� �9%��������;�]N����ڃA#]��i�WwH����Mm���J.eV��77�H��#m��q��f*L�tU 5�������L�H�a�ʳ�ŕ�t��|�UUUUTJ(��������$&�vV֠��gJ֩$)4R��a�)X����u��o����s�=���RE�j�tƇl�)T�*�ğy4$e�,���E���ѭ�2�K�v��^��=
��x�i�=�ZH��W��Cɪ�d#�C�yˎ��n ���r�,�Q��%F�L'A(:6�I��hS�C�;ϫ�O3���n�N�YpI��-5f�}��:*-���0A6��\C�$�s-to8�x��w�����Q;��V�㞈�[��I�3rB���s���}(!�yW*#=�i-l�C���~	a����j�A穈Ox{x�!AA�����w7l�����M<g�ւ��]z�[%��+!�_q�{.����L�����8)`h��d �4i/�I�(ߗ�*��=�����r]�fm��\�mmT�8 mv�VŦ��C.#�0^ɲ ΡT���t���}~G��͓7LLIZ���O�<��IM'2Sn�I[	��F_�խv_����>�`����?Rz�Z�Q���X��h�n�]�k#km�n*��_~~~}������g�͘K�LP���ݚǔ���aP�Hcͫl���ݼ@v���<�����Y]Ǉٰ�n�Fʜ�=�*�u:�l��ծ�y8�3�2nt�r�2�b��͸�\�v�]��0v8�rs>w�4���ܮ���}��#�ߪ���d;�'ڹ�\��>i:��Jg�ãe����Y��`b�֑�C�xҺ����m��!��z�o8�Z��a{�N�i�
>#���r���p"���V�jx{��&"i��N��<�e�7ʸ�~;��j9�sYL�kn9&Ÿ���$��{}�˫:�d~m'$����M�6D�4l�
\5�_WLN�m�"
g�����������D���T���g�o�IŰ�|FL�7���zY(��9��X�*�����_>�y�q�}����U�7Z���z9lܿ�~-����)mQut�$
�p�[!?z���X����=*5�#i{�z�D 'f�z[j�7ލ�P*N�U�b��f�G�Ғ�4�^���ަ��Ӿ�7���2z�:����Bra�ϡ�P�=�O���T�Ϙ.(��o�z��hyى��i��o2G��UUE�S��%�):N'�����o�l�0����/Ë�ܛ�(S�����:�صQ�c�w���ϩ��=��"|/�NMS}��
����Dt.�a��y��QN�C����V_&����O�a�cd.'�ċո�$X�z�;V��.�?�.8=Ӳ��Ơ|������VtK����m�)�5�mvT\���
m��!���LW���f�u����q�B��h�Ж��S���C�X�M_���`��C��zy���n)�R���y���*���  ��Wg0�[4��R�[�����co�̠{����Xl�w��Ӥ�^�u>B��]gA�ƏI��q��B���<Pܓ\v�H�Ð�j�ńn�xR�l��mu��
!<���N?~'��mAb��7��]�w��.�sEۋЋ���ٱ�B9"�f{���OW���5'�H��T~c0P�/ޤ&�i�bR�1��������R��fǄqUx�:�J*�I�oL��p�Z.0ZN�)D�I�Irh��9-1���+��iP�����U����Wˈ��
,�Q
6oZ�����S�Z��+��_a�-�f�݅�YR�κ�}"�Iw�T]���1���Og��Y���q'o���x��"�z,0q����j�z��V�O��}�:'��2��t��P1�J�@`Ȇ���/&[#1�}��7����}�\Y���e(K�E�7�bk�%޷�͑��Si��dz�9�E����>N��+�/s�[ܔ�u�|K�9#����h�Wq�Ѥi��5�ȍH�'�ߩ�zZ�����6<t/h*T*j%e�\m�,+{�9Y��̅�F���n��ِhd�F*�f:r�S�ة�Ejީ�.(�=��%<�D�I��+�-'�`�ͮif��F*�*�m�긍ିV��S���gn!��=�8Н@�Ť!O�-��/�뒅�(�^�ܝ�k��<F)t�6�r��w��>����/r���H
2F���i��4�R���7�lbһ��Ehc��^<O�
�y<��{$OO�hM�M6Um6I����%v�%0�Q����v�����y�r�@}ʪ��}ON�\��{��*�"I�ջ7���_,QU�"�dA5b�\1R�� ᐒ>�D��%M�4���5�Fd�R�릭yj㶛{�إ)�.y����������ӗ?�����<������~;�Ӌ�H����zx����z�2U 3?Z��{�����^��mϺz��@~?~r�wtl{���{��K���������yP�̈*�C"	�R`�a$��I�R���:w�YT���O������=}|=˓��xc���U 4ftk��/g���Ô��v���o��p�i�M{�Rw<���_�W/�
�U 6��g�UUZ9����P�K���aZ�_���?���{�i�Ɔ�YT������U <'��o��m��9�qc��}�զ���<D�ӯ�E�Y��*�=�^.ޟ}wc�gg�ٷ�ө�{^^���ϷY��������*�X��WV:�unq�v����Ǜ���� 7��p�z��庪�����i<����1AY&SYr���c_�pY��=�ݐ?���a-�{�     �J�    |              9  @                7=�  z
    ��UmU��ԓ 5U�QU�UU�UQ�B� CUb�Tɨ 2  	  ���@; �ͩU�U+&�` mB��Ҍ�VmP� ��P   (uUf�T��U��@  ��EX��D�j� &�fjVZ��e+6�, U� $��@�@�  :     0"�!� t:#J���@A�uVmPd22@A��Va��Mh V@	@�        ��]��2� $� j�h��UF@	 � :�閨�C,���� 24mL�)�h` �k&�caFl� �  t    (tت����H:�D ��L�$0  �CC ɠ` @hV@5�X  �k62�'�     �$B4 ��Q1OMG��z�����&iR�H�      9�&4��#   ��~�UR��*       "��UJj4���4  1FjM&iRJ z�S  @ 9�����޼<�?���9t�˧y��~]�d����V���I�
�(N�BR��Tʪ�[E��W��`��x�b3!�[�QK5���IKYR̨���u��y�i߻f����k\�(��ە�~��mw���7w������%���;�����{�;��E&�$R)�FH����d�)) S ����H(���Eb��AT"��JB��YH��V)
a)"đ`
(��@ZJT��0U�R"��TS�)�ȰR(��5B��
�������� �)"���BdUAX
�D�,QE�EQ�U�Ad( ��D`�X�%%*1`��!)B���T�+`RAH,ȠE`�AA���#�"�E�����2A�	L��*�F�%0PE��d)ED��dX� ��X@U���"�dX��"+QDQ�V�B���@Td�H,F�Ҡ��A`ƅjBR��RE�Q@A��B��E��T1dXU�0`�	E# #U(X�M"�"��"�F��
�E�� �VP��2E� (�R
��Q2I`�,��"� (�
PH�EUZ!�EV* �(�EH!HIL�("ȲQ ����Q�Q#PYQX,�X�Ņ0�db��
4�E���,��ADI	R�a%!%%1T�ET$RF�"��1�"�H��Y!D�"�Tc��ADE �����Db �*"��cFA`���VAJJ@��b�Dd�B(*("+�!�BER�*���S	$��ILR�H� ���T����k)��̢k�C2$U���,0�b�*+�A�H��TH� @TF��)"���U	CdbDVEj�"1Ad��PTH,HP�Ԋ�!HТ��,�QX"RP,DX*+M"��PŒH�0�F�jS#U�dX(��$) RJ֖�MR�T�kBZ��S$b
F(ăL��M�c@R(D@��)$%"�H�HR��2@b
��!����"��,R	FJ*QMU1D�""DDR�%"�����1b1���¨�5Y
RQKcY�eIk	3��LUS)�)���
��
U�P�$$�5 ��J`���k
�a,P��L��cX� DI"�U$`BJbkEE�U32�jkXř�(@X� B�((%2�V��@ֵfSZ�V��0ı�,�b$$Q�Y"�!R�"%"�"���X��)))��""�B�B��*!d� R%*���� 4QUDFAb�I�e�(dj����
�Xʂ"UM1h��P����
J����*H*0A�*�P)
`1��R!B�)B
I��JH���@h���X��L���B�,�a�JQdQ�#% JB���)����(TdUPb�`(I�	#R
4"ʩEJ��TU*�0�)�LX1�`��(F P(�F �P,�I"�@RS)A�XIH�J��U"���"�dX����Š����Ti���E!H�����J�j��R(�R�@QH�QeT
T�P
RH�B)�PT0�(�"HERI���������PRR@XRH�X�XDI)
`��ADH(��X�)���@��%FDQ�E�(�"�L��c��� �h�C�R�������"
JdD���Db,��	CJň��#�U�,��~�ܟ���h&�
4h�K� � �����������eh��٣�g���ݰB���R��
��
�� �*�@  � UT�� �l�� *�m�� ���j슫dEP dUrҠ���
�Un��P�__@
� d    ���q�R� ��U  )�U  �P  ��T�*��@Sb�T�>�m��      T *����*�6�m�B�W�e�ϥJ����l��w  P
�P
� @e�Un���M�U   �Ped�*�`*����@�@gun�WɱJ��� �  +(��l� ���cq
�V��׬� �m
�VQT    �V֘*�B�@�@�[E5Su�P�  ?�W�蹀��N킨  �U  @P
�6�wWT�[jB���UUݶή�Tx�h�`     *�`w
��  �k)U�ؠ  P
�6�@�@ *�� ����   � *���R��@  @�   � @ U�UX��ϼ����m�����   P
�  
�    **�P�*��@
�eU�.�@ ���R���2�-�YJ�� � �T� 
�  �v�m�  n�   U �mܪ��wT l*�P]�]��w�h�������g-     T          *����͐
̠  �@    8M�� 
�  *���� ~��   l�      ��� P � ��@              
�    *�P 6�     @ @� �       m��� *� �}        *�m�        �         T ����uZ�ڞVPU
�T�5B��.���6�       � 
��l�m��P�S�@ P F�U  ��m��l�����x^a�ʶ.ݻ��b���r��wv�nPng;s��[gvͨ  s�WL{vmݖɰؕ+��� UTPd
���p  � �*�( �   ���* Ee�pP;��H�ڥ]�R��T*�T �mP��ꭓ��˸e۽��.j�y�U}��J���[  
� w�m�z���   V֍]��J��+(�[L�*��_~��h�
ʽU]i�o^�5UQT R� �U�Wڕ@� ��UU  
l�(� @ B�  �  -��C���e���*�P ۻp�U�*�]Ͷ��X�J��U�� x���{����m*��� @ 6�<�ۻ�7��|�iz�귘Y�0�۶�V����R ��,8{�or�tw^ʭ�ov����w7�Σy���D⫻l�w^�]u����*Y�^;������rv�f�c�.���{m��V�lS�j6ʬb� �^u�i���W�v�h���v�[��s����2��ˮ{�uv����,ݭ{;5�j��.x�u��}�����;���2��[[Ee۹ܪ��.\Ͷ��[e����C���7��yom����v��E��m��� �J�b����p  �۴�ض[z�[̸��QYM�U�W�lP
�q���[�]�\�*��5�*�Qz�v�Z�ש�u /k�ݽ�����ws��!M��{���S޺Vmm����l�R��YB�/l|lq�,���$���,�I�ʻ���[��Wn������u����M����Y�9�S��oZ�`��M��M�u�k]�o��uU⯍ݓ��ڭ�   ],Sx���ۡe^����.)��]�쭪�ff�^���d8J���^� r˷^���]UT�m筅P 6��+s���޽յ3ض:����[wV��w���ح�^�3���T   ��} 6�-� �i[6�z���ۦ�ݣl  T�]V��   �� �} ���  m�*��  w,ʮ�S�k�N�   /m��    �    �  l\�  PW>qT }�   � =��s�w�akv�  U��7���U   ��� �@   ;��l��w����5n�Xm��/l��Z�ծ�6=�Ư��n�{�S�                �          l            
��                       �     
��UZ�m;����    �*�6�  � @            z�            �@         s     �                ���          P    
��>�  
��l)��s����[n����P�wu�Q�uP*T            ?A�             �          �� �       �P �n%��W{�k� 
�    p   ��
��h  @        �}                     x                        �P �](     �   U [    �@   *�                           T                                    ��             �           �         ��E�    
�   
��         j��V�}m�       �U �z��  �   
�R�      )�TU 
�  Y@ w  {�Tu�T� w         �@� {(J� ���J���m����U���v���� �y���U�l@ U�ss��{J�@                 � �P      ��u���eUM�Pl� �*Uz��հ�7�P ��m�ˍ�{`6�         ֕�{���e�e @  *�*��{d��  � *��      � �b���ۮի.�"�H���ݚ��a�� !!?`�Z����'.���7S����������Ͷ�M�(����������������Z>����{����h��-&�m�X� *�
���U �P
�K2[M�j�@ �6�bT*�۷b�;��</U� m�[m���3 
�T 
�Զ���`�Q]�
�   ��� ���P� 
�6�� U' U��@�m���p�   -���U  *�@   EP   Y�� 
�   �YV�\�©T���Ʈ���kv�n����s�=�� 6�T[!Tp��� M����en#u��� �l+( 
���.�������*�{q��,ݶ��ۋ6ٵukr��,60>z�U�^�{ �w��Kz<��`ؖ���WMKme
�v����p�le��ZN��M�lλ����']�N����K\���/h�r�du��G ���g�"`�{7K�ٵ�*Uݶ����-t�PU>U{��@
�m���6(|m6K����@�����eM�    P P    �R����� �        �  P ��uul�@ T    
� �VP �d ��   �    ;�pPU@     �      
� �  � �� ;� � +2�l � U�  ��m�GqOowe:�K   T ��lP�P�)� 7\�h
��P  �l�߯~~����=��z�~��Y��պ�UQܩ̻#l�lS:�����/l�� wFتQl������v�+B��ex�7�{i����ޛ�6g�)�+���ގ��^�ժ���ot�Owc��;�@�*��R����eV�;��*�m�*�U[j�&�o9��6����c;n���j���^��o.f8�i���iy��Nl�¯[�z[��s��}��E?���M�1����O/��~otw�},���'u�&-�M�٬�kS���
ǥV��b���BC�	X�|IS�4�o�M�j�0�_!�vilU�G�wY��^�W�xD�t"�-6� ��&��m����f��L�/��vk�䄥I��-��C)����w�_Y�ӗ��>m3_v�뿟���ͨ�ڛ����ɻ[ڭ�{��Y[� �mT ����k�p��ћnO��l��ܭw���]޵4��tk��׬�w���h�vb&���[I|j��
ў
�z�Ͻ~m�����Q���y��nCX>��Ě�L�mJA���`vjf�\��;Mm�h�8o]���~Ms�������r�2Y�W�m��A����n�������1��מ@�cE1��H�0�h��dh�kG�ob�)�<4)ITh�Kv�F��V�y��C����@�n��ݼV޷+{�`]��˻l�WZ�ڧ�����|����m뿨����=KN鯞���z��
�'l�!��d���h�Qn���[�jq���ӹZĶu�k���h��7J�����)�[.��N�U��o޼o*����{�}h��Am�j�B�1��kx�2�{�э�v���sOi�5���9zy4敶�Z/Z���z�����u��s�OS��58�u��\u�l���Ϋ-v���V�k�]��wn���7v�� 
���I��MRM�4Ҩ��X���oߵ��=v�f����-���
1��ID�i��H6��cExA<k'[{��^�>e��y�z�/���&�{U���]]�鶺�:Ν����x�����:�3�k=N������u�5���m�]n
c����,h����c0}����h�jخ
cF
��M��n�A��
[��h�7ƠB�1�s�^1�U,Sױ$��+tT;��&�w�U7��w+PTm��q����[ckut�5�sOSi�5���9�wW������9������ZQ �e��l�+G��*
c�Ntco_�����x���v����浦�A��4��Lh��e�P}��/C+���{\�pW��h�yV��]Z��]��޻K���������q�9���6��;���:�k3zִ�-)$ZU����aCZ ��'X�B�;���X����
cp�m$�i!Tp*�M�ݵ��ժ(����lڶ�� ��P  �*m�������e빵�l�f�{Z��sͩ��]K�6n��׺���n�{�w0Wwu���ͭ�\�m���R�B�Wt 
� `U*�6� wmV�
������{��
��� ��*�&���k����W��s{��`V�Ed�w;��Zj�Rh�(��@�A�2q�)�)�)�h��Ɗ��|j5�i��M66�e���nE�b�Ֆ�c�e��S,j�M@���:�g[L��OS��51���}��[ı���;���M���4ZM���;��-滗O]�Y�빭�[׏w���A��
[��h�
��i��TL�ˣ'[{��^�>e��y�z�/���
�X���X>ɯ�d��D��Iu9G�N�����;�5�mS� *V�b�{����li+W��6���yGY��9�����n�� �v�*��!&R�S	�޵ej��z���~l������oO]�X��71�����*k�!m��m�J7���[<�+C�1\��m�P1��<{O�0U�Y� [��i����u��_��So]�o4u�m3�k4V���+G�Ix�L�M���&���>u�2�����s��\��o��=v֏����4`z�m�j�	Bm(y�rm{��s�lֵ�*mR�w�j��m{�4�-���h�[��cExVO*���ǵ�Wx|�qTh�Y��6�+��j��������q�>��{�|��f�V��1S%(�Z&�+�e7L���s�_��w��&���֌m��W{�!���մ4X�l���%��I::�%�x����i��*�����i�
�ǔ����>b�ؒL0U&�(�[э�v���sOo��p�}��SoG�K��}����Z�A��I6�4KL=z��m����{w���@����U�{v|�F��x��q��\�ӯ����ol��Lƅ@��
ž�0S�$�A���D7u��N�U��o޼suxQ���w�豢� �PAZ�I7�Ke$�a�w�O�n=�h�޻K���Oo��Y�}f�W��5�!�M��)*��i��X��u�s,�I����淉��-�<+P��l�[%&l]1������h�wa�)�6y[5h�[��cExM~h���H�)��Wy���Uۻ�י�N�T���U�ݛmc�b�1��+��)�6��b�=�H`�C�`���Se0�6�T�n�W��&o4u:�g0�:z�o\�1�u���q\b�&�-D���i�I&�@Ƌ�|1���մ4X���71���j��(�!y[i�A�oC+� �{\�pW�1܋ZŴ|�i��oB���w]��7z��=~L�h�:�G��h�d@�h�⍠M�Km�VP7\ֺ�-��Y�����;����k� �� ������c�w���z�x� ��g�V�m����<��w�s�8[��WZ��K{h���3l������Um��m��UU n�Vت�� 6� w)VڥA�m���}��l�[[l�M�x �tgwn�������+"�)e <���M�m�`6�H2��
�����6*4X�[��c1�hh�(���$~E�ʤ�m��qm��um�*M~�<�ׇ�A�@Ƌ#��"�W�M���ޚ�_S�]�o4u�m5��p!��(�QE&�m��!Z<��ol����.�v��9��ܷ�o��=+G��I+Al HM3pS0l��ь��{�}m�|����v��>�w���6�m(�[�𛲮5t�Y�og\�� *�N�ڷu{m]�w]��:޻K����������8f�W����ˊ�}�H���`��i�E�jآ�]���ol�����c����w��K{�%%`�� S#E���9%\ƌgۭλMw�W�ާ�;Lq:�wz�6ۦ�l�[e��+�� ۊ�cE�y}.i�m���8�������y�5���M��e���nTZ֭�-��qG�[[-G�ӳ�$�m��D��m��Ȳri^�����8[T�@*���u��l󶲎������r����IW1���j��E�[��h�V~R�l�K%��@�hc5�W�Zgw�co]���\������q�ڀ
i �I:�ڽ�e�z�˕��I BC�=9�o�"JBy��������a-	��6ɿ�}����US�
`�Y8�Hez��5U�۪�ִ٫�kd�0�
d�RC�D��h`�Y-���Q:�L5̼7
d�RCuD�
`�Y/]��ϒ� ��)�0�N���/�V�)�
`�Y1�����������[iz�޷���6�HeQ8�L=_:�Ɍ����)��l)���w[�$=TAN S�ɶRC՟{[ ��)��S&2�US}��,Ke$;TAO�)��wZ�,�k%J��qܜ��vv�gom�{���B���ڭW�ZV��UWz�p�Le$>��%E�_ڹ��j�)�
a�)��RA��ՐS)��d�RCuD����aL�e$2��� S�{f�c)!uD�
a���{��UvkZ/Www�Wz��!�
|�I�����z�d�0��2c)!ʢ
w6�H,��Hv���@���7
d�RC�
c]fz�	�%����	W���W��U]��a<���|��g��:���O��3IUS)�ҹ��u�<�q�&�IV}�l��@�aL��H}TAN续sZ����Wwuz6���NUAN SS'I� �P) ��/�o�2|�Hz��Y1����\��s��0�aL�e$=TAO�)��^����Ej�ꩺ��&2�TN!���^�Cl	��g���n��'�N�n�M<��]�a:�m	��u����n�w�j����jw���m�:�W�th w�V�6�ۭ�m]ֲj��Z��&z�)�
a�)����}���$Le$>� ��z���ɶRC*�)�
a��P�O2�� � S����w_y�8�I�l����5��Z�n��Zn���
y
ێ�}TAN��7R�� �P)�F��RC�wD�������m!�D�
a�)��S����c	�&k��KVSw�hӫ�p�B[	�M����l&0�Bc	�%�7��&!6��0�N��}���l)�IU��ѫ)!ڢ
u�<���tӢ�V���VnɌ���D�.�=[���)�
a�)�������V�)�
H,��H}TAK��Xa�)�l��US�����L�e'���U�����ȒHae$�,����C�D� ��{G��l)�I��)��@ZAd�RC�D�0�8�Hv���@���oW��L@�8�Hn���޵�]� ��dv⺊Vf[nݭ�T7Y�����ܭ�.`  e\����uk�ͨ ��K���]����7v�++l�����w�mf���^�ݲkf���6��Ul�� �  ��wT � ;���� *�����_Aml< ~�����U[j ��w{�W[u-˶��� ���we���m�4����y;�<����F�)��ϿF����S&�I� ���w�ٸ,��H]Q1�q�2o3�ks䇪�)�0X,�e$/��삞@�aL��Hr���o��UmӪ�֮��6�&�I� ��÷��S'�I��)��`�^�=[�$=TAM�SaL�e$=���AO S�Ɍ�������(��i6c�[�s�^e�wyf6��s]54�8�~|v���@�����UZ�j��֪�V���C*�)�
a�)����ｫ � S�Ɍ���)���6�<6�HeQ>@�����d�RB�)�Ì��}�oɶ|�ٯ�U�kTi��WEӫ�d�0�
d�RC�D�JL&�I�S�����p�Le$>� � S��z��n|��Q6�L1�2u���}��<�L&2�UR��J���\�T;���Sz�;{]��ywpl�օP �(4&�#h��쥧ӻ�c��眲m��ʢ
q�z�u�IUS)��S'3~�>Hz���@��l���>��AO S��Le$>� �ol%��� �P)��*�.�SWwsp�Le$7TAL@��_ڹ��UO~T�M S0�N2��?5d�0X,�e$7TAO���6�<6�HeQ>@����u���Q:�L>aL�����ݚ�Z��M֯[�$2��� S���RB��oN�)�
a�Ɍ��*�)ܔ�,M2�� �P)�ח��L��H}TAL@���y�nןw޿�����ۤ��R��[rX�
�ǔ����>b��4X�� 0�] �&C
�i�m���8���}N�v����u�ŗ*�cEX��I�KH6�f�m$�x>,�����6 �*�w*<�n�u��H=v�:�u�}��[�m�>�3��y�>�K�e����c��c�&�MM�b�G���Mw�W��|�i�'~��o�i͸�TB �M �U��b�6��`�C?b���>u��QSR���͢�eެ�'R�j��i>v��o��|Ϟ��[��X��G�<+��ؙ�I$I	�����oަ]k
:�;Mr�5��Z�1�ȉ�m��I$�)6ۤ��>.�r����ͪw
�l榌�Zםر��������n���驧�ǂq>g�k���^�i��L��%$�e7Z>��{OE`�5�jq���|��}Kgκw/I��i���$�a��I6��#EX��LV����%�LoXh�8�5�����N9����CMM$%�ȧ����hb��M�H`�e~��PV���P�(�̖�uI5~O�������һ}/�ķZ�4�;^e��LW��*$�!&Q4�m��:c�0�=Q���m�m�*�m����͞vQPtSF�!V+��<+��,�LV
�v���[-6kE`�[�a1I7M4���N8����g���|�q��G[qج[J��X1� 4�,��m��b�V�V�
�E�����8��0U��V+�G��*i��	�z*�x��n��~N�QO�o�����j�ܭ�Lh��A���h�S�PV�
ݻ��xh�X�hc��+��)�6�;�{~~~~�VUP<**�]��m��m�G���ޭݥR�   n�n:�]]��u}�]�x�@�ۉ���7;�/:��hgWw;�vګ]�[]�,�`��wX�m��k���`�*�T�P��  � 6��@� �T��UE���w6���*������[Y�'[%G=�>rY���6����P w�Wus�m������|�>�'�u�_S�]�~o,�u��kV1�/S6�%4�!��o�v��N�7n;z���O���tz�:��p�h�-6� S71���5�<+Vڂ�X�^O�
�ǵ�R�m�_�(2�Z��b���feEkwX�qh�C�.x S�IQj�4U��N4�v��o������y�i���';*S��~��~��S����ځ����w�ӻon��j�ڧpU]�mr݊��,�����{����n
cF	<���)m=��1��A<j+Cx��ƋI$�	�pW��A�'�r��ջ����V�u�֒@�1@��L��ކ(��z�V��+�^o+}O����co_��}�k�M�n��칹OR�k5��i�j�ܭ�[׎n��P}��-���E���VB�Km�L�V�3\�pW��A�@Ƌ�i|�
��<0V��u�R�Sd�[Ij	ɷ�ҍa���f��B� 6�λ�>[wSbH���(ˎ�}��8���0U��}���a�.�V>���v"P!��5ej������eJx�w���i�j�ܫ��тYr�A���(���e"�H4����	�P!��1\��m榞6�k�������j�JkWw5�ӌ�/ER����1Gt��1����� �S��3��Y[-e�>�,|ϖ+�����2�I�Bm0p;�&�kV�'�����U*�E^�۹ѽ�0�m�I�5�,R���H`�6��U�r�
�������j�c�AR,�����[{縬ṯr�p�_�$R;E��$�j�y员1X��G�,|ϖ+�d>I�-��@6���5Y��;Ma}͔�>q�Q�Ho�<�
����.RIRM$�ڨ+C�MM?'��'���}N��{�U�g[O�����m����z;f�-�iٷ]�=��3���� ��"Y*�i$�:b�E&�ut��4ՃӜ�I����[��>y��c��ӽJ��+�W��A��HcE���ױ\�mˬg]��}�vi�|�ܣ'S_kI A��m��m7pW��A.*��1X���xW�����D�H��%��d4̽c����էuE2�}�ʄ���c�R�,&RM�"��0U�k���Y��r��i�Y�λMt��i�|�Ay�	$�M�0�~oZֽ���eU 
�f-�
���dT�l�U�Ue*��s  � ��Al���r��U��b���J��
���o+(�WV��f�R���H-���E6�� U ���J�U�� 
�EJ�9�>��շ�l��A��  �U.��;�  LR�.`w*� 
�J�(   � T         8�k�p� ���CmU��a*�tk��f	�@���T*�@-�� �V+�hVP�c�U�R�7  `U � 6�j���qyYm\x��4�R�=�ډ�"g:��7�v�!��Lg�N:^ѻz��-o\�4VcS{n�����56ڥM����T�u**�\��]Gq��o7m�:��W['��7I�rٰ��mwf�Ƽ��^0�����n�P�.�l��A���}��@R��w�;�Ul��U ��w��J�[��'U\�       �     �'����@ �        �    l^����U       6�T[= 
�m� �    w    �6�@       P C�       � � {( ;�  �lP m�� �wAT *WuV�P�gH����    �Om�Jc-Yh v� m�Y@;�u~{翯�����_�T`[� Ums|V��r�@m���wSu�;�P�  UBsm�h��*�}M���T
�ݭ��[Nv�u�ݚov�����+��[�|�O�������v���Um���Um�UB�� U*��� 6� wTj� 7;�*]նmmZ�6���*��v7��8��fE[il�oe]�w˸�%4@�ٯ�+��9R��&�Ŵ�C¼0x`�,�
�)��m 7��*ӹ�6u�m+���?%��;s������c��Q��a��M�5h�s��?'���u��5�fkx�O�o0��,TL� 1")&趋H`�6'S��>��>e���F'[J�MJ~OY�S�H2E���+G�+/AM;��gY�ҹ},��[�s�:�:��w�����+@�<��g�����V��p ;�T�m	d�Hl���m*!��
���������R�<N;�u���5]�}M8<5Z�H�I�E��*������z���}F:N����kx�2�{�э��Y�ډmRT�m��_�A^�!��3_U�c�һ�5gY�i\�������F��I6B-��A��Ѕh�{��G��}���v���9�R��_���=wtu��sZօѭ޵�ޫx�q��w���h�L�D��{\�y"��|�w�~�W�J[m���]�N����t��w@ Sm�VW��t���nb��;��Tr�ji�u�=�gs_j�1�i]Ϛu��+^�k�Q$��Up1!�r����}��[̣�q�y��co_�����Z(�j	�i4�h6�-���;��4����vu�~��g޽���Q�B�U��!���RI3M��a�|���G[z��9}54�:�����'g�������*d"�L��O���e,f�����`�y.+�ׇ���@Əx�ɑ��-�D$X	��Hu�4��{[���ۣܙ˚��M��[uTy7)ķ��z���/�u���o�K������p1!��It[I��`��+C�b���}a��4_�,�ԧ������u�ϭ촽][�U:�V�<(��.�}��=�U�mc�[���vZ&Ca�� SME���(�x�v�ޭѧ:��۔d�=S�V�d��A�Mi�Ȕ�:�n۳2�Z�shfY� �T��g�sr�޺�n� x
�J�nD��D�d�m�Z�촶m�S�n��ke��uo���2�m"�iSR_���qo�u�9�>ݭ����ӷ���)��h&�k�-��E&	=j=���壗"��]2�!"�,P�R�&��5$�;<��ǵ�v�Y�L$�M�AE7�|�\R\�)O(�ך�j�n^�X��F�%��m����I��u���ZܵH^�a�����Wt� U �U �K\ow��
m۳��j�vwZ���X����+[���n緛\����<��c��mf���s�m�ܪ�UT   U@���� �*�P����n�a�nb�[+u��d.�ݷ<*\�vo=��l��@��j�޶�;�{�2��gE�r�����v�Iy/^Oy$���M�%��Ç+3��Z��̀��&$(ϘM$[i��iG+s�5ɷ��G�V��V,��ii4�I �L��N�y���Õ�-��eۭ`ad�d��-4*���m�Ѕ&k}��#��+0ׇۋK�F�5Ye��<U���v��n�޷.���d� ���lǜ��%����`�j�z+0Ն���>��n\�^`��Ѕc4�	��`�uz��R�ni�y��Iz���w��x��m%X>��V���X(�f�A��m2SmV��16y�5c�)e�Ѕ&k}��#��+0ׇ��z�AM��h ٹ��򻎴u�c�t��9F�ﻳ���n\�V>�R ש2ZL�M1Z4��Q��|����Rq����O��V�����������W�l��l��<m�ݘ ��)Q��mU��Ӻ�ޣ<���{��i���6�7���I��G%��*S6����&��W���BZq�ܺ�&=c��Y�q���K�q-5��κN?<̼A�T�m�w����hm�X�*����`�b�F��b�Aoɲ�i*3��YZ���ח��bF�u^FaQ"hSi��Bkk|�5�����^1�kqfm�$��-�E�I&�����<����[k� *Mݪ�uR��v�]�z�:�8��{��R��׵�GKM��_!��E�hQ��f�Y!�i$�B�4�:޲��8��;�����Oo4u��X�墘�
W��@2)&�(�[U��i�qԧ��O��}ܽ_S�X�7Vq�m3��;�n۪�֮��Դ�f��Lۮ󹾥��kn��I{�ji���(��i��m2(���@�}��%���<++nz�`�qW�12
Ko�f� ��v��۹�=�Y3زsfҡM��h�IRi$�D����2E��o���xUz�xU��TO�(����t�-$��ˬx1G6��Z)�R[�����z)��6��!HU����
�$�A����ef]%'��s�8�u�ݜg��,���+E`Z� �H6�M�i�^}o�޸��:w�ji-3�jS�	���ߩY)$�)^��|62��Q��pV��#uX[�/G��h��m��iP��1m����m�vR�J��lm���b�@   �m��{uP*�ܨ�*��s&˺���w:t���n�Y�5�K\��yY��;zlNnv�p�w*TU*T*��  �@�@ m��*�PV��z�g�}+mm����2 �wMwV��v|R��w��� �-�U���������!������R��|���sGՙ��V���Ŋ�(�)��Mj��[����m��o\aM;�54��q|������m�C鱗��
u���w6\V�T>��z�I0�M�W�7Z��owZf��u�Ӷe}˦N{!x>��t&h�m6����1^���ï5�m������SHo��u{[ ���k]���w�wwse�wV� 
��nݬ�e��I��7�*���c�/�����V���pW�uD�A[m���3n��͓o8�T�!}멧l���L�w���!M�i4�4oG�+BQ}V�Wsw�y���l�.����W�c�ֵ�ӫ�M!�sR����]ϵ3�9�p�I^�LLP,$�-0S�*���@���3sL��=�3H_z��1�wUU�j���* q���{�-���ޖAsPw;��R���it֮����q���Ou�1�?'*]�HhǪ����� �t�m4��S�354�}����[�U�ϓ�]&Pi��a2ۭx!If˂�«��1�s�g�BI�4����~n,���!T�p�u2�,��YW�>�f�C�w����%v��c>~N���w6�6��m2�mׅ������0^b�
����<>�����4�m&�%�M�T�x���V�����m� �TإF�u�W]����ɶ�%���
�kG�QY�઱G{�c�m�s3qf�=^��Kn��Uf�Zf�ϲ�rߙ��n����q���]�eTxxR@mH��I6�5z*���:�[�S����˚C>�ni��Us�˻-u����P���ʿ��=��gΒ�}˃������$�	.��-6���3o9�i�B�ח-�����3��7���~U�䬥��ZT�뺭zq�������Wu� -� �L��?���)��A���eK��z�����n]N2���.i��UXiSI��e���YB���������#u��(��pU1��ba�L:%4�j�c�m�gsr�����!|�˖�̮vȪ��d%�K!��h%W��u(*���3{�!��/�>m��oS�����[�W5n���M�ަ��9���x�*bm������#.�}��-r6�-��I6Nm���uk7��v�@m���w�l�ݪ�`   �Ǳ�T�*��~���T�(����v̻{4���WGrw�]��U۩ۂʮ�m�mz�>��w-�m�U@�`U� �P m� ��*�T�����l�m"�lxܸT����͛�;��n�U�Ɨ�M���;�}�=s��V�j�ۯ����L۬����g�{�!��<я�0UMI$(oͶ�.�l���s���4�5��kF3��λ�_S�`�z���o��"<�M�B�+��4�3GM����n[��:'S�?s�}M)H�,�R`"�l�.��Q�%\��)-ŞRK�y�W��z46�M��I�K,d؎I��Ú�������³9��=��6�vln�wB��m�*7ym��[�.0�?o��?_ͷ۸���G.mo�3FU�i4���h�fy�X۞���Z�^9��A��o�Z���E�2lG$�P��P��D� 	��M'L���qKÊxN{<Y�dG.b�%S�]��l�ӳ�^��pǶ��Qo��m$�-��m�-@�5���s�^�v�e�wM��������2�4�I��kV�v�Ǘ�Cu��'�Z��t��@�)�i�	)���[mk���^�.l֎I�|��Rl2�j-������ׯ�zƽ�-��� �L�ۤ����l��}�mbǸ��݇nTZ�i��`�tPi�2�N�ձE���z���Ս���alI"C�su6oom���sewv�旳 [�z��U#E��&�^얢ӵ{�=�庰�/�$H�)��E�
q���Vd�Zw۶��C1�`qS-$RD�M֬kd��}���[=q���xY݉$1��Mۗ�����j-��X͞ST(�)2�L��	�̼ad�m��TVrlZ��OZX���QY-T�*m���;ׯ]�u��� 6�lR�<��ڷ�T�i��!��`�+V5�V��y��}r��{HJA�PM�MbR9�Z9!�ݒ�Zv#�R0E�i5@��Xݖ��l�o\��3`վ� 	I��d��ic�Cq��:����l�\1�(����.�N=cv���9�Z9!�ݒ�ZF�m��I��m$�� R��c�cln ��wm���ݻ� @@�Î^� ������w;>Ъ�+>v�|�u[g�n�'6�[m�yΦ�F�GSj�sk��A�����l�eUP 9{P�@U�  � ;�����-�!T�6�
���VQ슣Y��̇�إF�َ�S���^����l�*m��.��i2�-��޾[�n�Q�6E���Q_�m�%&�m��Zw�)�qz!��F�X��f<+���I�IPi���ʞ������͚��\�A�
�m�E7�0�g�l��q��/bI0�T�i"C-�Vf�t爛���!��F�X�����-6m�*��k�9��������δ<*��.{;�R����@��9������BI�L�lZ�RJ6YD2��͒��#��:�b�e��5Cl�m$�"޼�$�l��1^��K����jA�S-��m�uaݬ�>ǫs�a���&�ıa1|���!)h̐���h�	�f�S�?>��9qx �mkf󭱻u�wv�@)�[�����Ƨ
;)�?wo�������r+3d:o2\o#d��e��-"�)edصaݭ�9�N�j���4�"��l0�Զ9�E�{�Z9�%���Z`��i,�5KR�"Ӳ5���(��$��X4�����8�̯y�,9����d��m�m�������x���{+��� ��m��ҝ�x��@��L��}r�|���"}�}y$�vid��S	�[g�~�kqx��~Bd�i���䅤]6��i4���.���C��3,�G2��y�l�,2�n�,�\��z��\^nG���Y!���J�*T�h4�p����[��6��$�N�IT�I"J�I����L����޷m��zYͶ ��j�˦��7��Vl;��.���C��3,�Y�I��a|�6K 7[�i(��k6\{[�/7����m�iR�l�����ק3ZW��mf/�/�l�)Ja4�i��[#�D��C�{�v���^�a�I�)�H&�9��? �۞�/o*I~'*�n�-Fm���qA[j� Wr�*��UEQ� r��f�P  �J�Ru��B����R���E��Sj�
��^�EPu��ۊm��5@ 
mT���� :u��
� ��UR��6¨�U� +m��vٰ  
� ��@U  *�P  *� T   � �   �xzUs< 
�wR���Z��5�ޞqܕ����U��7QT ��� ����@Us{�`��C��   @R�� ^��5�U�-�q�=���=s\�|�M�mvw|l�y���ε��9ŶMq�8���ڝ�tҶ��u��ق��:]i[m�������r����;���g>96�{��R�;wGp=��V�[t6Uܮ���7���Su�㫭� ��v퐻$*�w m�[�Pol\���{u�AOlVcs��;����uz�             n�     ;�    �    ��  U�m{j    T J� U�  � @   �      Y@      `         
� � +m@Up  Sl � �
�Ur�@ Uꪨ��ްYt     F�wxUi�  �
̠[  U㥟��_��������+���< ��6-���[[br�/]�բ�^�    	�\8�jNP��\�gUSl9��C��s��uy���;��Z�Y��w���kSW{[v�m�<��lʶҩR� x� fP�J�� <�U*ll��5��.UU'����f�<�{��s����5��ov� w*lR��u�i6�,��M�����}y5�n7���ya��HPi����g�zlכp�!������=�i$�PI��!��nÈfW��G�^�z��)�)��m5�=�D�t��kӇ��; ��	��2�Ն9O��I/N��V}���������?�Q�*
�Pno9���kM�^�9l�36mm���ݬ��^~�y{�V$s+�~H��^��	Q�)�����l�����5�ם�N`Ӡ���h6�o�Z�^9�_���=;#Q^͞A�M�ۤ;�$�K��3�4n�Ďe{��f:PD�� �a���%�l���wpn���ƒL6���P<nn鲽�m�y���]ۥ�x��Ƈla��TZm��������|sl��6C��(��)��e�.z�9���V�Fs4n��3�m$�h�v�1��/�T��.�74�X���d��N�v��ӯnd�����lD�����$�I�Q������[5���bm�mk].�*�pv�䝻{U��W�����p
(��m��m4]4��x�{^�L�+2D��I��*2I$5�$��V^��ּo��@��:&�e�߈�!��T^#!�{�o�CM"K��KZ�_���f����!o�;�׏�>�rЙÈ �6[m��f�!U���@��uX+z7P!����°S�:�H��T��|���wn����`�m�
�%wV۹���[�J%��C'w��xh`��+��U�b��H]^28���ТSwU��F��`���=޾��])h�c+b��ѣ��>y
%4��)
��^*�q����u�h�#.�1��b@� �� ��l|�
�5wu��G��:�b���u򇻂J�e�m�I���瞚�N�I&	���W�?���� m���P��n���e6U�=��<�ʡT   �67��k۞<�*�)8����]7�MZ:)�֘[Q���]��Q�V��;:�w6m9��k��nø�w*��*�*���
�U*�w� � � m�*wn�h���ҋE6m�wZ��m�{f��v�7Vnw����T �I2]$	m@4�o�}��]vN̞;�t�왃v|A�?�-AF�N���ּ��k�"�ݼ��a��m�{�n3Xk*�e��̽�t+���9�\DE���ƈ	)*x,}c+b�\ �N9�X�+�x�{��z��E�� ��w��y�2m�%�rK�[�%���m���T�og����z�܊��
����m��+�.�71����?��Zv��n�v��H��Ȣ^T�M$�A75+;�T��4�/̇VԒB��Im4oo;&��:�z^��'���K��B�L������(�%���>=X<7fy\Aak0�9�@ZM�B7Z,h�\���1X}Դp���4�W ��c����N�H�i��-��[b��˻����HM���mmml�I�F�	��d���b��z8V�N��0),����DV����m�j�c�9���Sx��sOY�e�ߛz�tת��?<��4�5M� �ڸ>���:�cC�}�����5)`��[
�PAG^��E�I�6޵n�޻J�}W��g*�}v�v޻�p}���0W+0l��m��{����{[���7�on#�ߍ�1��9��|*
�_[�J%/�$����oml�ws�{׍օ� 
�����VJ�t�g�xT?~�� cg�X�+����a�J��1l�CH��i'I���AR+\.����G{��Z)�O^���Y�E!��y�BT���h&�����{����޿����m�<����u��*(=ɊIQ)��A4��+��^�S�� cg��s�a�N�  ��I"BǕ�2�^�������Y��1\TY ��m�uA���l��{k�v�V���UP n[n�umw�T�e��ei�S\�g$97�)�qx̓os\I*a��D�)����M�ڌ�g���Z�`�ƌؒCA?6�h�i��v��գٙ^.=������z�J�*� ּadÍn=�g$97�)�q{TQ�%4I�[lm�Mr�Ƴe��:��L����$�m����I �G�)Z�T{�
��U]�K�d�U۷u�[*�T /Y^%ؽ�ȫj�u�UP�fׂ1��׷u���^�b�N�[�N�H:V��jP�r�wA�c�lw� �Ul�    �  �� �*T[ R���T��{U*���)Qm��6�y����۽�koe�U6�M�v�����I&�d!�n�;5���~����q�|mD!�l��&{�ALjq�X,5��4x>ۗP1^��� �r��l���M�Z�Ӆ�|�>����޻K��տ&'g����h��%y��h
;�����0:봴���~|�m�w)8��q:�4��>T(�J��wPxh���Ky����q�z篩�������&ә�yT�uݨ�ާ�'N��\�Qwjw@A^��d��4�m�M������tE`����~f#�<��i}�}�&'���*e�[L�M�����K�(�,l��妓������=�,�|����n�ۦ�m���#=f뇆gy��'�E��[��R<9^�*�D��(�!V3�ɲ��6���Tx�eL�m�����I=z����M�d��wy��-��%$���9��v���k� �UP n�6�fS�Uܘ�K%�����GA���KWPXт����Z)��^�+��;)m�H'pRx>��P1^��h�A{����[8�
����Isa�AI&C-�<��i~�}[���=��>zjJ�y����G)����ߒ�ӷ����λKN糔Qd��@ �_*�[)���AGhѵ���﷕��}��@6(��m�x��Ín=�y!ɻ�y$J�M��,sm�;���njW-ݺ�vo`]��ɷ����tâ��@����E�n�;�;Q�L��׫Z�iDJ�I6�̔1)���h����h�fW�oo=�m�>h�@��)����6�N5��U�&�� l�����������TX��+w�iC�Z�� JL��$�S�od>��*Mh����=��$�m����m�4��5�;�ۋ�S� P��;H��A
I��)����g1x�ݼad�gq���5�m��m����H�����Q�9Sd$(I�-�Ц���ݞ��6jIrjG6��fm3E KM��&u�k����xjݿ0�n?ka���h&�^�rn����{S\������m�)��m�m��P*��qL[J̕����N�ٓ���²�U   ��ms���x�U �O_%@6޻��={N��x۷]=v�
�zN�t=UG��l��m����S�Pwnj��J��  U l
� j�U*�R�������mY��!Y���A�������ݻ���� 6*� 7;��kt��uJ�)�만�gݞ�z�k̓�S�}O�*ĸyx�I��m�J���m.+��S�w������W}�_S�o5����Z,�9
�>-��H2��!��}uO���k��L}��5�I���sռM����f��kZ֦�vl�o]����[�bq��_'^>����Ӎ��<l봴�B8PS�m4]4�����5��X-ᬭq:�5Ӿ޶c������K{y��ئک����f[b{��ճ=�7�
��S���D�R$�$�H&�
�a��v��5^t97v)�qL�(�:l&�`���ښ�E�d����(}3�)�u�Mc-2JI2�cRK5��^��o1�\N�Ms��[:��Ŀ[�kF�6�m�S7ALj��´Xky�Hh�y.]Ab�+{���
�\�~C�?2Q(�������P�}W\�b��y_
��)O��´`�׍$�I�v��U��{;��v��3��]ywjx Y�Ʊ�vA4�;�LAcg�X�+��U��S�+��
�Z4V�"Q��E��N�j�0Q��z+E1�\�<+E�����6̺��xT��$�f�M�M�bq��b�B�0s��5���u���W'a�°r}� �d��iI���kF	;}|*�:�Z,U�����^�S�+E�t�D���iP\�Y�]�7������Xq�������o��_��8�n� ;�vs��^�jk�V�*T �w[��Pݭ���$Q��^9���8PR���1��jNԎ C��m�
f�W
���/���s=߷���os�jλM�{~/ϟq�8�^J�I$"���c7���ׄ*{��xW��$����R��٬3r&� �6�a���8R��َ���{ڿ'�G�_����n����5c��$X@��E&C-��)�ӛ8�
�XS��#X<&�z�U����*�c�I$���-2�-6�$����V�g^wv������d� ZI�I��$���Wq�ΧDV�m�5�J�������.
��[-$�U6�!&�ճX,E'_
C�)+�,W�N�
�<y��w�9a�h	�	��Y{Z�[�4��Ƭ�͖�Ä�TiE6�P8��{[��ͬ9s[.I�j_W�kd�4�	4�M���
��][5���9_
c�)+�4`�����\
��� ��
�n��ͮ�]s:��
�l��ڪ�@   ��՛�laT�ب�SeR�ޱ�]�R�κ�^l��=�׷k]����qz�9���wa��;��R� 7Z� �m�;�l��m� ��m�l
�]͠[� t[:;�V����.�Ӈ{n���S� M"@) [ ���o��w����X8Xj{���i윯�+�:�kG���C��Z-&�-�|+Ål��E����*CV�OB��!��c�<l�T��e�S7\<+�5�18��j�K�f�X�{��S)H�]AcF
�qq%"�-�[e5|+��}~�׿;N�{�{�����m�>�ͥ�i�8�8V	:��Z��M�b�ٮ�=�������{�뷯��o�̣a���!Z<)��ʹXL4趒m�c�b��[��4絯AP;�T ͵[om=�����*�C�������^���*ƭ���kE���|)����,&]�mں�ƌ��>]Ƹ}�|�5we�5�������m��5; �h�
�M$�m3|���u����;��
���0xTW�
�Ս��$�y��	U�C���kÇ���1Wf��}�n][5����H�H?�l�i���
2>WPX����O�w�g_��Z,j�˜k�?%�$�m��R�t�n���z�[i���n�� T��m۵b�h"I
�M�%jM��M	��8�%��.�P%O��
�U$|�pz���kÇ��u���t�\AV$��)xI	��f�X�����|����kf;d����_�ޣ�k=�V���H�Ii6I��X8Xj{���i�8�8V�Xu�֏��;�^<9�Re d��4�
�xW.�pp�5�nu8�<&���5�ï��˜���ƒM"�!JM��o[>�d��wʹ[T� tͥv��s�;ؿcv淶�lQN��Y� �R>O���\9v��h4�%2���'b�Ƽ8x5=�u��/_wa�p����s5�&���,$�@���;u�<+�x>;�x[�N*	��s�xp����'��L��f녈3)0���n�8.����]���G���H�MP)��QI�;��w�����U�����Axj���c�g??���oY�����rov7ww���l����T[�
� �-m�wGz��ۯM��M�ǎk=�ߓo���q�<�����������:�T�x�e�M6ۢ78ׇ���u������AV6�8-����u>Æ�s%I$�dQw\,A����;�p<��b���v�k纮�1���Յ$�-��A���C�`}R���j�o��;u�<(��>;�x%8�L|�D4�d4]_*��5�Å���b�JL. ����Px{�{R'W�P  �J��p�T�UT�   
�  �U-�j�  �Y[b�=l �*l��ʪ�=�
�e
�V������ p�  �T�@��  Tw   Kb�Z��  U Vgt�[v�U� T� ��    �       �U        ^6+�U  
��P =���!�x�zv��[+eUTm� WSj�6-ր��ַ��[�-�͋iUY@ ��*�۫*l��mS 7��yZ7Ϊ�j��u���mݭ�wi�u�ojun���M�s��ǻm[���W{��z��,ڭ�֖N �yUp�]�6�۹�h�-���) ���WV�q���b��j�<�[+���k��Y{���l�/s  �+��m���.g	y�Tb{�U ��ڀol-�����U�M   x          �kh    �        l T V��(�       * l��PU��T    ;�   ��   @    �         � l �   �p ��� T�+n�hm� �P�l��p
�  � 8Mu ��l�@ +���   �k�����߯���� U 
˺����7-��mT�Q�x(`6����T  f9��ݪ�����ۋlmݺ;��^{e��m��٭�j۲��\��nݼ�'{�u��f�n�wU�Gp`s��UT*��` 
� w � � ;���T�
�5P��ت�}�������0;����{gn�op�톀lJ�ӻ̒�$�J�&Ia���^09�����b��1�k��_+��A᫽�s�`��w;̑A��e"�%:����S��w���K/GY�0J��w¼8xl�� 𬏖�I
U�����g����ߵ~M�������n?!���cEXz�HL�[M�W����\ ��W\,A���� ���|�<"�G�0PI��e�پ������6�ļ����Ӊ��������x���w���#ĒM��{�6� ]1��=���X6U �涬m���ͻ��cu�َ�v����|�m�g����|�
��3�녈<*(|h�
�	4�)�p1X��p1PX��>�wy]pb#��@���A
)��n�l�
����_
������1
}������p�}c%��DT�)��TRn�X���cCgu88A����o�qc��\�Q"�$٧E5�.j�X�/q#�T�`s���CG�v�;�����T;����^���{�y���Qn�*����	i�O��JA$SW|'Yz8W]��{��3u����m������N'�N�H���hQf�1�����pW���kr޶�׼^>q���x�:����(�D4�(2�������cG�r���S}�>aN�|+�7��4C��m�Kj�cG�ts��b�|^����v+����u����4Yt�%�Zw�+��x?�k�	^��|*���7PxAb�_S��qO$�����]�`m��j�0v�{�{@�J���ݶ����I&�C��vH=g^��=��/uk!�b�O��- �3l�,��M�5�p�~�<e��SͥH  tr��j-;GO��ջ�{��9xv$H���6�l4��R9[yY�c̒����K;�&�$�ެx�^{���a�Ǟ�s�kRL�I$(*�w.��N��7|�6�� ���ε�*�͉6I��h�ȷ�d���ܼ��[y�9�R\IL��m[7PxA���������kx�~p������_x�>���)���@(4�m�����;n=v�o*�=~}�{����fVo׾�z�=W�M0�)�ɤQ�@���Wxh��κ��)��+���j�
���d$�%��M��4X;���}ϩA�EX}��|>���>�� ���.m� �� �q�`S[UFJڷ�m\������V��VP� ��ʛyۻ]�ee�Kԥ@*�2�ή�m��v��	nvsmN����w8��V����m�02Z��m�ݶT�P � @ �_�}@;� �ٶ�,�۾���w
�[�>�}�6�6��8��.�z[�oS�ow�d\�T��4��M0�0�M�3Ɨx,>c2��5����/� ����W\,A�Ed�|�m�m�$5��د��1�w��5����^�݊�1����a
��-�B�.�0J�߯sn;k��S���_�c�2��߷�~A�{��2�t�m��J�����޺��y������o��{����.c��}�@#�[I6�-���Ə��s�,H~w���C���q�	K��xk�ĺ�bln/wm����jx�vj�7� x
�[g52I�,%I��h��x)\�z��}��]�q���y�ͽf{Ʊ�R��|��	��$Ju|>��'���{�PXў4��!�z�]��{8��D!m��f���N�1�����	�.�hc���~��nsm!N�e�u/_we�C�+���?xnÜo�Xų���h�7�6�"�֍^���̩W��3�λ��[�Tǭ���u3Ɨy`��=6cD�	JM��8ٲ�<�`��r��]�mr݊�Z��o���z�y����}Zܷ��u�^���'?+���58�R`�	2�A��}S�k7���|�~���:g�[�_>�}ᵳ9�� ��Ɉ��ɢ�I�M0nm�=���eJ���~M�Ɏ��;��쯠���޺���]��,!4�	$�J��4�������}���������l�"�w���_1�A�l�ۤ7��0j�������^�݊�1����`�5�9��I$�i&�	������x]�c�^h\�T��l�\��zb�t�n�b[8�< ��R������_��R�}xA����)��2��b�<g��n�hl֋�����t��P1��p�J_Z4�H���!�>/��@d�+�k����^���|��vx�mP`��\�0J��w��<1l�n����}J�;��}�W4Q)�E27�ׄ.ug��X�<iO��̽z.�h�|_�A����$6���L�	��o+�۷M�{v���@�J��eݶ�3Y�m�i���,p��_�pX��b�@Ʃ�78�<��Axk�zs
��Y-�j�1����`�5	S������8+�< ��R����;�� Zd��f�}*_+�k����A�5���f^�f�x�ċg��i��M�����J녈>�_;��CX}��}�x��X ���q4X�J�A7g�q�(��[�|����c�{�^��0l}�]A��ڡ�d��I��I�A]��UN��TU����p�����T Y@ݔ�f��l ܪU6ˍ�]���n���Z����͏l��n�q�*��ww[��k';Q��;�@U*� .[@ l������� �*UUR��S���R�S� �u��l��ykm�]vB�2��)��gt �ګ:�R B��������^
�~�TT�W�kÆ���򾹙���Q��L o[�z��RKJ=�����#�Z�҈6�e��lS=-�Qk�[!�{��:'�	S-8*�cE�#A&I6�-�u��Ԡ��k�o��oͳom�{[�����~=ϵ�o_��ݱ8�AP��m�H�>���vkG���p}��y+�,h�\���1�k���T�*fW�A�x��n�N���Ym�TVۻ�(��m�R�4Y)�p1���o��>x޳��z��z�ޭ���x����u�|�@�e��-�W��5N�7Z<5�=�k>�5�����6�s��z��=yx���a��h6n�X��j?�*�o����¸p����]p�
���G�4�M��|<;�`=�_*�a��X8x5=�u��/[���!°r���Km&J�/��0H2˂�A�fu��Ԡ��k�^�U�b��;=ͤ�,���I&�`:k.��E:�� �U*�V�[wl�̧X����X���<���a��V� ����Px\|_
��W9����-2i�u��*)�w��q����Ac��^xr����+g���Ii6�i;��+��>����V�}t�8~�g�����������߆��}~��ZXTA�"S���h�{�A�J��u�+��h�2z=>c��I* ҥ�%H5W¼ �/���CG�j��pX����|���_������D����n�+xۉ�{{����w���� ���έCn,��L�-��4X���+�\g�ugSo_�k��so[Nu��f�ֵ�W�~~q����i�����[�1�R�y]AcF
=k)��iD���M�*��gp���;��{��b����b�X��.!Pe4�@!Wu�3��o��m���﷎�O�4�����=Ə��@�A�Qi:	��ͽm=���3U�xߛN�o��~~��}�u��F
;=�Ri*m��kd+)����]ھi�2l[ 3�]֗�Jݒd�pxALo{�>al��W0K����[���|�����e3|�9N�|+�����1�s����% `��h�� =M�i�M%�M���^������k8�j����A����U�0t�R(RM�tSW\,A����A��d�pX�,K|�
�	}�w�d|x�m�Ym2�I7._I���2�÷*-jl�;|f�8�I�����UU�[�s�������+��VPVwUM�l�P -^<�|��8/W���@�Q�����4͙׷��.��Ss�-����]�z���n�wJ����ɽv��6��
�l��  R�l�� 7��~���[hU����T����]v�P7�N��I�T��{����w��m�� �R�Cm�$�KM
m�`��
���O�ŗ�� �_��A�
�^wU�b������H�m�L�
�	S��u��e��c'���Ab[��W0l�=ESI��I��A�QOs�,A^݅�b���{��<9Ou]pb���M$(*E�ZM�+�RD�F�>Ao]�׳��~q�{~5��M����EQi��)���A��/��`�=�w\< �FO��c'���Ac�<�%m�Vځw;�[��ٹ�ݻ�-���TM���Q"� �&�H&��0K����*)�w�+û��T1N�|+���E�%�� ���Ab��. �4�8�z��w��[���qُ�;K��.N�4�L��U|,AV���b���K�|*���W\,A���/C*Č�JT(& 	7pX�,K|��_r����;�b
���/����$I��[���,r����K�z�8�9��q:����W���ms����m��n!��1���Ǻ�ٵޮh\6� 0�$ -�e]4�M��b�,WoƱ���xߛLx�c�V��q�xgy]p�
kx�I�$�l0����o{�*>/�p��ܮ�!�E=��X��'{��䨰,�M���Aor��o���k>�ͳ��W��O�H �8� �L6�i.
b?=׽�f?8�=���&����ߛL~\�|��C�u|Zi�mG��qc���ֵC&�Mr��a�J6��q�Mًt����n� ;�lR�m�mU�ݚm0M�
:��1k���/\;r�ֶC�oNJC�*h&�M'HE�����_�����v�ߍc�m_=�~m�y��A�iSM�ФھbT�+��wx�h�%���cm�p}��'��*H��%4��h�O�8��;���o��r������g�74���z�G�TI��m��W}(��
��*?'��h�]0K��V�걊�4�l��,��̇����6���j��P���`�6�Um���z��I��k߃����o�X��;�녈0Q���cEX���PX��z� $�J�,�
����;�A���\A^���Ac�7¼ �_D�!�E�-&)�� �MN�p!`��u��׽~�_So_�k��f?8�;��+�"�H�_*�Rq�<���	S��u��d�z�Vm���e�C`���Aa���\ �#�;�xS���PW�t�|�>���l���;�w�{��s[�m��zU<�	�Sl�櫺 �@*��w���C�c���T (�nމGq��ީ�l�ʖ��m�;����m�4��m��ݧi��]�N�6���T
�R�� T �*� ��������bͷw9ѕ*Zf�ڥ[��*�;����9��j��v�:�/R� m��vb�|����W�?/߰�pb���r���J@��Vm���h�cz�4�,���Z<4X��J
�L%���h����)�*u�wսb�%�-&Jl�AV7�Θ�l|�
�G�n�4`����PW��Đx��m��)���h��{��xAc�v�S��+��+�AX0d�̤��(�޷����|����i��N����+�������� ��ؼ�t�	P+�۬x��[7[Ӷ���� ��إF�-���zQB�l�!3u����cE��Z�\ztu��т�\\J?&�H$B.�����{�=���o5�s~O�m���U�)�S{��b
����M�	%�V�~zk���[��f|������X�F܆�b�`�s�)�i�]|)<��n�X�
�<^�4U�����H���
�J��*m6�E7u0>�$��g���cv_
���S�W\����~o���66N��u������Wv�Jw|��u�� 
�j����ݮ�S+;^�����q�M�x�\��Է���|���ǯ��0V�C�H�I��	;Ї�.��XY�a��b�+��t�
c�G�����&)��i2�l�
�уo���A���^����t�1N�|+;D�d�Z����u�͸�=���=N�4��Z�YYm<c�]0]AP1K��*�L��h4����VNp!PxK|��X�����`���0S�!I��P��ks�cwVn��oE��T �5W[,Ў�WZ��;LMf�W���~���<)N��!��;��p�y���m$�%��-&o�xS��n�1�����c���ׯN��_So_���Miֽ�XM&�e�u�+��88AV�\m1�ͽߵ�&�x�ﵳ��x��s��i6� Q���o{�*%�b���1�)�����:`���4SI�����v���ʋX�+N��C7/�4�&C��j�m����{�۱�ɭ��d ;��JUw]��[V�7V�&y�xd�����mn������$Vh��ERm]p�
2x�h����AaǼ��1	}�w\�t~D��!I6�%��+û�A ��v�^X�݆�X�����]D{�4�M�A����T�Z)�<��.>/�{Z݇VߵA��t�E���6��-�����8�ٶu�X�)�?w�^���g�  UAT
�Ҥ�T
�TU� �ڪ�n� UT6-�b������ ��2*��� m�2���[YU
���� �����@�R��PʠU  AScd�  s-����:�
��[`UA��� m�UP*�F0  m�@    @ ��*  
�� �/T)��T�� 
ɹǷ��^]���vwW�V�5@�qT �� `m��������*�U��l���F�\�@
� �U  -�P�Qջ�Ҝ��T4��z�w�����������d+I�w�����wߪ�m�wN�QV�Y��;3����+(
�r�7]��ι-�{��q�ۺ�As'w�����Pg�׻V��Y޽�������V��ٷx��[[y���@V���ml� ��r��A��l����� 6�� x*�.Z��.��s�@    P      ^@
�T�   �  
� <�  �    �{��u�P       *� ��T
��R�     l    �m�       >��P         ` � p   �P S�T� �
�iM�P�@U
��[�� n    ��pv� �6m�� m[� 
�� �Yu��������W�T����U�w+L���<U�-�l��ʠU U
��ln9'��j�m��󹸪���{v�뵨����eE�d��|+����7	ʛZ�Eww[ڎv����w�ʠ*�*@� �U m�lT� �j���
��Vm`f۸ƪ��e-ݷ�6x��m�rowS��{Wum� ���]vj�u�!�#����������}�|bW6x�������y
lSm��\A�a�
��p�h�����~z�=���󉶻�֖�V5cm�(�}aml�|*���W\,A��~OE�c��� ����@�I4�"SW���;�A���\A^���A`��W¬A`���m�4�h6S\���N �%��+G����Ƌ�`���b�w�6B`"KU6Ý���c���^]��b6@3�۸��UkJލ���ۛ�j�']��w�ߓl�s�u0Q��z+E0�m()A�����<+E��������U�Y�:CX����Rt!R�i��f���ߓ�{��g����~.q8���
�RT��HR
�=E�Yi:	�,�[i�x�����YI��;~���er��uh�Z���&�tKI��f��Hs^������k=�&��߽{1�J�q�]��}�����+4FU���mt�m���\��[iJ��[Uk��u�Av��w��Cvr��^��u´<5���`ڍxHkEN�D�!��M�M��DR�`7�wWn���n�(�_}�`KԘ��4覮���K{����96\�V���_
B�t��]A����ē^,�Re�i��3Mx9���vq�ư|�w��
����+��3a�e�e4��oG�kEC~��)-���u�i;���<�N�]��}������j�f�T��w+g^׫my�]�ͅw]�Rm���]j�ܵ�W=����o���s�u��g�)�`�1M���RN��xIc4Aa��l�ѿ����!�~��B�T;8�q�
&u���><XL�t�-
Fm��{O&{��Z�n���ChRJ�m�
'ٕSt�F�{�v^g#�z4�_��&�A�/c���٠�Vf�����p�h��-��T;��ޞۻ�t�owzZ�4.j� �wsu���AQ�S39��(+EhR��֌�k���X�3�{��<*�.��HP�E"������\T�k�}=5��Z��;�qc��$�>M�@ ����[�+��f-����b�l�XH�m��-''������ՙ�ܼ�آ��$`�)&)�yr)[�$gD1I�q�OZ�}$�$���)��n�I�U�[[U�x *�����Y�G��     <�xe�5q�e��-��
�9o.S]��u���
^mSỺ�[�u���y��)d�ғa��`�UU
��� P ;�� � �����UU xe;u��α�ow%[�� w����5/Un��V�R�v��V�����i6� Q�Ϗ��g�آӻמS`�z��[��M&Jlŏ��ѣ'�J�6�n��7r�d$ �e�mѦ�3�e��%I"����h�sx���xp��U��٢�m4�6��X�xԓ��*Ʃ0�[5���9_
c�q}��pcG�N~D�A I��7»�`�~O���c9�_q�,5=�u�k:R���{󿟟�o�ۃ���z����v�;�כЮ� *Y[j���]˽x�cn�w�>���һ��Hp��{��<+��|�5�����<3���)�M��i������<��U�3)0���j���5�����1��\�>t�-6�)�n�1�98�w�za|�,����xp�k�� �5����Z�e��p������;�8�����p��¹N���\�ǘa�@�]"R��<�|��ׇ���u�����\AV5I��~5���Ҧ5��P��l�fF�;���
�P���C$�(��m�H��8`�܋�A�O'���XL/��S��q�<�%� �4�i�CI��Axk\�T�����]��8X�=��޻N���/�Ӫ�u�~t��/޺��+G�����W���u���Lp!0�Z$P��-�m3pz�����O�>߽��������2���Y��n�$�6RI��)��?p�c꺁����/PB�o�o���Z��!��M�eo*��l����nۼ��uU�J���nݮݞ�m�i:	�^=9��un��-eG���k�\[0�頝�d��L�;m�݆)��D��H��a�H��m��LŎ�2Fb����xj������0�H~�����-��-���R,j��X�b��N$?9z�����q����&rII6i�M]AcFa��ALj���?X{'+�Lp��܋�+�� ���,���-6�L ���c�7u�����w@M�mU�^m�꘲WH{�c�������b�X�;��X\���4^��p1xd~D�0��T��~��^��HAc��Ƌ�p!!�����h��}�7M"Km�����h��_��3ƗLp!0vL7��Òq�����@6M�A_�h��}�_���Ogկ6�v�Y�V��MV_���xj?q��L0M* ��\+Øaxw�;�c����[�o��I���?7����ߧ�P ;�m�ʧr�m'�v2� <U%h�*�ʻ��z�
��  �썐y��@]ԯ^���׳V�w���z�;���V����5ۭo���mLK(�l�efڨUT  @ �   m��+�_O��{��ou���� 
�[%[!AU�om8�]�ܷ^���u��й�ʠ��v��w;��ߨ�<���_q�/���녈3)0���j���5�{��a��E �f�S0u�"�xT���C���W*gc��^<'<H� )4M	��Axj��8���	A�T�O�X�c��xS�H����H�u|�5�����<�|o�ׇ�3�녈3)0���I0�<���M\f��'�Lp��܋�A�No���X:a\�,/�=��l���]ʠ�e7n띮��v��J��R�G��]Ē�m0)ZM��^�5���������7���m5�_=�~zw;��m�+<e6
i��!ں�bS�����1K[K9H�9�Ƿ�B2�i6�&b��;om�آ��@��^�"��^�m�i2�kó�g���*-~x��m��=��x� �"E�[B�J���n���w\�OT��+�k°~}ߖ��%�Kmh��m�U+ʫz����ooe�u� T�w6�ۻu���t��K�E��,W�k���CE1�v�f�T2~7�����+G�r|O&ۤm�
¤5��˂����s�X�Ou]pb��<�N����#�)�B@�B�٭L��r����{[<��3�ٶ]~l�&x����h���!S
�m�H&�Պ���,W��I��!3v��h���w�V���I6�)4M�h�oq|*CX'x�hc˻��k��������������ڨ�o�v������;�@  -֫��;��J���wϽ�<������/���8���ճ����_�Hj��0�M�-�%��������S��]���Y�����If�z�`��m �y��;����Ⱥ��Q�n���
�������xAA�K�K!�L������k��p}CjbCX0t����Ž��G�Vl7�6�%PJ�!!�:����2r��� ��=w�=f�w���[m�a��)6���{�:��׹�[$ m�lT�.��.n�E�p]���jN��<"��n�1Tf���l¾�7x��p���ھ�q5^�۔���{7���:ۙG>��몁��%��¢�I�Im��]ӟ$5β��2����4_Wg��4z�k�Ǖ4�`�d����V�w���5����WU�]���4|���bCX/��G|�a���T�t��kwe�F��]�)��V��֌~��l*YOA�n��j嵹j�TB�+@���� � ]�Q�����m�[6ު��mw{9��uܯ�����Y�nf|�˷w;w�M�-�B����oaM��t;��qT
�J�P� �m@`U � �j����}�����4�@ �Ъn�.�f[�;˷[X��{v"s� T�ʷ�\�]6Sv����]�l�+�>�9�BCP\�.
��NW�ׄ��&��f�	��4z�,�/CY$�=f�xZ�����/�]p���"p �RM��d���Ć�N¸U!}��}�'�����֫�h%��[m
c.�ݵ->�"��6w$5��pUXՓ�%�L�H:)��k��3��=f������x��Z<-l�uPxou�I&`I4�M��0a�sY�w��g��և� USg����304���\��|[��bCX'a\*���}Ƽ �j{��4?�����I4U�b���=�:����a��v��l���g�ΜN��ǋ ��m���*�j9_
cF�;��<(���1U����:��>Qi��h�7U�ú_U�4|���cExox�*�����6?siRa��.�W{�z�{����+�]|�8����;��9ou�A�w4��I��i�{�>w۬ok�\�<J w*T�<�۪��>2�D�]\h�wS��
V�+�V4`}S�u��0Q���c�7@�U	iI�SW���Rq����{�U� �I��cExI�_�b'��-��%�����9Nˮ@�=r��>��hX4V����h��<`�
�I�A��gS�������>��V�O�Xѡ�N�� �Ojw�eS-��l1���f�s��o�&�3չ��Ͻ�����'���\�$�m����m��k�m���fս��j� T�k�ki��®�K%�|>�S�o�xS;��1O\�H|ǴhX4V���.����D|Jn�������
��3�Ř�N��Z�k�^b�%��N�qo��w��Z��O�umnn���l"Q����M>�-KRI�u,[E_�5�
��E������/�I&�*y�wڣ���mݹ���d�w;s�kF�x��\�@Cm��l� m��ť��${{��/}�v��O�L��T�"Zm�SF�>^����e�jl�QkͰ�,�!��-�8�Ja`��T����4X���PTW)��CEh3�ņ��D�[��0J����V��ӕ� �FOH`��a�,T�������
f�-�Ǿ��g�Mfz���O�{9~t���v�5��G|���m"�m��ll�����J����*��P��m��^�]�     <�x���[�m��y��۰��{%��j��d�X�Z�C�EwJ��6[�1�w�� m�U@� U ��  � ��P�������ij�����s2���śoP�ù�v�u��\��x
�P�6�����Ȕ�L�׫�c�����t���%0�Hj
�Ի�LAc���*�_0�D����BCZ-�u´xmk��5��ړ��4g�-�/���iF�Sm�M���kE	s��!��ԟՂ�v����Έ�o	�QC������=�f�0^��pT�0�$?xJ��c�{�>鶓d��W��b�l��l���xes��?AJR���1�<k}=ͤ�I��&�M����.��=�����oe�U6�P��m��j��^|�{�-�|+�!w���?XrN��:�1X+�ap1!���	�m&�L�!X�g�?ʡ_�#����4^��x(�/	����� a4�*�w����W��b��S�	�6]AX<2��r���+�i�i�N�j�4g�.��B
`�1\g�zr��]ȿ�Ѣ�	(���m�Zi����T}���-������v�^�չ���Gm�>����,����V�l:,M�r���������C�� �k������w������O��??;���m�~�ͼv��}x�̩z�xf�+�:A��L���h}O���0z�.�. �L�7�֏[8��`��~f�,2�l2���ƌ�s��q��'����N�}ưp�k�����:�6X�2W.=D_vzmL�#î��vC$.2�(��h5[w���#���d=|$�W٭��}�~m�~��2 <��S�c����_*�r�l�۞�vN�U�-��o��O<}�oZ��޽K�z������g5~m��{�_q�<'a')xѦ�P)��ƻnS�����0t�گ���,u�<+��HVR�QH�w�	ƴ_]������˺��}��CG�����b�(�>I2R "��=f�xZ���}Ïr�U�v��_���O�Y���W�l���$�&��I6M��5����:���էH�����1�\m$�	&�[ol���wog��M�[�Nj�T�6���M�E��L Q��Ə
�9�C������g�N���F�q���枿n�wl��F�I��a�������W٭��7��0o>��h�K�8�k?O��l�,���c�3{ܯ��
�]=���vܣ�rb��
�-��ku�p�h�\��$5��G�7G!��e�) p
a��I�M_�h��[�F=J�s���;�K���:��/Y��~�H�b���PQEU+!	
Z���QK�Lx��^[~��(��Q)�QD�,�� t4h��rl��L�Y���,eR8�ĥ;2�LU%&2��PXʂ�DLb��
�2�B��I���©�)5�Mb��(5�3!Z�Y����-2)��%�F���j�xo�;rR�]'^�����?�<\�[wt����p��!�C�b|��t��N�0��wz1."�j���e(����ϧ����ʗ���_!`�j�R�ʼ�����{�􇼚�uC��z0�臢���IE.���o�P��و�8Mq������r}O������ܗ8{���̌�U��6���;���՞��Y�	�TJh���RQ�ت�ޙD��6��a��Ō��Hvm��w���{�/e%����]�>���u_`;N�uC��..���ޖ� �ie�����g��2|s
QKю:g5y���'�S��n϶z�V��p��z���į��|}�W���Ûƒ�\���þ���|_\�×(p������L���J^xz�(���u��W��c׉��-!���\\Q�]m�|ju5J%-�9!�W_�]\j�R�[q�i�<67�mo��4�e��^�#��)E.������Q'�`����=%_�k��O���~~/Z?.�h��ۭg�;?'���7�I(���{���IE/���C������$񮣁;.�L�՚0Z'�!�����p�*��ڷ�9w��(��S�M�;�Ϩ�t�G_��q��n��h�#x9C��2��_���͟��Bk�����^𡹭���j�!�Fq��{�,n��f�Eˠ����H�
L�=�