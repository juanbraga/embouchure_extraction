BZh91AY&SY&M��ؖ߀`p���2� ����bF���K�f��li,V���H�u�lA�C�:���"����d���,�Qu�	�	 M�6�УCe����vSA�@5� d�� -� AB������ݎ���(@g`j� ((�m�
Ӑ Qѫcx     �T�h�D��mRS�p �`:׃�  @(  � �p   @ �  k�GG{9� /{�@Qհ{��AݚSG��^{��(��=t�V����oRТ���N��uB�u����GZ;��n��d��ӻm��vt 
ȭPh(��@�i݅	Q\-Wvt�;V��ْF��)IUJ�eB$�j#9�kU5��M1�6ڵƔ�"Ơ�Z1 cV�[@IT�l�d���m�a�ŦX�@9�B��]���NP��Z`��6�kcU�M�m�5(͐ҙ�e��mT��۲�iKj�)0[mRm����օ*
6VŁ�T`mhj̶��S�S��P5f�vʹ�h4P�)��BWM��mTb��J�)*Y���[)U��-��jK[f���@�jT�Fm0��bm,�%B�B��ՕZқm��q�McM�������.�m��ݚݎ�Y&��m�hkPZ���(��;b�
̡�`.��M����D-�0 6�٬uv��Zkb�MVX�k�]�@�aY]AD��1 ��C�@tc�WL��w���:u�b��*�J,h����X6��j���t8��[6+fV���[6�*�lժ1a��m
)�Vh��TbN��R
!Pt��H4�*�ٵX�����U��L[�R�i��i�Xe����hXa��mk0�6�m������a4ʲ���e�&PfU5��hM�[24��h�vѲ��l�һ�fu��J�*��M,���Em�VT�d���f
�6��e���fT+Y�i�*k��E��H�5M6�wU��TWq�� ��4
�ӻ9�e[Vb�t�U����Y�I�B�в�h��-S몮j�+V�X�ZZj�,U��'A�Z�e�L��Ŭ�2 @t���	t�*F�E��f����6�h�f��b�	�h�J4���b���v�m�@E�M�j��.��ـɖ�j���Kg�]m"���� |E?OER�     "��I*UC `           "���I@Ѡ C@ ��hj&S�I�2hF�~�i�ޥ=4z@IQT0 &   ��{��|�c�����]w�#F��Y޹.�u�]w�}o�Y��w�|q�������ǜ����(��`���{ �"�0DDW_�""+�X������~r
"+���DW���Z���'̧3 �$�u��f"&��A � BH$� i� ���3Z��Z�={�o;�3z��5ƨ�)X���7�Dt�R&��d�����$
(��p��		��Y�jV%����nݛU��1��\���d��� &/��v,�זm�5�Q+Q�F7u+I�m�æ�]-Ie��S�A�WH���nk�Q��Fާ9V�=��ݹ����6�B#�H"B���s��-VDYJ�.���׆�dԢ��{�f�C�f�d�"$2emE��(�ژk���o(� �F���ؼ;�a�&YUXF�	�ۏu��I)t�3"�Hƌc�ڲ�1��)�͊*�7b�0���n���v�1�kg^����wx����
D*�rC��)
54Y�P�7x�T`�ohh� Ɠ����7�*��3��`n5t ��uʚ,�S&�4獧��NL���ma*ow7To,�X[B+�����Eei�a�ӹ�k�j��V��xSǸ
�U�"G��6����-��Y�.��{�_c��P�of{fI�]�&��摺)]��nMf��Ǩ-pG�j��Y��̓6z5��\��	�Ɖ�Miԁ�:D������?!�lӨ����G�v�@��&�H�@4tН��g)êx�c���n�_W"uf��Dl	T��Y.�C`��L�!v� �u.[��B��%"tAT���JȎ�� @$!F	8@  \�
R�$�kn��E���cu\̛2�d&ךΝ�F���Tde�����SV��(nL��)�َ���Y���W8��0	b���ee%]�/�.��g^�������Q��ʉRe��f~��Y��j�� _L��v�X^Z��![GB[*�.��Ȣ�.��Z�t�4#:�Ʋ�,s{]�L��˝����4���̚�1%��&2�-Ah	U��X.a6\�X*�E��ոʉF+�r��V�C��ՙu����{<�e��1+��f���$�e���"�9����p8�fVa��Hm�S13{��pm�яn̷�or6P��F$�U��Y6U>.qI��2b��/&,٬`+����^f�+���ej��un�t������dFF`+��ҋ�.��*e9z�����U����&��l��d��Mge�u2zL��N�O;R!L�6�2K����P2\-�q�v�*�Yw�C�&�w�Yy-��uf�c6�*�:Լ���`]��x(�����r�!;q;���N�bctX��Y���U�z%��miuw7cְ�k�Vź2�8e-z��2f�`�A�u�;X�P�/r�k���eb�kZ�]%sZ�n�{���Q|���/�1,*��דC�E%�УKc6����e��صN#&��,�ҩ�LH��ײKt誅����K���P�J���4Jȩ;o�˸n	�m�&�cXj-�����fj�ͽ��V=��dM7S*�k3]��DQӶ�*�Xk��mfOu�,�\������P"#�w*;p�Da	Q����$V2��BUnHK��J\b��'rBn����kHP�Ek�&�b��"g չ�\��Ɩ��S�?l����f��K�mb.��Ĳ�%X�y{�TJ1�T����u!a)Aj��	 ��-�o-^����+u&J��&)��
:h�}}��n�-:w����ܹ���ӯ�i^E��7�+ls*n�q�V�J��B���.�/��v��Z�d��:u}�8��s[��v�I<�]UV8��x2u�#������S��j�ɕ�����J��	�M���;@i����ua���)�C8�O^��&��&����J+FD;f�F`��wU�3UK����e�x�j)��	��6em����,~1c���9/1A6���]i��a�ԡ���vc��w�M
w�,��m���.�VAqV��v����]Se]ū+(�� ;�������w�/�1�GI����o�ҝ(L#�ifT¼.����ͨ-�1�
��U�,8�TYY��+ov�;�����YB̎�����ٗ��%Z�� ʲ �ӇD�¥C46�
�H���*�)�ꭱ`�W�?�l'j�&��ZX_��sr^��W,�|j���|M&
��S'���˼/2��I�ɹ�9���-6q���k�񓕢�6ӷ8_]^�-OXo�+.Î�髰Y��a�-��b�kb��A\����gE�c�����ʜ��S;;�YUΧ�H��joLq�@!�!$�!Cl1�!�d2 "  � A!B
"�K!2��
�2�$���C	�HDwI9}%v�W;��u��i����+`�+[���/!��;�	�4P��&h�F�d�� u��c³j�藱b��M���h�C5�,R��Q�+ZOvRyo1�Y9eFIwe#Si([��$��K&j�v��D茋U������h�.NP�h�%�+	�rڹ��̒fi�t�f�6Q�Q�]�R��t�p�b�A٧f`�-�v��lCR�V�%�f�y�R҆�3 ����� �/K�ZxE��R�Mڥ]gutق�6�x^J̚��lX�'E�mݵwr���C���\�jeq����ft��j\�UV�.�BI��Jm7f����T���Lۂ��j�I9382����5��4�l�a7�`���W����jK���z�XԷ�%�
�H�g�t�7&��Z0�����0���l����d����4*{#�{����3�uu�e��U;oS�<fY�y+��r�wZ3\җNs/iNai��B��i�b��"F��b����6"m�W�[/0�A��c갲��Ԅ��#�T.~E���6�U�9��dJ�x��Yz(�[��/0[8�̱�0-�
����!	"��Y�75@�bW�SS]�r�D[*be�W��-�7p��m�V�Da%�הl:o-
˭�'Gp�t켬+����ə�&Tes(�xf�,ki�u���h�)��xpU�S�Iv��5?�ޚx��[Ai%�Tg[f�e�n���T-�W�䞤o4�;҉T�����G�զә��{�����e>uZV�:�]ܕˑ|��5��7�n���A\�]N�S4طr�d��*���9����X�Qi:V���͕�n ��JP�&1%�%�JN�K6�w,��ɻy�e`�Q
�Y	H����5�u,�	���A6E��v�E��-����t�zRbVn-6�;3�
�p�����2�g-^*�'Ky��V-�^
R�U�3Lt�)��`&f�;G���]�hSfa�{nː��J��v+)vq4��j����;J׵"��u�nayp��,[ʴ�s.R��*�69Y��e#i����cR1X�
�T�oN�LVB�B\D�ۄ�)!;��&�2�!QS�A����4�P��h�B4�Mh�9�9��	���n;���&�i)���+UU3:����%GUvٛ���� а�6�v�(vU`A�4��ֈupJS���w#z+s�[�3/ynX�`��
��	1D4!Y��*�I�M���f�gPf��x�8�Ƥ�*����Sd��LG0nK�0mS�f�H��̺R���ok4�����Q���1���r0�њE�Z�2��7A��˻���*P�	Y�� �����J��$��R,�+r<wk�5$��ݭ��TJ4k����1��h��sPY�a�/i��؉�m�MR�ٖUn˛�K^�K��s��uJ�+�)��M����+�&�^RӴ5������e��أ)���Z���[;r��X6)���+d)E@�\^:*������P�G*�Ř�<�E�>���}�uY6X@�S�dһX�m�+V����x�J��sF޲u�T2�82����f[���YeJіt��j=�7��)��xn���B�r�%�0�ݞ\�so�ы9Xg*����}���
�.z���b�ܸ�ǙX�ڠ�B;�/+,h�թ�����"��-�%]"1IR��5Paa9��A�-<�K�+"[�P�db�I���he^]�j�X��ejY�0��Jˌ�%�o���^d���˩�V9�eѮWb�y�\���oVӽ�Wk̵4#�b]��n7eUeݘ#Bv� ��T�d�� ���"�8�Iux.V��`�����k-��6���f�wE,&��7`�q7P�R�]arѲ$��լ���+F���4�3�\�/;�AOVn��Jѱ���֦^�)��Al��7Mb�.^^�ˇt�"Q(&n�H@a�MH%��*�B�P�0e*�A�V�H�s��s�9x7Z�Y�}q��i������7$,��P��r�+.�#��oH;�̖�����xÒM5e=�+)8�t$��Q� /v�.�Y��uJ�r��J!$
"2V�F�(!Ԡd%!K$D!@�B�W�Xr���5p��"G��+h����L������R�2�(����&-z�Z��\��G���m�+7�ì]8�4��U�;æZol� ����X)E\]��I��[�e��<�]b�;����VK��z��*���zh�yS���D�3";"F�Z�v�����)��3j��ŻY�.��j�2�Ct�{��B�ʣ1u:������4R��3��ٌ!,i&��$B)U껪��4��!�Ȇ��)�o7�X7�8D5���p���-�2U�M[۷��l�˴�awB	�!U/dX�����c�uWr��]2nЉ������Id�Ιuw�3�����cg)��E�OV��vg.����Y3t�
۹i<�6���q�y.͒��F��2�Z�y5��a6��d,�V[����t��ڍ���z�e��,��$�+2��U�7Cn��R��;ˬ��)չmroE����Z�U2�c��ʕ;�,����� ��c�B��֤�u���4r�62���.�:��~��ܶ��i �-F�	���Z��n9X,��:��^8�䖝���-�:@h;.�6wpK���\��H�v�)���[�a�r��ʍ��sY��.��X����)��p�FR��CU'? t���/&iK��g.�dS�	�t(ێ�@��Q&[�����Lb�t�ǍȎ
�j��Q�eܫr𽙗M�åmy�)b8�1p�"<)N���R9�ZU����4j�&��&���zƤ�h�OoY{y�^�+2Qܼ�de�.s��1p�Ҥ_>��.���{N�P�h�:�6�f�m���d��GuM��cT�[j��ڕ�m��n�J�pm�Yr3�3?LU�Ar\��s!�r�&�Aӽ���F\�R�+�-��[v����2k��z��������$_	2��eڨÛ�4��5w�S� %��R�[�nsm`,��[56����ݎɭع:$�<�]�uf�έ"��/6�UK�dC�v+QV�oFI�-��a����.�]�Ս[� ]Q,M��)c)bA♺8�����c��N�Y�eI"V(�"A�*�9�W�o�s	WQD)](Y���Y�W3��%M<��|d쓜��Ɗދb�7r���y�s�y���B�W*��&1�4[���%\n�N�,7�b[$����<_��K�E;�\`ܵ0����e^�U6�aB��҇������B�����G4�2��td{�Y�=ӎ�� �D��l��'LCF�/YM�3cn�քM����̽B�hʝ�2���ju��t5h�$XsV2�*P���SR�8wPt� p̵� �W��B+i���2��#�$\N���p`�E8$�l�r/(�D*�\® ���D-�]u��*�4�5/q�Z֩��X��w�by*�V��t`cMu5ڭu�+obV�eqbowfX�t��SI�vU�uvr���n�z�@�sA��Q���W��.MX��{gEj�r�4�+p@P�W�S��K6��}:��<�t�k�[�ە��;!O�14r�2.�n�j�،����5��TQ�5]W��.�Rq�8�,����A	F^�1+s]�v�ܰ��Y	�C��,NIb2�W���$Ʈ�]�oHW
ٺȌ�&f�I{B�mh%��E.�n�k��YY��jV�4BH���(M�)��0�j@9
�Y%2�Vmlf:Pę��krZ��K�{[�T$�fg�8�p�O�0(:���4���_}9%Mo��ۃvQ� ���h��Y���i�1�i{]S�¨�q�����T;3SW�����W�ג�lTsp���R�?�1╶�	��DV1d5�<1���+F�z,��,��Ȓ��M��VU�Ԍ�e�(��ۗ_��B>������E�����=���/͇'p\`ɪ���jS�5q�$
R�U�vV׊v,�?�ۍ���t�R߻�FQ�ʌ2�?���e9=�ݥ��˺2�����5|�M����K�Of�>6��O�l�X�R�KU��d�7��8V,���x���l�J2��$��4��nU�+8&u5��]�=q������n#�������Q/��i,����SZ������n`�[�Wt��+��dH�=:cV枎��pfe�Ub˥`3Es`������B����i�:�&�K1��[R&-B�'u��>^b̷(��l�]�H��D�KXVN_�_PEmK�+ں��$�p$0�GV�C6���2څh��>w�уH�va��4��Y��K'>���k�ҙ�%e�N����ܬ|����9���xe3L���D��y6�����P�@���Jf5�-���Ac�!��L�*��sʳ�z��{2���u8sF0�6Q�\L��q�l{'b;53��Z��S�k.�ffr$�7n�;[+�<k8K�o[2
s�f5o�3l�λ�2֥2"Fa)[��\�b�9��P�[�t����q��Qp�
�5���Е�t▜k��칖���骼�6�Q�_=�^5o%9o���~�XM��ӥ��b�>L�ۅ��F@b}xbwؔ����:B�]�yԲ�m�ݾv�����z+^���=�erl��M�����s��^n��j��XJ�w������A���v(��U�^�
rG��})���Qfh�v�ΡKC�43Jf�$�H�e2�v�t���\a�{-~�Jv��G��aj�e,�E]}�KvM�:'����2���FC�e_�"t��
A-f�˧/r�����>�%��.�KG�:�d=�gJ5}��	���ږ� .�u�ٺ�8tq�WW��6'�f��z���P)evt���<`ܬ	��J�"eE�"���|䣛�v5`���(�J��[�ӉN��w=�a��oTYέV$͊ZL�D g^b��R��l;״���F1zxS�Y$�]��u��"F+q�P����{^�����/n"��֕/�X���5K4~2�p�wg��6k�|�/����䳵f�rt3��Wr�o�nL6*�ܦ���dZ7o/�nSU�NZ�J�b����&$���[�Q�͘�Y���:�v�9�Bc5�Y(��aN�-+u���Ư{D�S��qJ*]��8�0�h\Ո����n�ݺe(�l�3 tiQJn�3s���k��MC�Ε�n\�NA�=�s���W�Ǉ�_^��.5�-�+�ݾy�u�zp���D���:�5r��U�̩��o9�=@�`���W8�~�2&�e���Y���x0�P麉V�����rS@��扽�Ι�lڳw;���9hph度��{�Opk\q�K�25��!��
r3֝���H�Zt�/!V1�h��36�`�w�U'����⺻�H�V�����H�)g.���륻;�e�B�4���4Z�����ݗ��<��սX7�v�p���d��T��TH�X ֔��ڭ�������`j��p^VF�`�yA���u��y��i��ɷ��3��P���{�
к�/7R��Z�9u���k�w*�h��� �4HS�Ύ�m��5�1{��>��y��g���Ni\�Z7\7�ŉW9��"V5�4X�Ϩd����������yo�6���(.c�K6:.�\!�����X`P�Z'B{�0�Ra��QX~c�0��oN�Ԕlm�(��މ����귦@\áu㩯�(^l7֡�e�S{_v��mee�Q|�3c�=�_U���Wqw,�4�!�;��9r�nq��XCʏ-"�Uxg7rVr�z���$w���J+&�쾡�]����^�I����J�"u[�S��NU�DT��׎[,=*��픪W����gAw��6���1���)哸e��y�q]�����tr`!n7�������vۂ!F�f���թ�N�M��G���5�nH�r�S���;/�k,dC'%��A�R�=�98L���p �X��`��Q��7�U�;}3��[�vq��-�u�_ ��_>Z]=�Q`G��o9' ۺ�Y�,�Vj㝙�D�Y�9E���������eД�`a��eK�����uZZ̚e�����.�fv�I���y�f���0]��"�:�@�u�W����t7��+$�E��**Z�JDn�*��ڟ<r�/]���ͤHԫ����U���g_�V�q�z�1��f����eѥ��~�ݲI�wkz6<&�yKy���f�U�A�G�!�N��>�\�[z.v]-�[X��LJ���o3�n��D�0�m��b�WFe[͒����!NToK��=Svvɗ�ve��9�
`"��u�n���y����x��~��N>:��Yt"R�E�>�ڒ���s�̡&]J\g�JY����<�ث��s�-���a3I�W�� �J+n��k Ʌ���ٕ��O;3������8h��v٘��ܥW�wr�z�[z@�^�a��۩W
����h�ٹћ�Nچa�9ZK�7G���Qɚ�l�j�c��g�d�g\��jA���\�#�I�V$ѝ���/�ϫD�B���;���C%X�u�#CE(��[�[[��n�����o"����\����%^!�p����� ��h{(]�i�a�N[���fk����F�gY+xl
�b�@d�0��:���틚[��U%��E��ъ�����l#@��W:y�g�3}KzR�j�⌕L�^y���,���T����a[��˽Yv��8mYn������S����_���05f55.�27`���Fٰ��):�δ����5"�vwn�T��N�z�]��x�J�Dک����j+������FMۛV�8�n+�P��3�bc�V�.��f��B���Įԣ�A���n  y�sju�V�OB�$�.��f��w���=��)���-��6��k���j뫢B�Z�k)P�/%
h��˷�z�j%��S�\$KE����K��3�����5�6r�<�hul�����%�t!mJ1έw�{i��U���=̾z"����ʸf���-B�4�I���{kRY��X77�%8��Ho���L���w�`g�%��:�7�d�S��'��ޑf�p}�� ���hR�4�������K-�_r2ZE
��y+�9�I���"�ym/Fej�������zA���̮�ˑ��iW�ܳ�f�}Z�Q�*~9j���i���U�չC�ٵ�R�?�Q�F�R�w���]��LdK��3�]B7�MNO`���-�v��H�0K��f:ꔮ�����V�SŤmt���G�긺�&9S[V���L^h��-J���¢f^RʨL����L���
��j����}J�w�3z����[Y�/m>Z����Ħ����#�)�mf�ɷ� 1���{+mUz�y�>����w��㱪WT�r�e��;g]�?Dkw���-�|���oo�t�EO��&G�U��Pro+5Y�w��{{9T��ܺ3Az����E��n�
%��x�9[R��U���MHN��GvK�\k���E��䶝	?^�u?3����u����]�*�2���&������:k&rv
���{����j,f�MT�;�K5���+[7ﷰ�n����X�YZ�i7�n���8�k�M�����/�5�����Y+gA�X#y;ʁ�5W�
g,�R醺�ԣIէ���l�f�{^��~�����u �<ځ˕vp�Z7I4q�d��[��w�K�%^�����𮨮��S�:ɺ��^]��̕����Pֲ�գ*y�n9L>�T3�z�h4P���]�G�
ܨ�=�%u+�8z�b}ռ�b�wX�l����8�Tf�_!��	�����-E��:��T�s+��뺖M�-��2vȻk�,*Ĕ�Kj���L��>��K%�$�#���%��L����C3���q��:�z6��b���wAS�^��.�u�Q���(�x��q"�}۸z��t8��?;�o����x�W
��[Q���̫<�\j�����3tv��]^�9~Fg�h̺}M����P!߱Ѻn���;8e዆�"�{��;���:���#��n>͛bkU�fdjr��:�H�Ɯ$�	�xE�iVBN-���aۜ]�����p�$GCq�<���|w�3G7k H�\4)���Bh��,v>��o9۩�E"����	�Oъ�.�B�_�+e�:Αu�i+�d��/?v��Kw�s���F�f��vq�*8�yo���R�d�y�n��}�8���"���)�صL��*��,Y��#rcv���h�**��r����]
x�IT\����h���4ي�
I����F�p��[�b�:vV������yb��7-�I�#TUpP�ꛚ1�Z9��ዧ4���t@H��ʂ�����l���Ox_Rĩ!3�
�Oη��Gs�Q�s]�i�WC��o$��.L����x400o-x��b�f�h�mcޱ�<�s\��e��Ֆ�LƵ�6�y�H����`§[y3LRC��K�3�S��ُ�4c�Ѹ#��L?Y�[�*fUno�i'�k�t#���K=MkG�z��h"�I�opczPHj�OV1?6�tW}�_!�JwJ띪ٯFfv�Y$�����@�`�M��K��XRjN��t`ݼt��{9gn^��\H��3����D���t�f�g8����g�Y��t�PN�k���T]*E��k'j�|C��r��FNOF�]U�:��	�ٹ�j�w�j���G9�Y:�uH)�_	��D��ZԈS�@sgEr5>��3ֶǩ��L��-W����S#�w���_nt�K�ٳb�ٰ���醻CBcvP����&����Ns�U
�ܨ��QރN(34\��{�������NJ��(Gw����P��i�(ĭ��f�8��7�Q���B�����Ŏ�V���gV.W`�[�v����T�\غK)$�՝�*���"^������Sʢ��"�g~�qEsܢ�ݜ��G��х�u3�D�;l]M�Yu��Pޙ��2�K#�Ͳ�l�S�j�P[��x��=��o:#���'!�.�qV�Ux�
�e�t��1?�^��dβr��n��wz̫�Y5Kw,�DUX�� �k�ܹ�A|wG;S�J�(�w!+v�ͨ��<���2vdɱpX6.�Y��t�t�;�'��R�#Std�<�b����-�Rͷˇ&�1�ƻ��;}g��9E*�JZ�%�C���۽�A]���Ra[�ɹ6v]��k���'sx Ghef����L����g4��G���b�Sס� (��Y����p�O
�Wq!oU�BC�v�m|�оw��,�2K�e����H��E+؎Z�<c J���t����]J�:�Q���݋$�<�W1AZ8 �C]WF�WIL��xi�L��\����ѹڎ�|��pɪK�����K"�U���d��������#7Z����)\�b��m�8��oZ����ۥ;`6����v�3*l�,�
q�]J�-��]����6��I�>�6(A��c^��sw]*�bȈ�����C}��Hfm.`W`��o(՚���hf0�#�<�3�`��W�`����7 �f�+�j�;6fr��뻓g�g!���UJù0��;�+�<0��3*��3y�-��<Ӳ��H��­{���������j˅-gK�h��Y��:������Wj舺ni-1����
���J�&S��I�^c#u6/;p\�U|��:�us���Ĭ]̆Ϧ�6�PRt�K$��	^\�hf�ɱ��2���w{[�-���Z�t�09cN���-�yi�Qӷ��NYI,l$h�tn���b,�+�2���B��8@�8bZ*hR����鼠�)j��WA�4	��N�f6����ӛͭG�U3F��13y�R�wMB�j��fuh'L�ۜb&�����j�/�$�ɹ�kL��.��׋��jk��Φ9[{��}̍���M�K�;G^-Dݥbc��0j]4f*����.8���t��ub���h��e���xљk(/�枆�e�%���̛�!<�� a�G_a��D��!P�D�Z�lJbdd�jf�,�s�������in���K���a���2Q��0 �Kx0�=qU��)C�qѣ��7���Ca*D�ǧL�G��z����v��U��ҙ3s�L����]�M�;$^�
�vUSFh���[3^�N�v���8+#����ZRg�R��ʹ��kF�[P�udS0m�0�u���(�X酶��Xx��/��G��㇈{9҇7�
�l
�+A.u�m�����A�Sn&o,0r�v�I�p�]j��g"����ݜw�sw0ҵ�b�{8�٩�e
�l��8`.pO��
�$�38c�n�;zr� ��u�� 4��c�jk]�Ϝ��Ѧa}jC9\�U`<5�U��}�ȥ��s�]�p�9�ge��e��[qT��x���{^��kt���E:��f�v���0b��`�C7{�%�w&�۶��d�Y>B&�++̞ס�[XW.�**7.R�t����Y�yl�gk�%��Y�.�Xnt7��B�N���"!7X�T|�u�aT���9$�/��ؕ�����ӻ��il��,D,���X��
XX�3���f�w��<��V��-��P��YR�Ssr��ی���9)փQP�H>�h���h�`���w�����ux��v�������r�u�un®�H�P�Ý]m^��Wս��߇�̋��z��wT��k�T��ⓢ�~F���4Az �R�*�A��/V���
N��5�v���+6]kv�"��b�'���c;R�][֔�Ĩ4�:�B���5��{i5�8�ڳ0�_��(P+������?w���"� ��������(<`	��H��J�H�d#܀s(��T�:�x� ��p	̪�L��@L�rD^�r �(��^$;�ֱ$C=�CP��q � y#�4Pw+��2QMɨ�5R��� Ї̨jT���@���D�3�P8��C7���@�	��EwI�;��<��QޱrU7"g��P<�n�w��:�
Q)ܩ�Q�%3�H��5=���(JC8�9�9� %�O:��w���Aԡ�;�))w/>`�y���α7j$S$��P%#�=B��|�\�2N�8��Rf�|�
pr�C�+�`��&�C��S���H�8���0��;�܈u'����{�y�N�2 �W$22�\�%)�8�
�!K��J�)A�9 v@9(��#$�(T�� 7!�+���q��\��䡐���2^�S�@� d���>@��zWP!��q�� 8�� 8�2Nw&Ię)��<��q�8� ��:���	�9+�u�f�ܺ�܋�� 랴9	�J ԡ̾u��=AԵԚ��B�*���C�#@u(u'0�AO�#ԯ�b�.�
P�MC�d:�r��A�0E�9�)�Eܔ�T'�H����N�0S%`^����@�+u���:�w!��rS�3R'2��w	ǘ��y�s��=Ja�ɸ� g�Y�q��N!)S���M6��@��]ʗx	�#%M@d4��w/Q�Ԧ�z�|�����9�s��vJ���R�U�Z�!$@j �S�g7��"n5�����1S�z���c��0ZL����@�2A��pn��J@:�5&���2�09��P��)�c��� ��)V+�!N��hZMBd�I̚�Z�)N@�)��WP��Y���4w�8��/$%�q��u�R�D�[ݥ�C^b�o �/Y�����<�:��''���y�]Hu�{֍��ܼ����� �P�E�@�J]�*a^`�[�瘽Hu/RP�d7X���zѨ9��jL���q#���xF��m�V�
 �vb�@ny��$��)#2Y�JİRB�48��xй�
9��4&Z��9�(�P�iE�@)"D�����sހܜFAW��өB� �2��a7R	�%��FN�V(Y�eTI����2�i1���	!IE���Gp�9�Fa����`�h�*�7
(@�<1H�I2�j���P�\+#Ȉ�@BZB�+���l�8�s�kx�SֳrPn��x�:i*RzB�.ʖ$�(�椌��n8\,sZ�R�i0�M5OmY>R��P�𶞞������V'�yZ��1����K�`��Kǂ5��\�Bx���TŞ��!{ސY�8<�,=2�
���̥^k&%s�t\G�&��YZ�2�e[���J?�B⤴�ne�u��E	f�3-xd'z:�R���;3���������LAf5o|���ǫ��r�
i�|������(��v�WM:!1*s]=��VoN+'���+�NMͪ�4L�&�z�OI#)�9d�ŝKjf
i��bg��jڨ0$�$ØR��b��y!�;9��B�۽@T���+�%��,��^֥D�eކؚxD�Z�z�6o6�3UcX�rW\�.�� ���fnV�9*�ln��M\��z�{E�5�/Dd��t	w�+үgn D��T��2L��}5�R�U�[�0Tt4N���tw�1�b�-��!ǎ���<������^I����r.�^]��$A���Fӂ��� 0���L1HF�S{h��ꦌi_ "�*C�@k�.�U�y��+��g�X':*�C�u_2�س!+�q��t~{(��&����G���r8��hZ��APWHK��q*n���k��ɶ*�l�ә*�%o:�6�[�-eb�U�[��f���x��M��:�ݕ)N�U��w���=K4�~����rr�gu��	�B��nK �`'��d�UR��!	H����[rU���E�t���&:<�v��F��I��k�+�{�Gn����6]r�*\멜�:eU��c�Q�v�Nr�zń�m��%���Eb3�Yq-%t��1tZ�I��fM�7K�(��Nr�B��S�ޛ=�؜��B��_�u�4��B�$�q�{��ѷZ�q ��)7.��Ռem�Tթ�`�N�����V�R�oR�����Z�}�K��*)��J�[��L,r�2��[')R��[��Xa&��I+��T���ӛ[.Xkjnh�F9z�x2��Ki^�B������e;ԯ���z�9�+j�b��C�c���hk�P�r���kt^�R�X	dcf=���h:��h�c����A�s���������={�=���|���=��K^�N���eT�.�g^��o*�ԫjP��%�H��չP*gj�+�,��.��S��7������ �V>�3��}����e�i5f�N���畉�S�/q��0��2���V�o�˴w�ה$���;k:R����mLu|�H�gJ��9G�h��rm:M��`��ƨ���� D�v����;u�N��X{<=��[DT��!j�=�X�>64���i�o�<`��5�Yܽr�!��M�H؋5^U���,�sb�(x�ܸl��Xt�Hѳol��2��#pS��{G�-�vm��-�tW���`����5�wl�}F�$��E<���HWAEM�.��%an�Vi��u�x����T"WWH����NѦ�L�e��}�]���k'{AѲ��u���}D�"�������٤9��vc�C���k+[�SDU�/�I:��j��	rLY�V^-�Еd�엁E�*�<8�u*&�jf�𕗴l_\�
�կ{��es�[�[��)5��x�[Y!#Uf�ݩ�pc�浔�U�6��\�/J��"�"��b ��3�峬vn+S���3
��iVcП 29{ux�����L)bdՙs�Y�ȱ��"	�]�P�c�;Nca@�s�u�9g�iq��h�󺖹u��uc[��=x,�[k{2��@m��}W[y����1�c�c�g�w�f�[E��ܙu��Z���4���y1�[��gז~B�Q	(�vzg}���yskz��PZnQ������kU6�S��e�]T�/H�R��� '1Vةx��^���#�yo�a}H��/	ھ=7_U��:����s�k��<�M�(�8�S�9�F�^�D7(�4�ܨ�*�p"y+��ζ�� /ĩ�@x����2��s�!N`�9�z<�Ӣ$����wp�~�����;�)��|��  ( � $$��@��Hb@" �LB F�뚤B� �<�B� �  �P@!�T�$��DB�S
� B�� !$�(q� ��0 _4�@@ ���C��A@� � ��-i�@xhD �-�0 A $!#D�! �� �BC �
A @)���W Sb �   @�	x` H@%�� �H ����
 �	@! 2�(�@B�@ ��8"  �&� �� E��D�$��D!�` A �	$ !^�0�B� \����$ @$�@�ƙ
��>҅�'^���w}�6q�3+�FB B@�B	! B��B�� A ���p� �b! !�$�#�8��B ��y� @�B"9���B��� � �! Hl@S@� zf H� "0M B+X`5�DQ3�RP��R��	 @ 	��  HH@�z�Q�@�^mHHBnuv{4@��!  y�  ��޴�H@�,b*m A
 A�/����Iu�C�=�7��9  H� ��hU�Q@�B �?��!  B 6ԈB@@�� �h�K���͉��h�d� $ ̀!e�(��!X�	ZΕP!�pX�CM�X�4����s�i �Aqg��	�8H   BiI"B�8��N A�JR �c<4 DS�m6�DA !
�k����snu�u�7��}�j���1��B��\�c9�i�QD�FF��	]�饢�p !HB�e*A
F������RB! �Sa�0�ÈBA��8%x��I	 D��p� 	=)Ā ��   "߽qi�.	`�� �p/�>!�$	WY�}�-�a����M}:�۹r����"��8bD �f]l4qn" H5SR�h Q�����ۥ0A�d��B>/d}J��@Ȇ���8��˃�/X̂�^m�E@B^lD[Ul@���A�W[t/� !�D{g��ɺ`@�Bi̢��˞�*���������@u9B c����s�@@�	0Cp�!�=i1BA�����\� ��*��� �"G�>�� %����ƟV�P�BE�+�LQM��H� ��_T4A$Ĵh���-.��@ �i����[5���/m��s8�f�"@8�a )���f	�[p� @&!�0"��0" ��>����T�%�x��J`�xl|�}�` 	D�)z]@��&B{��f� L�(m�^p��A���,��_>��ԩﳃ��=�iB�M �x�$P��뵥!XЈ8<8�f� �����"�;-\G�m9i�*��K�������V��T�,�B ���@� D#�M$LG�e	dMJT -c��(h
��uا�W�;��WW�<p�@A_n{7�t����}*P \�>�ff��!� E�2$ !�.&a�p4AS ��[O����V	hR�0;�P-p��3��]��@�)@��n���[o
9ګh,SiQ.�Jܩ�����s�.�z��Ol� �����V�M<��bC:wh�w���=�N��])�o��������!�׆��Dd%蜘M���U^v�e�{u�w-�9=a~يڮv;*�5Iuu�}���� ��2�9줸V�L�5 zg�T�?50|�0� ?q��ؐy��{4@�Ɓbi��yMդ�>#���������Щ8p �˟��@$  �j�}�G޹�����b�{�2��4�{��!%���"�Դ��b|&��i��ȃ͑4�I��7OmZ)��a0B ����h !g�":\�0z��! �e}L@ P��*B|`� ��-����}>_.�_���������Be�9�!��94�i���W�QC��BSg}׍� ����P-m��hi���K��� ��дb'��|�P1�+���+ �7B��o�岶�c�nC�����v����$Q�_
�͠6u�Ҵx�$�����H�3'��X�!p��"@�pǮ�/��
ĸz��� 5s�]3$ ��*�"W���3͐ G���[WS��.Ϩ�W;�Ӄ��H9�y?Zd !0M'��_�0�_K���P%�99��ww����٭R���d���4�6�i���(��R(��O۫\",Lm�#�:��J�X�o�k�~���{w�l��8��(��w��	� 6NZ�S�,�ʻ�褀��>�����4�fL*(! �OI��R�}{J���͙�A8r�$_���k��uz��幛3(o�>�"a����XA��Ajj=�}I��}K��5
��D���$ ��_������"l�шm4_8�xt.�����je�m�	��JR^^oQ�Y>�ݼ����^4����>�R�f�.�!ͭ��m�����*�
GS,S�B���1 ��" �J�]إ]sS|�Z��chB@��j��Y
�\5#@ ��+Y�~����w��v�Զ�>�g�L_�%�=�Jb|&��Uy��]\��7a�B�v����A-�eȁH� �Hͣ�!ޮ��A�@��/eX(�>�����:�η���{�K\���)��)�8L��K�/�)�i�O��1�|'���y�-\� Q���u2�bA�ܻ�Ԃ#�۱JmB�3ھt�_4⧦��Ji}��w+h{��������B��p9����Tx~25d�q�s�ִ�ajD��:]	E�}�ҥqWWO9dq��G��+qP�S��>�~u"��3��	Re��v����Ž��RͽWG�9�i\�������D�p�&��������b�3U1"
i��d2D�}�����)!��b!��hаL ڟ!|Ґ^m�7.�/�� 9���ѫ�$"�� ���˻��i�6O��nX��^�{ӑ�@�i
<���Z` ��R�D�@w�~f}~�VT�>i��U�о��8��1Ǥ�HD�U�h�& D��D�t�@S[-?��۫|}s3�����;q߾���"c�z���pА���>��Bpc��جB.�O)�P�V�/��L�\�^��Q�c�I��RUl�@ Bwʾ$��e)"���u,��O%�޾���b	��Ѣ��:�QM=�WPۆ�]z���r�HoӢ���	��m�3zU @�u1�i�,r��/\,B#���Z_�+�{5ٸ+w�&e&D���uiL�j�\Q �}NQ���4�p
�Ⱦ��!'�`����G�;4���|�'��`ys�;垏�m��v����>̼ƅc<Y��@H��}w�\������!- �a	$�0I�]��X���C�Z;m���D��zS��v�����J}��r���~0b
vuX�o~/�5��j�*���!�;�B������*�7z�<�*ٮT��č�gU: HB��ۿKQ� �b��P� ^T�����a�D[^���`��l��X��+��v�jP�� _6|�=_y��`kVC�7��%��>U��9�q�]��x�c�t���Z�
ܖ�J߹|B*��V ���pA�g|Է�&w�V�,�j���dL�����v�di!���h��U�[h�3��!�k.{uN��o�ڗ1�X`���&�fy�����#�֍o�[��3�~h��i?jd��q��)`� �iHs�kΩ��/��`G��`޵���^�����u�X�m���7tq]�9�u�L:�݈wj`���ܥ!u)dnR���U3�bRr��hկyk-ٵ���1\���U��z�`�$�wjA�`.�u�wՖ9�ח�o�J̓*͔���)廢9��=Y�I�/�Z�y�����>jO�pɧ�2{)�"_�1`)�mNe]�����=��԰�ݩ"�Dq��B��B����8�J�}�Zԫ#�~�S��nwv'w�UJ\���Ӎ(pchB)z���*�袹�/������um�{2��r� C�>+�mtߨ�[��dk�~O�]�#R��~n��>&D&i��<0t� $��ƃd�u�γg�
8���;0�Xk8��bRҶ��
}�^,�Orj�dd�/���Z��eGv�z(t���r���U�6����ŵ[��c ��U AM���s �}��U��{�P���\%���$\���VH�l��ʿ��4��	�;,nhT9H������=��_8��&|ӻ߭X�5�����Q�NB�*Y�X�1�Ĳ)	�
�hD��'T2F�G=O՞ϯ��k�J��u}��6�YK�J�]�m6�M
����bPs[�=+j������5f=��^Sg�r%���%�C�^'.�7O�ꝼ��õ�}~%}�(}��B����_m;#��F����sV��1��@M����쩙�\L��!
�h���g�!�U�+������1�>����L�^�ڇ��\��u"j\?}T�B ���M
EZ�J����h� ��s^�d�E���=mtQ�j�5YC6�z�ǯ��$d�޹�Ks�EuT_��'�/L�,���
��R���E�,�c�aq��ß�N�t��B LR����fw���~���;��F
�-Y]Ց�m��U� ����->��N�4$��z�  ת�(@n�+*{�.:\t@,y�*� ��U�ʡa�h@N+}�&Z�d�l����ޯV��[b��%Nx�x��.e�(v��\��7y��7&pza@!�[
n�'X�%�1�):�=�1���*�P���*M�	�����6������*k���X����L�Hμ�dy���-������>�:6�qRgl���W�Q�!a��/�@�G�$��4[S\��j����]�����L�=L�̫�y�'S�rV��t�^�m�Ĥ	}ĿM/Y���qP#� .9�Dz���k3���s�}lٻzbמ�լ�X*c'u��ֶU�>����R�籺��R/>k�`O�r�J�5~��:���;x����_$�����Tj6v�֨1|���q`�4�o�D�A�����i������p+�3���zWk�6�F�-t!3$�T�.��+M@3$�H�A}X>,�楃>���JE���! ��\X�&���|6x�c�P$���/Bm��]xy\��m_��q#/�tc5껪}:��_��W�EkT),_~O+Ȓ{v����=���j��M* m�������D~�r_��-f�tGF��64�Ep�eg�e.�M\B�zҕM��_ŏ�]i�~kҳ��'T�Q�kU&�"��`���L�4cф����)�캬�Z*�ϖ
Kƪ�h�v���>�1�	��0�?Gΐc�#%��j���"�1���]�CY�Ed����L�:T-?�#��p����C0s��1��N}�6����]�i��\N}�G�J�����p$�ֲ�v~Ɂ0#������"�9����W�>ɐ�']k��x3�0�ʨm^��>g�8�ʭ��+*�ָ�a�emV۱l���¸b�J�T:�ZT�:�_;s��!��;i�ݼ�>�]S�c��}�؄����.���7�9mH��s	�L�R�mK���S��9B����&�R���Z^���R6
�OxY�GV��B��)�T_�>��!�H��W~u��
:��S�wuq��s<FH�'��pL�%P� HP�k��ǜf�ם���������=o��w�j�]H�0"�� ����&���kG2��&��ɫ��*=z=fi�tn��}u�]�#�	̇�=J� �	��Qľ�M��z���Q�XBZ(��-$�����OO_�s룸��Iʽ��wgd��ݺ�(�,n&�bs���^�	�Ԅ&�lۦ%]�����\����]�ԯ�xb KzY92�����U�$)��O�&�zbɍOX�LN[�}U����տ�ڳjRf]]'[3����F����Zr ��d�ji����D�	���An~�[2Gӷ�'��pIJE�Z%��*Ӈ�q�<l/����X�����n��W����h�ȧ8{�톾>��? 8�Lr�8@�`I?"ȲI�1��ڭaR�Mz�r����B�u&Z���_A�RV�w}���s_�V�)x��W��[k�?���zZ-4�ڦ:`��xF9#z���fa�0��t����>�a]b�7�������S��*m?\�ؕ}�m��� O׹�x����
���>�@�.���T�Z|�u*R�b��R`����W����.�w����)���he{�
5w��-HI�"~�Hʟ�g���܃���}�%������uiZڵ���m�R������.�I�MvC���_I�WX�q^>��QDEv��_
��z|����m5h�B�m���d��Şn�L�?Q���n����Y�yx@� De�(�u�y�'��/L4�W5��V�L�T�D���$<���1�NHt�P�i2��쫴��w��9�������2N�_sC�Z�mF��'�h]��H){(�����b�Is�b�����.5cq���5����@�9U��������7K^b�9�{�+�&�A��}4$��y�˓�J�6��6"��bf�/g(Z�w�7��f}8$SL��#`���C���;��f�ݖ���?0�B@�e�x/^cԀ�=��A=G���\h��{� Ԁs��g���{}s��	x��=��}��_�ކ_۰��=n"A딣��挿�v}��_c�	PԆ�R+�Q�/���n�k]��{�Z2�!Y�w����6�Y��w.D��OY�k�e ��Q�Bbj�3$��̲�w{,�g�a�VR�Vf�o�]h��זw&����8ξ�#���[I�X�5�}�1L��r��l+\�����&��]H!�M�7��߱.HG��ÏT�<��`p��o���"nO���抎a���w.�y��_&RB>��TG�b�������'��J�W"b#=��PP�qĪ@�1�%Pb��OmX��w4[pH\�|�~�Z=�\��\>S11C��eNP���g隙R��OJI�ۼ�Q�ޖ~�e����qd�g_T���y��):"��gw���\)�{T� B�~� Í}���r�,"�i�`��Ҩ4iUe���"[I�ID�vg������)�ЫmB��� 	�s��=�0�Fu35P#pf?�偍4�N�g���:�*cW��3C=7��n'I�FNӛ}k����cz����DY��ڑ5]2G�eA�h�"W���_���^���\�A��}udC�¡pL &�\ɋ=
�'
����nwի�����\���ۨg��ﶫCD�F�B�`�Ffʉ�<ޛ�%��fﭽ����*֘�!;�;(�8�jx��vN>O��XA1��
��['�)|E�ȣ_	4�և�)��Q�e�ޭ���{1�XҢ��[Bfb8e��)��]]�Nm|н��Od3<�$�\�ǟ������\H�+�z�|,�n
޶
�KT�#��l��>�_��mϟ�x�? ]�j~�Yn~����eB�v"-�z	��Ƿ��,D�5��+�Y�R__���ӵk�=� �����h����?��˼��8������I%�!3H�#�I��a	�x�B\Aɩ�<2c�*:�}���R���" q���[�P�s��nBQ�4����Γ�I����D(�N+�=�������8�����{z�J�믈TBTiG����Q�tu���4���4��P�"f~߾믴Ԉq��r�K�0]�WS�۶��hm�@��6��:� m�VTʽc�RYD�V�4�TM�q)�8�:�U+-)�i�n�w{*}��i�A�іg�̀��\j��JϚ�:�����b�cȳ�M���p�&��˺�("k�N�~�oJ�7�W3�g�q6�/5��zS�WWkA^�<)([�{,�IB�zmL�397���sd�HDJo�|��ݬ�J�q+����t�Ĵ!�y;_WϦբ�g��s���7�+ն�]�g�,��^�KƑa� ��W�(@a�x��f�q�c��G˯k����],�h��|TY4��r/�w;���(Q�f?52��,�@(Ϻ�<��eV���U�}�W�kU���zm���~�H��p��o¿���h�_��G{pE�K�֪g꘽j{6�uJ��q�`��9�J#�"B���UM�(���J9Y�x��%5�&3� ����H<-߬�so�S隀��Y��3*$Wm4D�s�11�T\�s<'�Enr��V�vW���;p�f��h�TT���\I�����A��0��*ɩt2�qS�-��|�j߉T6_vm�ފ~�Ak��]g?%��V�Q�8�����3 ߽����H���*���*p~�(V!x�T�%�M��>O�d�{��,�/n�'b���{��8�l���׮��ᑢ��Ё�I����Bt�
m7Y+\u���ʔ��>�.�}��uW�r��_w�3�~"���j��/c�I��m�����s��������(`��mO�j�w�vJv����(����C���^�ŗn4��R]�ö�s�������V�}O���KJ�ў���|M	ԝ��(�Y�:ڇ<����=;K�S��= '}��|��g_�m�믵�w�n���cԼ�ۑ3~�.�<D��eJ�WM�����G�����DcFj��J�ӀG����;u:�մ�{��S�3r���|N�����+���J�u��bZ?6_U����Cɘ/�Ő7[��B"���BF�9���?LD�t��Ǥ��@�"�Q�[ޙ����W�ߣ��{�|�x���C$AVy���ʜM^
�%{�_\��0�9�11S.N�1}�}b�u=�ǭ{,&+,v*ө����t) �=����T�~lt��D��&,F���t��=�K̯+q뼚�9��6��yF�v� b>U�l+��O��.Z�i�t�\���Җ)��Ӟ��`��zqO��洲�9�L<��'>��V�j'3�����^�qF:B7�K���y��X���@��߯��J�X)��Ss�[X%��i
�h�M陿t�^����Z��t�Ak7z�\8�v�1�O��A$C��5��j-V:�̙��
����m�ᢙ�ڏ��8���Q�/i6��O{�㓯���/{�[ޫ���}�n��(]/�R�m-s7�Th�׻f� 1L����R�U� /���J����UK�m<^�k�w��u؀B��u8��s�B�!l�B��+	$T�ʪ�>�xe�I*�j��p
`U^�É�eЏ�G���V�8*�N庋Լuo��4X������
F/
g=R����*���U2��)OK�h!�������"ϲ�R�p�����0wJp#}"2�ڲb��i�=Rl����Mh��qu��<�W�v"UU|�岫��OOJm�B���b�7�3d���򹗉�F��IZD�m�Dv$҂"��&@!�L�V]<�7�<]CF*;�y2�!��א�xtK���#�8�[bi8�K�!X/ł����ע#�Ο��)���L���_V	݋��W}b�ȫe^I��K�ї�x5Yt9��ӥ�����y�WH�S]�'��oz�>V��W;�ٔ)ܨX&zg*�y 1T;kUD�#��H� ��U��C\�^���{�d*��CNVMfy�&�m
���;W��+��F�|,��}�K��r3~��h��e�<-E�S���W���=���of���&k�0/*n������l8����P�"�ӧ�I�>����ߨ���R��9����Wb�\�K�G�����X�D��m��}u�k�"��L��ʕ�:^��w�����d�T�uB�������4EI 0�Q7��J)榲���ǌ�dڷ�E.,���u+ծ��M����Z1gz���ޔ�J�s"B6��w���W֌o�3�r��*�
V����[ϴ�����.�|Q���Ģ�L������s 
ET�R&�  �>�IV�wx3�"��L1���WӢ0D-��sW�D���DLGTY\l;�ul�����;>�Y�
@Y^�ױ� ��;�#��ۇ,0�E0����L��$�Ც�Z'o�_��-)П�;7��xO���tݠLu�ב6�)��&�����{�ݥDO�`�h���I�:鍴f6���JC��_?W�����,�R�%��S,�����#ؾ��u�����j��Cp&;z�Ã�?��aȱ�$�;��Z��*���R,}������������S�!ס�k��#/؇9�u�<��yBq�"rzn	(Fx7�ڼ-�j�r�V������&����^�Yצ,�˅	O��VX��w�=
�^���0�.�'J�����̾�������#�X������J���i�'G���`6�om����m4`T����9����9��B|�O�8�U���`A��7�|�P��Q��'#[x���|�:��͖��5J&��lȮ�E����u��j��9C�f�&Tc��^�x��b%����2<^jح�;�4.X�uP�=���";z��IOv�IV+��z��=�V����׵ǻ�AG���WQ�F�?��xy�����ǚ��vڹ�L�SF7�\��}����
��k�آ�u��(��K/�y؞�`����6�V�R�Ū�$�kP}���S���Y{��;ڳ�kt3Xc�ee;�Q<�$��Ň[�\�5��%�$~iV��2�k��]W��#}su����:�P����-��X
4.w6CR�yNė]��#y��eu�j��̊�fd�w�D�M��y����+��ᷯ��0G�84�a��i�(���*B#�B*���@嵐��2�b9n��ԓr�ͭ���7M��+f��fLɊ�u�D���	NӍ��fK�4�T��׳�d��6�j'04� 8�����d�z��}�qAّ�i3�,X�<jj�:�-��ַJ������Y�y�V�K������Ut:��ɺ�^n-ٴ�dLT�I0�M�
]��Cl�1u<ޚS��F�R��x�گW�� ,C�x]FJl�
<���єRRP��׺Z��+��;
.2��M�0� j���ye�\4t�K-��Ac9n�Hm.�ׯ�`�;��/�����93a1��3\Mh׆�̝�&��o�)m�W�x^����vfsC;�*I�@�k���E�ȯb�]�H�nJ�(ڹ �����&T���� E+
���g�x��Փ6X3b�YF�T������P��U����KD��F�;6��v.J�n�2�,Ή9�H/���L6b �̛�N\��p�+u��z�u㫹�!5B��5C5x( ٘&eS쵳)a�2��c��kuf+�H��;?kj�I�]mgT�u��y+�۴4Y�ےݬ��d�4�;��q�؞К2���zW>�a<��U�1nK�����"���br</Gf���v:�9-\*WX�fK�KI:�q`R�4:M�����Z��ݫ9:l�w���W.��'/z�����8Z�ܓt�dJS���M�@�ڮn�����ܱ��v���M��^�c�>Q	B��1��_=���Lץ��k�I��O���ڙ�YF��=�˺���ի"g0�j]Z�}�����60��؇u��iv��]̏�=3��yW����Ь��A���P~�R��dD���iצ�l&�"��aɞ��h~P�C}��K����U��;�B���[�gkw�^���E׹nHx%O��+u����yP"���>�&@F3���F5ю䵼�\L�j��-����f�!=B$ޯGFz�b3R~�Z�`!�ffC�OM��*n���� s�Τ�S���0s���˭�t<*���en	�W�+�p,�ʈ�0�����ڳ�ٞ��܂��>�f$��16����)�D��m����s�d+�vC^�^]0=�F��<�eB.Oҽ�G7{�,�䘻���߽=!����1�
C�VcX��>0������{���^"��6˺HϽ/�"qC���s9{�,�����J����3f�����[G�����Z}�����EŸځ�+� �� �L���QR�ϲ�0Ǜ���W�VT4�Z
&�.���!�}i
��:װ8�m`��P������3�&`����u�Q�7+� �ʁ)#a�H��)�t�v�7&Lh�&t���x^�ۤ�^�&��i�D�(���a���5�ʺ���9:EBg��H�|��w�ӫ3�w�Bܠ>횻�K�vL�g�vì.NG�=t8z�G$���&�*�nz���<Q��s��51����Q&���ڱqh�Qrҭ���=3]Xq\UY�ww]<�cj��N �^�z`DӘ�說�]�k�e����iwP��F)�c�9n	���4T9�&��p��f�le�mb��f�" �#|;�����b�3��#�De��Tq8W�G:�Tp�"��1�N��:�4p�T�[%�����	�{3\�P����X�WQeJ�A"YV7Jog;z�js[}�fm�#Dg;�v�!��\/T���X�M^,���I�^�L4�D�*�B��a �VE�����FG0c�v�wt(�d����	���;�F
OM�Dfs�䬁QN��G��������F"m0�2$з6�"	$�T)v�W��2E">�ݦ�\�{�i�<�
{����K�v�G1�cƍ��s�����A-#63B��IU&V�2�?$�bZu���H�|��9���^!����dU�A/n'KX��/*�c�ꉏ;ۛ�Д>J]K)ɓ�;���rV�9[�X騧%A�`)�{�+|a�F.{Y��P���|b�{�/0!��ͤF�(��h�.��<ao&��V9A
�~��ld,�*`��0P���Q��P}C�輌>�
P3^��q)yڇ^��R�{�6��A���0/�F�'�| ���?�gۛ�b a�6 �24Py2;ٸ!���ݺ� ��m���L���֓�k�2�=KJ0=b�3*�ފWB�r*��Jv����8�F^ԪLkjv�R��:����*��*�.T����W2�����2;�k�'�sI�S|{'�VL��4`�ו
(
#�eB��kd�p(���g*� {��}�T�tS9G��dҖB�`[�޻��^��)z���_��~C�+�G;A�� Ta��)�;�%mُ=CY(�Z��JJO�y&�3lƖۇ&	�I��u���n\[j��wc��Rw�k�埊�M�x�՟�˲��;���n�ւl��Ġ�;�)0������$�����ABL{Y�IT��+����UKĺ�Ӛ��
���X��u,R���E�8��uF�qk��k��]���oo�n��Κ*%Y�:�dz��Zf��"��(Ks�L�)�8�E���S}{zEMM�`F��ֆ�7�Ga��Q���,�>�M��冴�����Q��(��v��.���D��y��u��/�i+O�!�5��'��9a8�'�I7��##�J��������R~�_�iص"Hv"Æ����9 F�Ǚ��Y괺��-K�r	[Yx�E	�q3�1T�/�!�0���*���y/��4�+��JjX��+�"�fE���2��B�*����2��@�Z�?&��~�����,EU��r��0���at����238�r����fGŲf����F���\K��W�80GpO�5N&�T�����&b�+���=�8�ɉ �	=���4�[�mg��ٝ�X)�־�rab���*�����b/��`�t/!E�,�� @�a�G�Mo���gާH
a�{n*��| <���*�J=�v���QM;��4��3�(�1�yt�^�f��ćK|����_,͒!r�H`�9K7�*�&{<��E@�IR�#5m�VPK�%<��{>T���$7ó�����3^ܯ*Q�;81Ao���GlĈ�v�e�\H��➬��?n|�!��D|� .p,N��XG+L7H�{��0;���Z:����%��D�NB���.Ni��##�ѥ�牭R%�Jhm�qu@!�y�s�g=�v~�V�j���������U�̋:�8@�V��^�f3�m�VM]u9��R���y�8������� F�"�#ģ���N`ή��J&�g��ӻև���l��.� �m��\���ۚb9�V�V�!^�{��������D��[OE����ʢ���̮��l���+�2�nd��^yM{:i̿x��:�����#��6m`��H�p�����[�֭��o\g�TY�6W�
�i�T����B��_9��SQ����6���K��=62�\�7����Z5q����\��IT�We�C2�5s�)�{,�̜oKm�f!�w�b['z��2�e "x��Ųl�s����}#{p�Wv��"�=�yq���S�16�s��Ń۹��$h��\="oUeq���߼;�с�����b(�����`���n��b;�^)-L%�T��N���S/e��`��{	���\]r͔�;ݦ���p��dɖ�{<�}o�Q]�W����+��.U������-��9�\�]�/�6����)�£g��Ê3�]�U@�أO%�Y���*w�wM�*Nt�d�������/�%yJ?u0DM�X�74��;�2���,��^4:�w��OB ���`�̭Jd0bY>�5-�q�Q��g��3���T�0x� l���{�샑���d#D����R���Y�>�I���L�qB�+>�exb��K�Kj�W����/y����'�)�t�SR������)�}�ƃ���5�'�yGuVԈ*F:b��QВ&#�ra[�g�ʡ�ܱ�QP��P�W*�M\(�N��g��j��O�Ekm�0����dO�j>U>䔉�)i0e�Rbw�*u�����x@Q�2��D��o��C���S�m��M.�����;��ޝ�<�;\Ϥ����M��DC�����B�wp�f ]wʲ��<�3u����BEw��r(=�k�7ح]�&���wA��b���.f��Ӊ�� :�ֈ�����Hx5 ��	.�	ݳ�@���{,�R�aS����[ݷ6�X^R�r�&13jK��U*;��3n�In�ܷ?	�)֍��u���[�Fw]e��6�_���]�B뽍#v��G�rX�/��2��M��j�gyzvI�ʗ�p7�_^[jw����NV���:��ǅ��7
��]bqQ��}�A�69�������&�FuR1E��7V�	d��h�Qk:�z}��bU|�H��(4ܦ>��R���[�=��I��]�cY��p kG�(=�Tg�ٺ��Q����פn/`���3�{�rfaX�/!�N�ѓQ��P�PS�%�����`��U �����m��)m�~���0eL�lЏˈ�[�|�	�9�PJP�Z��݌��Fχ�ڷ"R�l��Ys��Y�ۇ�+��é`���kG�1"�����ty���uF�(ʌr��[�}#�6��
ʣVnɄ�W��H�TH�H�H����鯻�,�����S���}�;j$�D�YUdpJ^�ݒ  �3�&ҽ��/��;7BD٫�S=�Tm�䨐��V��1�^����g���7lh� ��~L�Ж�.���G����1��##�UѠ"��l�Q�HF�a0��'�8�����T{��UO7Xמ�h|C�S��8�{��Vb=���M����gx;�&:q �u�nF�1��U8�/�	B�Kv.e�%��dO��k���a�����^����ILA`Ǉ��b��(O���"g���fba:K���ۦ��:=�����229/�<�A�6�,+��~��+h���w�}ʉ�ˌ�7�!/�qn��|�.V䏔o��ic�R�S޵��|�;�~4m#�Lb�_���8I���7�l����r|�ٵ���.��@}0�o��@�"c�1�aPP#Ҏ�U���˹�;�"��}q�{�Ξ=��I��w��G�2R�z����փӻ�Mrj����ӵ����b�@;[� ٙ�����t�	�,b��WV��UM��b�W+x�	Y����z��h�{��&�c�D���\��n��I�wL�v8��\�ۛ�f`]BT7��4!��	��O_lX�+�ʩ���((o�萊[)pVb��\�h!"([4��O�<��EH����c�#��m�.:F%�����l�K��k�wĴ�Kޮ7B��'�_r���){�f�!ϔHw�_E�(�Q.�_��W�L�[:1	�e���
j�߰LդD�t��wA��g噭K�=&�zj_�$5�?+�Fb�b����!̫Nri	<���q]�՚ٔ���#����s��"�<���V�P'�N�aUi$�u�Y��i��Z�>�Q�`L��>�`[[R�nQ���[E�$z a��e-�"����T�u˝A�9���oB��K��W���4o��2I�c�pHVU�R5פl��0�";�)�HՀdo�!|��o�Um�e���=?>	/������}��  �$��e
��0V�1�*��u@U�7Q�~����!c���(l�en{�ҡ`Cq�痷U���b%J��	��J*�vrϜھ�Q��@�} {��C�V�72���Q0�R[��_M*nI�Q|�za�Z�f��vx�$��}k��4�H1��D�;���a�<�X�M�LJ���ib7Ԥ�P�����1��W�%y��w6^1]�]:�be�p;P(A&��i�S�捻Lt-�j�P�SAYy�s���v�#��d%� ����g�3��� ,���Y��.��1�&s*R�c�7�7+Lyy�H)��W�����A��@�����p��蘽f+�gm`��"NW��l��U��ą���j0	y����aߦQ"-���+)Pڂ���}H�\�f��T۱����:�S���X4�beTO��v%¶���ۉ�y�Ί��Pb�$�c(�vE��eZ��>��»b�(�4.��g���o9��ǽ�=�,B��n����-���r�<�� Y�I�	]|���[T�+���� ��(UG�nW�c%*nT<��cǭ߭�^���$ܗd��g���[<�� �F�̚<a{�)��^ؕ;!L�x`�P�*V��,A�p��|z�]-�jsKv��|s˗��̕#���ե��w�jf��z�����"ߡ��+摽e9ȝ�y}�D'$���\�#m{=�,��;h��AgY�6��7�I�ӕW�>��y�R>��[�b	��R"�BQ=A�$���B2�b|D:y��7����E�]��>GoqX����b�
�Y���r�z�г��l��QF��mg���]X߲�������sG���S���߇�B�i��X�f�.K±ź7V����+�M�I�����p��x�e��b��EI�S<��~4���,�Gxf%�B6~ԟ┘Jɉ)T{��L�����|y��2<a��Eᨥ�<�\2�/�Q�*��� �3�0�&��L�c�|j���\Μ]��%j��J���s���Q�n�D��T��Q�QQ-�d�� =��)�����4����`! @m��C�|̞u�q���{�c3��Q�M�)��V��<�V?U#A}�^!�l��C^;�a��I3��+�4���xm�"� ��g��QMY?!�':5򫧶��̬s�����MS�Q'{0 n�����{�~���WLv��i\Y���7IR]ˣQ�/*RpB)VE�UFU�Hʎ��vs7ϩ�¨� �;7�]�r�'���V���t:@Z��X�o6q[�pH�M��/2��+&�6hl�K�,G��
�,�V$�yl�bfl�(-z�'GJ�����hs ��E�nn��k�@��3Y������v����o�<��v��}�	���\\ڷyt���2���K%у�i6�fN��ua2=b�$r�ˬ�{@Ώ��	����V)�j��O�a=k\j�'�C��o�v�J�b7>�n��#<�����}[�� ���59��ݙ9w~�.J�	d�h+`g�{��^d�}�V&&��d�8Wu�P&�����^:�����)�T}�L��*.��ъ=�z��J��Ajnޟwml�]lȚSMC��A�K@�[���	���'�N���XJ�r#Ƕig^�R�d�[�6�����u9����f-��t�~ڨ��u�H�ja�T+�ck��8���2:����6�&s�,�s��/=�������Bjɝp_��B��C��r8��J4�T̜�^�5C�ILl��a�P^!c\z!gY�����Û�OB��Fy�*�}���R+���Z���1����S)W�.I���� ��{�>��K"��g���R>ؾQ����W��8Qu��J29u���r�i��^PТO�	�`����сu��/Ի���f�V���,�ށ��6��ϯ��nxD�d�
�1��\�LU yn��k�:v���WZ�;)m�ze���{�suX�Eֽ��CJ���_��0�1�Q�G���ƩUP�TFG���5s9��G��7Ʀ�.C��S�}�����_pw豕��_�\rnLkF��U�bV0c��f��^��g3o�4�Lڧ���S8�r��Y����z�QzC�s,_8CW]���*�����{�u�sUJm)7T�;*U�z�kc��)v�Z��|8v,˳#��>��/�i��·d˝F�W3�:�j�5b���Ai�.����%���W"A1�f����Q��^UL�<��@A7�3�zy/T�a���<��	,�4��Ej��4k2c���P�E9���@A������he��'����-��M�(,�Y�vs;pz��ue'�m"��"��G�
�`[_zsoև��DL��]bo��_
4[^T�J2�QT�@�ؚw�3��Қ�g�F=�R�j�Eu���?b�R3.���P-ӯʬ�{���X���jx���-ıb5k�v�}ѳG�ʍ�P�Y��"�R3�W�*h.n(a����+�QB&����J��+�j��o.U�r_�s��k��i;oLeay�8�yA}<�'�ʫ����Nhu�]Ⴧ�2�{���?��l k��LЀ�4�y�&�s�↸.�֗5�ނ'��ymG7�t\�S����(��M��g �w���$^��~��Ina׊�G8��g�%.}��VC�/z�<�7낇fԫ�&h�3��`�M�]0&���"�(��ؔ-"��4aeb��{�����-F"�0�E��3���A��ȣ�>�P�E��qW�hL����e|�-�߯ל�n�t���y~��+Mp��\�'�F��8�"��0��Σ�漙0���Lj����"�'��C���n�`M�r�\��b�4k�������J��Na{,���0��^
�Ni�a�l�}���}��*�����~��9�x֌y�c�[Fu*�a*ԕ7��f���x�+��sqW.gu�k�pÒ��o1�?+�-��2k<ս�-(���KUn6�ڰ�K�H���u�yAw�S�L����{n۠�A���`��7O�Kt�a�E}���V\�?vڸaB�vVh���__vx�4��'\j@B|���p%���u�q0<��ON�{[����l�
OU�^S�o䶽��Fa.��,���շ��y�����`�P�/�F�}u������$�]�Z��b���#nm]b6��T��&�&ip�5[l�u��h���	����������䍃L10�;�[��!��.�ZtV� �7ꬑ�=��ࢣ�w![�G���b��H�jf��M�}N·=�w���ь��8y��
��|!i@�o��(�.0��B�=a#�3�$��t�1�=�����zP1�	��$�s����e,����WO�H\ӘG���Y�Hux�]i�~���NTޛ�iz���Z�����֢�/�O�<ķ F��T<v��Q�N�A���3�C�[�sS��|'j<��z�����;>�`�-�S��,�=�~�[>Ƿ<_�Sq3c�
��d�a����b��u��*��&ZqC�2Pu�!�!���	W�ۑ?����������ZI|*����P(��q���WR:�=y=��gJxlנ�ۼ'7&�}�L�e9���WYٜ��C��Fme��yi��2%��.o��=xIrw��nc������܋�"�kn��tJK ]���aT8ʶ��X����u ks5�]-Q[�Q��왡��q,5�c䀗�e��#,p�à����B��!5���S�Mx�������!�N�e� �]���:�;E-�z'������vk�1ٞ�D�t6���ۙ�|����K�������=ۜ��l�$1Gv���T��Պ�T1Sj�ܭͽQ�]�)� �1X7rO�7�.T��pk�ژ����]Nf.]y�K�s����Q,�҇e��٤�������p�\o��V<s��K�֞�w[�M����:�a�Ӽk���7����^�:�Ӛǩ��N���\[SP���ҍB�4��P2����f�u��	ū��k��}T	A��V'ht�5s�]��/��ߓk�.R�)�dݭ�ǿ��x�ɫ�&d�u�&Z	Ӫ4����d�n�\� � ������26r7hՀ�)�j-k�P-nL�#����ks�z���,�G���%�k��ġv,�MSܙ�[��:��v�3�qjw��-��ST�ݒ-�O�����e���L�j]	�Ǯ�V�����+@�Xڶ�)%u��Z^wq4�yÔ-��5�P�yva�$U�ӢF�	
�B�Zh�]��tۓktrc5-��� ��꾬Vn�o-瑉t6N}|s�:��L,pv�7]�:������9�*�E0>J��C�@P�&vw��	A��2��@��]�(Wr��A6���@$���{�����WP�S"����m�3r�E�/[�9xnRء6��"i�:���l�
��J�S�5��l�*y�J�p0��=�(��l���p��m)��4�3����H�.Z�IaZt4�e��gP�}�}t�x�Y|��{���s�yS6Z&iZ�p�R�ʜő"Մ�&R�^�Y7�O*C؛����x�^�W�`q5-j�����Wu*�C/j"]�.c�TF��SM��TQn-���ކw!&kG2��V3|)
*�Y��B/��x��V_���9K3�_�����v�}-���A��َe�j���_yҷx�Ey�v�W4�g����rR��sY����!��w�(�\Ժ��igR��o�y*�^�2�)�:#�76�	�nJb�^[�x���C����]��Z���	�"7j��g3wf�e��6T&Sb���H"��ЧK�y7j�FK��kj��u��Gn�ʺQ�Ur�9`��Y�<�Z�a2^��V��f��6�0=�5�Ӹ���7+�ﻊ��CWn�o_N��\Ggta�&��*��h�;\��Z�]�����ͪ2�5���b�aE;�����(l�r���s
���J��J����6{jV\Y;�& �%�+/��b:u�wo��R]s����[|XX8W��3:.W�vs��^z[}Qޑ�t������B�+���'�>�GeVԔ��+��Ǘg�$���W��:Z��o'&w��!&��ܢ�=}��n�M��>Ws�S)���L���v�eU�.÷3&��ũ�nk�}�FȫTjf]R��P��f�P��ң6�S�t7��
a�ݪ��扳���(��"|����EO�E6�����2���B����	-r'�����"*2-fe�V�n�Fd�h������j�Q�G�/�C���O&��P�LM(���"	�\l���	>���W��˾�@B�&�(�W��"=�BI�YWƱ,4//L �p)��a��R�\����Ͻ6Э�貥Ո�Mr�M�1W
��1�j�<_,�y��nt����y����_�R�+����Dâ��%5�^�9#=8bw�K��W��s8|��;�,MU�3� �{�}�·-�zw۟OvxD�l�p�"0z	��m�]v�J��4W�י���2�dľW<wGT��J���Վ�zv���J��89�;�WV;��t�� �!@�f;v�,�Dǥ�F'���r1)�ET5g��p_�Q���@]c�W��Q&VG�ޭ��+ޖd�Uۡ�=)�M�,t1�	M�*<��+n�afȘR�z�>=90��R��d�<�=��꺒r=�-�7���{�!>B��ʢ�����*�����Q$���xl��m/YRo=U�Ҏ���
̟|mS����r�xaa��Z�#�O;WPOHѺ�}��5�T�%�b��{7��_�a��~0s��\,@���I������j[�ȱJb�Ìs�ȸ�B2�!�7{�&U:��`�t�7Z���Ŏ��V̓6�IH�e�m�ɡ%ꎯ�6w	Ԏ��h�t�d�iܽ5�,�.ֵR��;����b�e��x�]f��vV1RE݃��ţ�dJ�6�);�9#<o'ێ<ňnG1cK~���ߵ=pj�T����}���U\��t�^e���½�,��"���� f�o}�#�*��!6��\�Q)!w�y�y_ܞ?N�y��i���t�Tޮ"�c`C��d�gy�2B>b�D.�l�}��E����T"��E�w���7B��Q�w�t�;p���$��ʍ��7\B��f�rh�u���)�����93V6�J)Y��WzpJy"�L�.d�:�W{���/=���>�ih�Dl��ٍ�f{s-̌��Wƙ�v���A�
\U��+�|��Y�=�w0I�xV~K�jm��(���6T����)��$���;�T8��{f�c�%���>���Y����N��]h={�o�.G��3�/y�T2&�0�Ӂ���x��D��-u�9�ά�e$1R�{s�=��#�H����h��G��Q�m_*���O��T
�1N�e��'�(�w=��]84'�[^��q�_����;g����~�7J.=kvZ�f�RN��	C�}���H*�m���.�o����I[�3�*l���E�͌:�@���u��j�#��8�����ɘ����C��og�9��q�E۷��A��;�Q���q�:�ʇ��7	OL:QY��XW�^|;�SI��d��kw7��,TRl1�0�ȩ��tUa���f8�M�q��R��fVy����Eԃ�+	Q�iҡnT���(f�ĵ����E�{�~�BN1�.�@���8赹�עk�� u��c6��A(�����1(�^�J��fފG�~�\Ϋ}Nn�e���9�Vu���&4@����TLQ���+��C�,h7�S�~�Z���
4�߲��߮��{S���ؔ��	�8�r�� �pڸC�n�3��>�0�6�D��˼~�~�^j��ܘ�BgT���s"��͎��T���ˇ�,q�)��M����y������9�G�<N�\W��3.<�-A,��*u���'�u�j�S�}�`��sl��!�ڇպ�dZ� ��Fu�س��{8ʺ���:��g;lǞ�����J��� ��	q��H�i����c�9��ޙ7^0�!aܿMZt�;���I���~ZoN��|�9DV�+���G(1�8hYr�I~���9�Ug׆l�R.��H�^]};�E���+�l�W�p��sK��@A�yxϮ��EWB�x�y�Q~�Ό�M3~�0����o������G��ѧ����H���y��;NOh���p��G�O����yir�������X�L)=k#z�$@�Q��.��F���?�}�Ե
����!�!z%�B��(�3\1U�9΄�`��`��%�΄ �ǲh{7ӕ����[87]��/�[�Q��s<����UR�����+�엎ps�ovu;�t�fє7V�nQM�S'Q�C+��Oq���H�o"ԷRqn\�ed�i|�U�I]�Ά$�a��v�W[��XTs�[�R��/YAiTuG*ʸb�q7�@WD�ޛ��}��������'����Uv���y�W�q5����f�?p
��'�xz���=�;��,O��m�Kו*���c�|>S& ��g�O��UϏ��>7�iN�U�s��?'3��:�������ǔe�
�f2SX�+/~��gbT!��=�n$���ϻ��_�u�ۻ/@���ˎ����kΰj��>��:��4��n<Ѭ(�F&�g���� �]�>�ǩ���U��gxʹr#4{ü.��/�ى���ө��c����e�c`
/}>\�4"�� �Udۢ"���-H9"�A�N5�Ķ��z3�f�+ܝ��Ǩ�q���e�B"p������{z����Co6ו�B�D����E^�b_�7@���UA�u���=j�9^���,�1d�tLFP�K\ʙ��T��D�|P���� �;��p
�DPM���LX��?zZ�����U�+��^��W��/
��ٱ���t��G���;�5q2f�{��}���ʸ&���ND��P��f�=� �����ݟ^��Gt�_��xT��(^1�Q�L`�;)�A����{�2ٓ�^�}���u@�%�꠩訝0����I��&~��F^G5�ԩ�HU��7wB����L���D��H�N�7+)��x^w3;�WQ�8�yq'�$���u\�[��U�q��A�6q���d�6-���e�:uXaQa~M {�c�4X"g��Jj��2�}�E���p#����0j�2,6���L5�nw���/# f�I-�t5�Qm�r���M��-�	������7)4ԯB����J%�UD%Qs㹹|k9R�^����̪���� \)=j�<RH����z�ko��r>�~ާ���k�>W��<ep�������GgP�vI�7W�e���x�ۺw���ĎPR�q���g�ݮ���&�{�-��"����<�J��-�*�Y!��Y����:����.���f�@�H~�����S�4��s�I���?jBT�?`�G�G[�������_fo��:��,�淎.`R��ğP�0q�ch�;v��X�xd��x��y[dP5�|`��{^~iM�U� |���Vǵ�b�~��«���eu��+U�똁��� ��|�u�؞�j�7YV��>�{F�n���b�z��8�LM`W|��w�}cϤ�o(V�aK_NE�q��p�>o7����<���W���Z7Hm��"Oi�eyZQY�g�u	=�M^�����%�J|T,z6����U��WI�-`����o��M\7OM������+1���Þ�u�V���G��M�O�8��5���|�5sb�?�n�5^
��uQ��"��l��I��S{�%�p����*7�}Q�u�03���^�� {.��S����2Г������t�`�5��������kq�Ƿ�j�,��ؘ�t��0�]Y�?��2�IJ�{K�f� �fU��]b�Ԧ��R�^Ӓ��]���}�+j���~�r�V�B�-�	��ܗK�U�ڏ����|�d�<M�{�W~z���/�v�B��kL.�pn=V��]++o�H��u�3��������OÍ�i�����������nB+ŧ�����G�;�E�(KU��:��<�_�``�%o��K=w�U�L�冢�wl��Aɑ����.��b[0���a�=�����)�����;f�/��c����'��Q[��ƛ���{�{� Q�D�U�CK��D�T��*�8��Bɭ�0���"c�b�wO3G�
��>pEz�*��5_ņ���]���W�?[ɴ�l�O����gs�j�����"a�πY�p˼.Է�=� ߸�S����ť��\���yUy7����V�`k>�jr�<����b��rgfq�i���<rj���0�������;�F�Q5fb�
�e��)����-�V�y��1I��E�F��ZMز�.�f	ʊ~Q�6x.L˲��Z�,Ltj�����Z�����p߳Mq�]>�<�~݊�q��ԥ
����) >���K�TB�t��I�鼘�Q�#)�jN��r�\'��	���f��\�dϟ��Mޣu��g��Cc����l���,�T�/Lx/�Ұ�ʋߜ_��iE�<~q���g�|��mG���q
��p���Ū:���;)�Wn�AGz�ޏ4c�!�S.���ڲ��%��@�����Ω��h�t�aT'��oD���i�ݱ�x��9�so*�D���k��j�2��7�s_,��_D�����������V%f>�{�0�{��À{���� ���!���Q��fGY���n�9��ǒ��{��}��kLWݷ����N(��H<afM�P_R=8Lo���#�sxs��3�d� �mRh���s>UY��هY6jl^v{0���D�{]TP�<���TW���dU��g.xE�1���/�w���o���o�)]޸��hH0F8Q�{���o�W�,�UT]"=�*�},N+�>�c��iE}�q���}�y��X��L-�k�'1�t� =���Q١>��i�Ƈ�fN�F c}�0C�zR��;��F�]E�*��˪��^':�7L��Pa|y��p�S;Ǣ�6�Vs�(� �E�9Dv}�%��duz8�y}⦶8P̃ڂ��[�T+����n��FF%�5Y��+M�P�D^k�;U}쌨0�h���qpFr��{%�MѴ�oÝD��+r_���%5>�Q�V�l>!��"#��*s�e�TZ��XT��M�1Bw���o�;p�j�=9X�.��G{�s�pѵ�3�*���nQ�C�,	��M��_mZ�z�wLi���m �	��kəR1��,�֮�Q��{�	ف�w5�
�r��h��|�O̬](ǱH�^�gB���`��(l�6�&�k�b�v�,��i?���ǒ�rL�6j��۶f�4rd:�F#Ix��Ad�E�i����B�}B�!d�Uu�*��v3(�n�27�?D�R��*^:y����.��d����c�X�`%Ȭ����UGb��S�d{8E}�����r�;O��z'�J���z��&����v+�k���7�Z/���Gey���b�f�G��ʶŧ�s*A���*L9�Q��2wl.ٽLu�z'�o����e��;�2�m�6c/�.9����U��wVq�SS�3���pB�C�pZYiyԣ����H����OH��&:r0�P����9�*�^5�F'�5����\d��/4I���C6]b=�v|�w"�=�J��/9����!��D���G�j�aы�<�
0��1�Q�;�v���쎩Û�*�F9WN��m:�"�oy)�'�Ȉ
Z�z��������g*>Rzr�
�P�\򽆷2.1(�]�s�_b�ga�s�҆O���ga���g�h�eI^ت�_�Ȋ��:����\a~];յ���Y�s���G��T��/f���3Md�5C�P��ra�C$n��몢:8 ��f\K�S`��]5FFy�������0+=���=�Oy/z%�9���%]���͌�B<�^x�s���L�6����O*�u)ݾ���Vٿ��z�Ђ�E���I�a�wX���qN��d���\6�x$�5��:��po�w�c[f+����5:x(�E�����Zzؓ ފG�����n�z}�"R���Q��ܽ�evVs2z�mm:ȡ�0좴���˳/LV6����2�ُ�~ΜU���n�] }R�א��Q�`u֫I����Bj1�U����p��M^u3U�w��u�sꝙ��}J��%��עgB��P���u+Ez��2]z��q��{樠�p7WX�٨6�	��'<��S���5Ҕu 񠟥D��:���}.`�`%��c�W(�'8��U�Z�*�#��2�����Y�����ڗ�-gn7d'�,��?�%"���{��.�>�44��jSA�bA������k�7�^����{��n[�u(��)����˞�żG�b����s����q��d��=]p�{y�E�FI�r0+;��G;�	����ֽ (�n`�Z^0���p_2�#}Y~N��~�#�;�UZ�ն���>���U�)I��?P��2�AN�B�y>#o���d5��b�^��5k:h�G����De�L�H��=^��Ί4bB��p�k���:��L�+�1��
I��x������}	�����3����"��y1Y�Pj��S}4�nڤTS�����3�~�x�'7�wb��x�λ��j�J�Z���k��?f�^�"tH�B_�� �y9y����K��L/�w�Ui�;q��n�άs��R-�,5��42$�u_^T����ܭ�jl1�,��+w����h=H���sT���y�Փ��W�er��®�!����]��t?���녙uh�pr�Ԯ�I�7kf�
CB��l_J��j��䬹0t]K�2V���&�Z��ۑ Fl��;t�#Wx��N�B�K5�����q��ĳ�-R�?�_����p{b�Y�9]�O����B�GQ�w����5`;���S�AR������w�"�E���@�^�5��⟳wO�I�{m���Wz<V����u�@:i`Ϗ�f?Jr���@�b{*FOe[�c�*n{ف�l�ë�6��3��j��@F3	y	��N��g7}	��i�R�����wJkνK�Ѱ��YUp�9�%16{g�՟{@�<#��u��8��Jb�K�W.�r;S )wZ䵾�����O��/u���Q��R�Ɣ��nM�U�}*u�u�9�DuCu��w*��=�gx+�[��������ۖ�[QOf��X�이�E��oyr���sz�Ղ�>�{X����D����뛙���s��t:�n��2,�HVP�N�˖~�'�/�����_{�m{�v::�FzzCX�j�Q�#��u�}r�¢�`�M�1u��	�wA����V�<'ϓ�j��o��ѹʈ��ڒ���z��_X:/�{�3=��W�c:�IAP�e�Ub�����j�w��n�u��5}hk��@2�gu2�ר˥�]ɕx37��''tu�����>y�5{�$��Ҫ���e TM$���5I]l9�M�8E���m�����)#��ݬV��N㤮w����y-_W�0��c�vN�6f��s!AY��%BL�=�a��[I�����/a@�C��s��X��n���ĺ;4�q��1�b=ٖtE�!��3�M] j�#E�t,
���M]�8p�`�Qs`����xݼ�I�I�-;H��WW70H��l,�g*w�:IqPL�K�T�A+����9Z�,�u��=�u�q7����Z���,��1L��~���J�aq��������ά]r�y\�79VV���2�S7�;nuY���E�����X%(�,�����U���n�ؙ�%iD��*ΈxL��]\#(��mN37��7���[s}[ֵ��D����s�q���w��b��D�O/,�w����uj�b���}�7��d:SXk,~"m�h5t� s쮏P�yʯo/��V�MaB��.���Gg���a^݌Ӕ�Hڱ��r����x��(��{���q꾭С���kw@��.ݲ�	PI�]1�t�Ey��VhM�Ӱ�i�ubȣujI��1���.�щ�����Vl�Ï#f�M=�Wo�85��u��C�������%gh4S��e;��fL��*�t��gW �%�%��js2����)�Ϊ���U�"4��X�/D܅:ڕ$�7�q�#���<���\���-�f�q:�N������ 	����{"����^��)F��5@`Bl���k���Z��bG"�h��[��-^)��J��yB����g�wid0�҉��`�0� �]�ovd~�@}9K�t�oB�gM-��	ÉCzX͘ó�T;X��/^�v���;L��?>p�Νre��Bo6ġVVA`�Y�s�y;F��_�fd�j)�2so�]Õ�L$�%�R�����Cᩛ��V���x��U�,��_F�E�\�-	��tG�R�Ry5�L�Y®�����+�E��&S]�S��[���4iٕ��x�EgR�@�D%>�e�B��,}S0o%Aۭ2�k��U9L~L`�C���mҦ�72wO��O���T��E��wq*�X�"������^��D񌞏o�D|�Q���l����bFn�[4�GX�0@+F�W,��&��^�jf�y2W���*���Aqsc�*����'X�y�N��TS7b5Ť�u:+n�"��A݈��L#7vu�Y��A�n�=!�^p�[�=�J�j�Q�D�[�H�v���ӻ4ѕн��4�;}�Y7�c�(��t�tn/�I�Ӹ�>2hh��F ���!�h�xT�jQ�~�XJ�B;���+���������d������&E^�\�GtV.Fު�v��RLl�hw]�>�,vegeus�6��h�Av�wfYЄ�P+$�'>Dq0'c�TaYƍ?�}�D}�xt���5��q*�y���i�$ȿw75S��.�+�oD���+Vnܜ�A�Xf�^6�fQ2
*�2�n[�Yx^��G��U��d�''�S�Υ���}��Hζ��EE�.J��=�b����O83�i]�\'�����Ϸ(�g[�;E��u��|=QAɊ1ǂ�$��������ש�+����7)�Lf�������.�x��+26��%-�9�1ΧX�n�V��}�^���K�Z��e��C��g^9��t���X�i����ya�y���2��/z:�MGf��J�p8X��b��/��<jK��"����m�e�9�u/<U����f���H1�0�N~�`뱓�Y+X��k4k��GB^˳~>+ᚒ�Q~Q���X�i�J���4�:�_{�a�Z�f��ɝ�Mԃ�r�U�j曘@/u�B�����gmf���񖵾:�T��/!��Pnю8�D�T��*�|�=_N�K���2�J��`�c���P����^�f���i�g�Uz2e��JMj�ݵ81��^��<��y��@��7?hdx�<�|�!Q��>CB�U���7�[*'��ox�mB$z���F�Z�Y>�l_y+��I'���`�5��7��,>|8���@f�7Ǚ\����K��}�i�ع᫢�.WұX�{f��ڏ`��5CI+!��ot`�^�Z�ٳ�� 6o��7��J���/9EqVV�d���s#]	�9�xYށ*�b(v����k��y+�����
�ѭ8�c���T�!1�~�e�8��t�gN8��7��5N�?<^*��8�m���P"�z��=Y�7=N�0<�}��ӫ���.�
7]M_��#��B�]�"=Y�D�m��J����9���)⨯BLO±����]�����g���ͫ�5�=�'&���D��6��ڄ���!�t*}���J2Zw��?	�+�lgyH���%z%Wb;G%@�(�v�:�s߇���tj���sB׎c�ps�z��FF�P�μ�h���9t�#
k�񇡝�ĝ�s�Vx������J����qC�/@uv�>�}t<�a��n�^!A� �߶z�B�Q�k�o�$���$'�с<>ChhI�+���*۞�Tz�u���s|(
$�����n�a�{9���^�G�+����wvM_�n�L_�4X���8AFx�{�����]׈k��Q>����s�s��u๻p�n
��
2Txм<Fc�{ /KG�*�砕��R$�R7�5Mqs�=�������A�"v'u�"��֨�w����1vc��|�OCr������g|��@�;,B��ؖ�k��Q,��ƍ��k������]�}`+Ó�KZu+G���<�C:�ՍY{���.�/��;�m=J(h.�ծ���:{t j����n�й�[m���`wP<Sm�L#�v�{��ݦ�[�I�������^��&xrY�S��,�؏]8�C0�.�*ZM
ލ,U��A]D<Ŋ% ��[�Cr=#�cN)&t���
���Y3�\����aQy��T��&����W��PSC�~~Y��3��ɤ�� `5 I�nmL�1'j��N7u�|��5��=��b�%�|��'��;0{,ӊ牷v*=���;���q�`��O(��M�,�l��%���r���3 ���lfI��<�5�~6:�z��}|Ι��J��'/c�N����p`#�����Ճs ��#4�D�/���A�:����9p���,;C�k�o��}G��_\�J�}0"�pmD��������U�eL��u�����۟�3_-��Y�r]p��^�}��x�|{6Toj�s=�J�ޣ�o�Wˑ�j�I��+a�K�~�%�!H$ %uYiq�w�v ���Ɏ���(U�C��>:��F8u��1�Ϭ��O�WajXY�%�Ĵ�+�����a���`�%g^��zJ����zo5X���V���1�+�@�q�!y{!��y�h�b�~��[����ڙ.z����s�m�+uu>(�p����QY1ԯ��6N^	����7��T��x�A�\��dZ�_W��q���co9�NdE^=8m���2�8�mvYG�#����{W%�"��+xd��VvsY�Rb�l�߮�b �Syf5�uK�lf�gsYo�S�`tiT�p�m�&�v\�{X]����P������\�C��HG�N���xOn��W�Q�Ŋ�Β_>g�;�u�{@���t��h��v�.�i-�xae@�]ڂK���s��{�5�$?
���D'�c�s��-����펜��.�<W�گs��ؙ��\�>M[]�8�U��?�֡.�|�3SE)ҷ��}R�3�l�똉rS�Zÿ}�a���(�N�����}�%;W8�< 쨛�������S�\�8����&Q���Gٞ�w��]a��ҙ��i��OS8����9� r�C�̫�յ�!�R�=]K�@��u > ��H�
!��G���V��9���7��oDs���aD\i�V���>�y'��?��5���sQ!_y.^xⴰER���ɞ,�ݏ2�w��8j����ꊱ�Y.V��������,jw
���J%֩>k+/�i�á���6R�'����+��8k:���!����י(��>��(H��P����d��UKՎ}g&��tB���1����,���+s?>����B(#�P��Vז�1M��q~��//{��*�ʚ�f��ϖ�Jp�P��{��h������	A 9-�2�Go��z�D�9������y�l���Ul�'�oMa�� ��Zk!�*��ኜ5�'u���<��P����\Jl=�����g���}o�i���������n�<yF7 ��vD��gCj+6�,�9��&Rs#��;��Vf� �S6�f`��v[Ƿ��0\����vג��fPk2��P��d� -�����5.o��K�?e�s��'Ӄg
�y��R�71q3yV�)^Y[��Л�P��wg�H�� �ŧrb�k��=�珣��t�&�1�pz��=����5��4UK�c��+[�[�W��>���S��)�b3��kT�2.�j2�a��qR��@�/wn�f��d9�Bm�bL��Enܽ=y4hӘ��u��r���z	������ي�T/=�3�v�cnWI|�h�Zx��B6&��R�KXWi� �-��=�UĞ��qX*����]��kL��
���^��]��)v+;]쐽��ԅL�����cj)@����L���R�!T��z�V�� �M��`��0�E���j���G��4����A�W����6 I),��G��F!���������F����ۑԤ��2mf�����Pq��q��L�g׎���J^�r�{�!��{�P�nZ�_��^~��2�<|���JwT5�q�h��v��}�M�	�� �Yy��6���S���38��[��s���������*B�T��W��E_����;�2�(vC���O�������6�Xn���`���e����C���%�'v�c��m��B�	�;��K�l�v_aM,��YV��s�{R��(����P	�Ɔu��EN�Ö�<�r8���qU���j�����Oz�gs�wۗ	f~X�W/E�s�T��c�Db��3�Ъ�<wV˫[d+�X�W�K���������*Dh�e��RU`���R��aV	>1��/�R1�y� ���ڻ��}qH�<n+��;Ӑ5�ʣX�Σb�ߧg�_fbd��Q�������ȉ1��Ҋ�˵��<⧸̠}~�aϡ�{�אkaW����!�F���G^�~���tv��+�ax�[�|��q�6w����w�����Ղ:Ȭ^>jfU��SH_6��Ɇ��b>zS{�Nf�"����T�J���Q2��au&�ͤ�.3�v1wm������|K���Ǧ�ؿ^��֋�F��p��ڋS��>rc�B�w�����~U]F�b����˶�e�nh2=��]=�	���ơ�:'s[qw�(+�{Īx��/)�(fED�)K�9H@9jh�����F���y�5	Q�[��y�'�_��>����/:�n܂S����`"s�˘���c�w���Yzr��)[%��b�b����$A�:���_<��gWd{�+����#i`�qH����7���i��4�9ftA0%�L;�e�R#�I)+���U�K�ZG<���z��Jݨ��yW}�O7��F�j�BHGi;���⣻�A�׬��}8'Y �l�ҏ%6r��_��P����
��݇k
B�I�%��L���A&��F�4��ѧ���
�oD��f��7�����/{��	���ꇇ����������x��"���~��x�J�>�z`>�ł�*���&m�l��I�7S�k�á�D��|�#����{�(�Aڄ�:��}�baT��X:F;ŝ�t��ME�=0a	�Oe��Û�@	#D[�/��5=�#�����=�z�� ��v9�����*��74�ʬ�xv���Y�&3zkƲ((�Q�]m�H���F�tz�Z�u��B]P�tD�kw�SGx���T:��^]� ��=��>oR���%y!�"W;��L�  �@��e�G��ѣ���ar��.�F�4��,�`��}�'zM�������c��|�'8����q�N�z�x~*�`K��ҼC���ϔ�cs�D�r=�d+�J=qnߝ��Lj�)�V��ޅFʰ��*�:m^�^�ȩ}W�g���]][C Z��uȅuz/s�9�ێ�5-�������=	�j�����5��W'MTR��s�8�k��0��՞��ٜ숹P��N�p��Aﺷ���-�Iݸ_tcvG���Z�z=W��+�h��g��0��*l�Ⱥr���|�]�׮��Y�!��h�������U.��,�uo>�;���*H#��1����b��D�F�LJ ��LS�/"����s3�u���У���
xG�RN��vC���aۖj+5O�k�(0��1|.j�X��.��}�җP��>�d+Z�B~��qCO��5�>���f��ă��6��/}�L[�6�.��FIL���o;�G�۪m��T��J21���R��;[��*k�{],Ăbh��Z�)T8�k�x����a�RCۨs��@J;�����&<{�l�nn쭓O�B����p�ފ�@� ��M
S����?Vxբ��w˲r����bTxt<�}�N���*7�Ͻ{4b�ʊ�W�x��'9�T�<U�(eMc�4>u��ν����z��A�Ag	Z�z��~+k�j�����,;=N��>$��S�\z��,�PJ��=~��.5�y!dh�&o�K3F��J�80ߨr���j�[���ֽ�vz���ҌAc5*oy+�z�O�Y��S��\V�*����0Q��:�/� DTN��^P1���4�N~iE��Oc�7&���ҹ����#rZ�;���7��T�0����l�KSt��Jόn�}���O\n���A"�c�y��~��ҕ�
s_���Ԉ���;�a�r}��T3E�
�	'�5B�&�w� ��[]�=��.��o���r.�b���##͗��2Q#c7!TkB�{n�Ѯaf�:��=�)�0d�'��7[�g�8��a���q����tu�u&w����'X�ǈ�4�D�yB�6��◂T�|��5jT��i�!��Yt��d�AV}�q�C�tq4s\��ܺ��j�/|�����w�(�u&�Dv��yC�1*�90bv�r�zy�Onm�-�#�x_�)���\ǹ��<|+�L�>�E�f����q0Fl�s3��NWe�������Ig��dG�_��L�¾Na�gӇ6%z{$�C3\9�t��R�d��o����[�$m|�D��8�B��;{b�A�^G�j�Fĸ�	�?Z��dQ��Y��aq�������L�S���pH9�Tį�z���ƶ}��v�e�8[�}c�+k{�N�1��O�R��:=��r�3�$��`ZӚiw�v{S�f3/����^�����J}��uMR�6[��#��[]=WkV[s��~���=^��,�{MP�6���TI?W+�#W��ö1H�zP#�����(>��#�ǽ�(�P�p�ʅ�X�-��'��.�[E��53Wy1H��^�TK�J?4B~��>�$�	>e��^��2 �Z.ƅb_���3�u9�����ȗodI�߼��K�g��]��)�YU�:���z!f@nLK�=���Z���c|{�(h�z�?;0s�QaÜ�?gq��V_�[�F+�S9�1�|�r�b�n���V@�$�Y�*�~62���X�3\�"�´ҩv ���l��fӇ�a�
�T�s�5��\ip����p�^�®�O�@4^ZEjB�n됙�ʵ*�(�����Ǘ�:s�/�L�D��f�qK�3�Bu	�|�i/��ƴ�f	վ��B�t���|�]�S>����=�w�QCez�ԯ%>�̾&v1;�]�!����w���{�U�X��
0�7�X1�h��P��㺼�vB32�KWQ{��Q8$Fh�����1P�ӓ�#{"��V_!8� �w��<s�ևK���⮐��J0�ܓ~
���w�:`�_=�����O}<�j�x���-�{�u@��� >mH�e I�22�j>��⫥�3 g��	qc:I��Oʼ�z��Rovt�TT�@@FQ�\�1-��7gQ����2e���GDgld��7W� *+l��飰�JMN(��5��_'�Π�ә�:)L�c��@����B&�y����<�	PF49��/�x�|��0�+
b�=�*���\K��`7ڛ�.�xx�-:�s���1�7Zi�g�6��=���R��{ȸ�Q�ptoCP {«��i��A�^B���|R[u��%w]m�,�-ۍӋ�7}�_vy������Sxc���f�ܑ&���B
*{u@�ntˁB	Z+8�[�qy.j�?.� ��U[��f�.��*)9��oY��N�N��@:���Cq��qX�&�]����V]����p
'8Y�&2\����N
��2�sӝzȒ��.��	�kB���7�ݬ�v��s1Z�+�*�k�;6����W�Q�5�������dW�ن�/w}][o7�"�r]k�]��P����	�>z�[��ݸ:��Lu��/&TV�`��#1Q�L��s�Y�F��V�VRι����uYk�:��͓j�O�{���Iʗ#z�ٓKOq��{.�+EEb��T�4P�Ξ�JM�t:����y��h�^�.�w����-����v&*|cجn��o���e<ZܛbT�j��e/n�/�%�e�HT�;�yb�����r��ƫp_n�{�78��*�v��~
P���a)9�uA�]�D4����Yx6�"�A2���U���L��|R�Q3�o��<���-kG���[ĺ��WEp�ō�rYm�^v�yyD��.Q��zY��5e�u���n�Q�dºw- �Ijsl8��A�TjY��}.d9���&��U��6mk{"�d8��uˏhP�ջ����(6�|�]����c=��lN���]P�{���o����8�t�wv��zsUf��.23u�95�r�����w�v����}H=JW+���K�"�=�bYnL�W5.-D�/��?Z�C�$��mEe���X}�����a@�X��m�ߕ<t��M�Y\�lbܸ�����]u�´&iov�/4�5�f�v���f��p�H�bs�xL���YyRa74������@C�a�Q~�~ʩ�&�B�hE���y<���n��q%Ƃ�-ZaK[��Dž�9u��`�����+%��-��zM|��+Q��X�5Č�v�����ET������J�m�>��d�����	�B/m	���D�fN�vQ�ji*�
�/s2u�f��W;0�ّ��h P	8��*�٪ X:��k�^f
�tۥ.�=ޥ����J�Y�7:�Rh�(\��A*0'���ܰ���9h�zf%��l�ڸ��Zq.�t
&���`�G�І=H�l�&�偶����J��y�K��E�G�8aj�y������5��Jt&C�	��p��@�s�ǰ0�&��8^�z��äb��l�V7:�N�	}��.j[L�ks7_l���-`yZ�=T�ڕ,ם&XyJ�A����������u�DWv�r�)�����FХ;{��0#��f��ufR�V����ݐnV9ah$�C���WK�<H	ԩkF�yS�(�!eerf]闍j4��6�䗫p��N%��ؗJ&�&�U�.+�yap(�s��{�3��ֱM4}�B�eub�e��L���n�u_BMuod&�f�3m9�EI(ir�3p**�I6���!�ܼ�c/E@Gr:��/-H�r@���n��8Ys-L�L�`({
M� �D$�"��[=�r�c4�g2��RG�'^7���_-u+2�V;�۾����[3&����"�j\��;{��B%gV�<�\���S0�m��<w��l�Ѽ�!�XZ��mX2�v�!�ӂ���2�q��ڽ�B�*���Bja��k���1��j��@GcJ��in4M0n������0A��n<w9�D��7��q�B�=d�ݞ�&���i���H������!�̸��0-�}4D��#b]�Oʚ�\[~��"��ezBJ����HA�p���J����{Yfm����`�b��/m0�^�����M���t�S���Ơ�l���NIu�j}��m��-/�G���%G+C�
���\`5j=-�J%Q"π�Y1�d�}b����G�­��bb)Iq�l^{^c��/:�Z� ����5���=�|;��D	�?% ρZ;}s�����J޿�#��Y�S����(�{�u�g�Һ0�T�
�G\C~q�2��1������E�c���S��x��>�)�ܷ�z_�+��_QqZ8���5��:,:���b�_�<w�
~��;�;���K1�Lw?72�t�"�:X���P�Q$`�*����3A*j�Dt�uS\ElM]�p�{Yk��c{A�b7FT ���0��e�ʋ�Y���m@�m��s��ȱ7�Ŏ�}w��ɻ@��bJVd��)�a�7��-��Z�b�b�4Ȝ*���L+�,kة/Օ�O����9
�y^��������l���I+���6WN�N[9m�!0�y�W`e��FEa2P«S#%l���+N_�Lo�&$@J{�d�hl̡i�����+o��%��}	�B����+�ܱ��~�ѕ�	C��jz���y��0�#�I��N����2̜�f���a�Q۬�Dh���}G�wf�h�Ȱ��$�(�S���4}��A��XQʬ��4�ߔ����z�,Q�<���f��RuQ ��*�1DLU�)�f_B�h7�T��}>����t����D��1�w�Kgt���TcJ��0��}��f�Kxc^�y�K+��=m���i��:Q���A�D�|��;m(�)��"�� �/:�?ws��=L�r{�:��Z�{���i�acR:�}��;�S ��)����ܥ&9V>kDU�����O�G|$^w�2��Fɪ�W�5y�͵�c���G/qPH�Fb� ��z�]7�UyB4.�t����ܹ|�U=�@;�x�$�U)����˵k.���uP���j�bvr�����qjޭ<�eT�t(�V��OuS[]5�2�m�뼑���7nD=�觕���;33���'�%P^�(���y��_L�_|~1,I��,ZP�Υn�	�a�HJ6�pn����	E⫧[�66c��:���R�V7�ut�n�_
�ܡ�uhr�n�^��8gk����^:&r�[8v�[�����0�F`�����pwvR���A�h��*)�1Q;tn;M��
װ{��f`[^��UL\ƞ�Я}�~�y�<t�8\x?ay�$hB�PD�GD��=�coآ�oc3<��H���D�9&��G�TH��#1��3�TnҀ˃���1SX:�g�ȳ��S�^�
�x�pR�S���2/<Y�qkTtΪ��$]
����6X	�N2u��Jɑ����h��a��\�VZ��>��4/Χ�
����L�y�]w�K�V��s>Fػȡ�Q:M@i�<�y�ب�UJ7�9ޏB-���lH�K�|hY��y��#�e)aUɯ3�����3��t���ϙ�p&�C���Ѽ��;4=�N_n!ݨס��[
�#1�~y���V�M�(�U�x��Z�e�.�4��^پ�/ZbB�]Z������УXM]qxk�8q6oU�c��^W��g
*4���ؕ���9�Gi_��l�߂���"m�3��e��5MY�<��7��(ꌹG\M�2��`#���k'��NpCb�w��E����i�D&S+r'����ص�L�j��.s�tE	$D�f3:n��[��߲�HO��nBK�Uu���v��w�s[�b���D2�qi$�3FWKΠ@����`��<UB���f-w}�u>�4/NnyS��$�FM�W%9[3��	LZ�79��B���ptK3N����ҚWLCZ���m�J�j=�3w9ˬ���q��#C��|o�旤F��Y7eƊ��x�p�z1 �`,��"�_$9nT����x9�H��Oz��ҹ��=tD81c�w�}}E�{�8*���p#x���Q��7��#H��p��J���#bٚ��c��BqɞWz�J-{�0�o%�n-Gww�H�u���*�ĳ탿y���p�����H���e�'.���+#EE���%�tՆ-�\Ưy�޿�_��h�g��@��Ac�&��2 T����=`V�G�
�����C���vh�_>ы���_s���E��fh�;�����x�`���3��V0?7Tqq
<`��Or����Y�42g��"�U:6�Ç�~��sr��O��֗fαj\���O�<�eW;�ax��p��
[sمQ����Pf<�ؔ�����d�n�(�'�Rף �x*`�["uڳ�'��(�53HQL/p���#�f;����dw��fQ �^��VG�MV����"�)�xrf9E�>���k&ЯB��8'E}�bzu�	t]�"�)F����u�vB;G����P��T�'�sv��nNy�w%�͕!≓�՝�<�V�|=�'�������[(ň�ҍ7�5�o �>�$���?d%ի��d�ޔ�>�[3]Ǳ����{0V�H�����w0R�3j������Je���n$,�y�s���Z�5���u��N�l��\���OEeuM��egN���u#�,������$o��rj��v��z��=	�K��^~r(��&�y�S�T�����vr%��?��w�ߍ�Fb�g=fLt� }7�(L����E�%�s�������c�{Y��k��R��I�G��]�#�E?�nA.xu�<^�]2'��S7f�ۗ
����*7�b^�f����G��`���Q�N]P@�E^:c����GÎ>PO?tN���a��Q���S�(x<��Cz�:�h��|�&�6d/� °]����F���o1^��W7���L�oӮR�!������v*G��V��֮f�}P���j�`�)�6�0Tnϩ�^��w��Ւ����&t^:ߦ ��U+d��q ;�{��,������lI#�p��eQ���D d�k��������[1N��\Q�B��W��4��\(��yo�^+=�w�"w���Jr��L�?���Ou����M���d�Gg%���3nl�����ǿ0�0��3+ً�˽
�k��$~�`�ڽ��U�����6�j�G��/z�Nu|$�g8�Sp��85����{�Ͻ�ī��Z��l^�5��V7\�鷺J�2�G��+f��(���6��Zr�5��K�*�]�2js�#^f���=U�j�����1&�:R��K��7y���w$��/)tS��/�&��sX���w�L?�eKwF�	hR/u%5wt���GL�3�6�_�O��h�ޥ=~�s�/��Q����|�׋'��=�^�B�z�#yxG�-�0� o���n���=���dϥm���I��g��{�,=⒛����#9\�wz�6�y�9՘���Q��{��%��;bT3���
�)��s}0�rS�9�na����Z��e�ʤU+�z���a�07���Ub&�s�Y\�h/u}�Qu<K��7N�!���m�_�����J�^�����r�\��4v���RjY���c0�����ED�L]�����Ur�\QQ�pa�����̘�3cw:ߨ�g�$��^�������S��#E��3�s���T7`���'"��Vrk:��� }�i8����b�0zj8����
9É�[��P�R�������ekh���yVxWZ�*��W�6Ny�	���p&����#�M�Ih{������/˱㣦ϨPt��o�����,��x�F�9�����D�����".Ŀ'1�b8�cq��q�\�+w�	�|8`��#�eh�'�d���n���Љ��v����'�:Bs�q��pLr���A����́�wMc}�"Un�V!Xuȧ�w�SWY��:�c|;\�E�pk 2�{k�u��ϐ��	�� e%@C5��u0��e���<�i7c��{�ܢ�eb�}H���-�<2�Bi]��<���n�\%���S����L����t�P�w/���B�!��>�:b�۝ާ(@���fP,�<�Ie��Q��#�(�v�{v�Y�$b�<�qC'�O�g����KWz�(���O2�#��sj�ປ4�_�e����=������̪c�b٩�ʕ�5=�>܎*:~�!����:+�蘞[��!��1�HI�^�c��[�*n��2BC�5q��Ӝ��g����\v�ȬZ���g���'��q�GB���;w
��G]$��mօҜ9%��~�1\�'j�1��z�Y�=6Sٗ��pW=��e4��$G���N3��P�?T��y
B��\��+��^Nx>��M�S�������[��1+�*3m�.��[<�h�1��X�h暂Wl"5gIտ�c]p���ԩ�~�1h��	�]�����W�}\�5�Q�j3wq}����U̐��y�XMy�~��u�@�⽽��U��:� �������T�4�`>�ư�d��s�`&�14�T��\����������`��\���hC�Q���n�/E���z�,�)e�|�15'�3�3uk&�Eh������r�jR��~	B��#x�`�e�q\�����^�X:j_�jYY�.�;�Ĩ�,MwX]�F�Ԯ���t�����.�Eă��W]�*Z�D�U�	Ľ;��7Ҋ��+VS9+Rʛ�s���넶�p������!'V��n�,�Q������V�zΘ"p�	�A��32}{v�t^���&�+�|��P�k�~�T�3J�!g۔n�Ov���Y� ��uf�E
-����>����=᳦x����(G��~y�{��RR�T�-%����)����ᛌG������Bc��*��-�9fa�7�g7�_�S�ڇ�u·��}�DhY�K$����rd�ɉȞ�< ���5�)x�p&��ؐ�z2q�qO0l��qS���/x�Wa���qp�� En�4#� v�ܸ�m���\�mLަ��"�x�W@V�����'�[����U$�ތ\�z.�̒�eYs0F$�Wu:��ʵ�y�(���r�ۉd��dݨ�U��l�00t�ytM+W��D��q�\��*��s�rF�<�$[ ��߻����9E""<=[�n�=��`|��U����t���>���<��(�뫹q<l�;B�-�G�<SYR���h�h�^WNf"b��;���ϓ�خ1�0hq��o�;�����2ǯz<hd ��ħ]W��I��e����SN��Ӡ�˙v���n�xʌ�+k��/7u�����	w�o�q�Xْg��h��C�6iqS=q��6�ђ��i���¯�·�Z��6A�77Wx�4��ק��O���jh��En�e.���׷���S�´]�ӳ�t/C�j<�z�6��C	� �U.���ȽQ�uN�];�L�'k��Afj!"w4�t]e!.���r٠-lY��A4�1V���sf��pս��0��Ǽ��ͻ�"�B�{�6`�E$Dk���9��V�����n�8�LO�h'[�^�� Ix���ޥ�`�˽�j?�\��#��w�W�}�fd�V�~����g��wrL�9Q�%z2����U)�Ͼ���GGf�Ĳ�L�3Ү����@�nϦ9����{~ü�LeP�4]��j>� tHׯg2��"Gh*uK�F�ț�ɹr]}1ϯ�7ok�s��otД1G�9#ڗ��[�t�e��m��,�$��~[y�׫���7t���觘v�\N�r���L{�_�F�(h��M������[�	��q��uW��#�2����:�z�;�f�sC�-~*g1l�B��≊�v:�]gUܮ�RT�*J�s`{��R0��|��q �L>�����ge�L�� 򍏩K�zCZ7��e�Od���%�"������z�R�(ݐpd��I�T�>Wj�n�3KG5�^cx�Y6s%D�ڰ"FZVe�;z���0�k�Y]qәp��3��gY���}Q1������ͥT9O� Č���ͮ�}���S0�8��v���;X6�s$�]f���v
�6��߷�8��"�h�S�:tԭu�$��c%�����m��n��7g�c-L4Ӛ�����(HP��Ǳ��u����S���ı�V��}p��1�d��z�T��{�^Np�A�o�]5�-��(�`�˖��\�I�V�Ra�(vb�����J0t��<������K�CV���B����l�T�(�ps�u�텱�X#L�ĸvL�u웯�w.ѿ�߮��|��P�w�2�7���P�d�,�N2���u�� �WLt����=Y{� j��vj�4
������7�c#X]P^���C<@͐�����foƹ����1��}\�����Q��Z%6����*���렊�?&<�b�Q(�<�3'���^u�����X3=���{�ꃙ7G ���;�yX����2aڥ�c�ЏTN��2���<�f�0����<F��K�Q�l�/�IB�t��Sh��Z�w�B�T{ݢ&x�����O�=fi�v����)��,��E��Op��Y�&�W�l׳:��+*�ױ�_Kk�L�-�e�S5{�SSغt���rN���'�]h.�����糳 ��"3r�^E��Z:��ۙ�`�B�hf�OWmI֌tݜ�xպ
2�q��3:���"��N�S p��J&=���y�R�-x^O���E[S6<U��</pbHw�hs{ej��ll�N�T�5�$ ���70�v�3�{�j��ն��*�z�%,Q��^뻔�y�6Liw5�J��ξ^;v
�xU����(R�y��i���Dո�MJ5
r�N�5i�rH�1��lLE��ef�sr�]���0��/��5�<<�ֳ|��w�D�.}ꖦPA��S- ��'en�ٛ!���RQ��0��IB��ͬ���K��+=�D$���;�u�՛�$�a[S�p�F�ۗ���7�o/O[&�y���+Y�6��[V.���׫��C�������G�(��׾��I-��I����t6�mݕ'<�PK��Ѝ�n5nZz�w��߸�����kb�$\B�H^n��Fh�Y҇3��*�VҞj,���%��5w�4�%���	x��Q�����F�2��=�!uod�`�D�2�t��/�,N�l�Ҿu��+%�+u�3Y�4͟u̡2��4�i�ݔ$�l����Z�k�����t�_��~�X�[����|f�`��Bw�k���$�8K��733[x^����)Aewu6���3gz���KhS����uuI\��޻Ýuw�
T�<�4u��I ,��OV�����.�v�(��I��8���[��3{�{�!C"	j.CT�֞�E�7D���Hn:k.��	lbU�V�c�ԌklW o��Nٹ�:7�o;��S/��u����׹�t�V���a�agm����iX�6Q-�)٘���֘���	F�9�u<Ʃ_EQ���o,LS2+�P�=)+؞�K�58��7�~^��N �*t��c�U�8cǹ�X����iY*�����O����@����g��u�L�4Y;*G�+����K-��e�4�i��{�OvW���DG]M	%�w���ꋦFO����&,�/qO���q�q`YE��Z�����u�\#ff��|�Vx&����ʝ�p.���u�c�,�iǇO<��&Ydu8x��H%���wl�Ɉ�]sR�m�u���;G6��N��cŜ�d,8=w#59)�u+l��&�]&��qRАn�P��C�*��,]ܖ�Kd�Su�Q�ɚ�.���F�#v��mAx�(��u�%���S��
�՜d��YR4r`���e=c ���N�.+�h�Ѧ��t��X����ڌvq_���'�ݠ�gJM]Y6p�+P`z?q�\���ڍ�so�Mo���;��H��XUk4P{V���p[��=�x�@i�澯��-n`�K<�n��׹إ�gBq�l�/=��]�S�W{;ڐ�}2V�FP�;	w�5����d�7���0���rnȆ1,\���7t���Sr�]w$�����w���ΩJ�0����h�/$ϼdD�˵�۵Y0Zy�Ve]���η`Z�C��jEeE]aK6Y˼�5��oe��"����7�R�wM���v�en7���ީ`u���{0��x�7�3$��4��;W��fʃ�c��w�iڕv�ֹ�L;J�fd���,�:��cU�l�S6�Y�s������sv�-YvcdRX����q\����L(. ���(����&�RR���[[c�}�\�Y��P+�����J����ݹf�K�`�#-������:�Y�[-Dˡ5�&�@R�T	Ӊ���VӲ�v�HV��;^�w���PޜNo9�cTN��}ܞl���lP�HǪ�彇%&�xI�m�Hp���G�}�w2�L�ͅ��� �~�,}����e�	b��W9]fkv�u��]#sy�N�a �9�S5�1��z�eɀ���p�V�t<�gi�ª�ʵU7KMz�~os�_~8�I���Hc3g�m�z��;2���Y�����fY�����R0#����^��{�(lg?Bo�V����s�k�|�a��T;�qU9��� qS����6wJ�"v�ɦ����Ψ����6͞K*�g�j�k�R�HAG��Ϫ����4��^���Zʊ��/i��Ӿ�Qû�B��	��}y�	t�R��-�tb�b�{k�Ԡ��x���X磏��(&�{�f�WH�QP�k=}u����K�6���B�-�Z©u�{��ރ������\s�F���팔"�F��Y�5�\�QU�}x��zr�*��p��B��I�!���Z=�����^����6q��m��>���B\\Pp���F��h>Tp�b���?vde�L�3�|�o��b��������ͫ`߱����©OϦ���9�\�8D��}�"����,��w��mo�*XݘT��'!�<ۙC�حc�~���@#���{\�l�4��3�
���N5�U��s�n<q[�}^��S�B�4�Z�Ō�Vy_>�b�N_s�9����!S�L[;M�����o�ohHԫ�ap��\�r�u����M9���ɘCT��5}9���[��R�r���+�*�wV���On46[�d��q�u.�t�C�[�E�r���Wt�z��j����}	� ��z��g�m]zb�gӃYW���p}��WM�3�,>E���w����Օ�қ�Z3w�����ҥ���f��D��;x�{��Q���gh��~�Gt;�oe�L�o�{���B�EY^|��K���pp��r��Ks�6(Ͷ<k�6���*����J���r��з[�]������2�>1����d��ش�;�����ER��$�r�E��>�n�7	�pK�H�3~��� Շԣ�x �x ��\߮V�ߠ���� ���Xyv���'c�4�
��]�u�X��23~�����n��R���6�܁,��@C�I����1m�����0�ݕ��ZQ��y��Z�:e�>t����n��v�M�v���Fb�6�F�B���0���[�9�`����:@Շ36u�U�����(`Lb���y���~����ϡ9�=w&�r}Ս&�Pލ���K¶�g*i��:�����T��_=��Ѭw����y~Ϲ]�����(q��޿���z�L�W�}y�D�g\�w��n�p��8���;�/GU�G]�˦h���թ��}�I��%�c�"�`�@����.~����L<aM�o��&p��wDz�jfiU��k;k��烳he���c䝲:���}�+4��F���Mu��y4:�l�V�Y����OkY+�n�x(٘ӻ賠����N,��VB��}�z
 ���Ʒ�{�a�o�B�1<� }�ۀc/��f����7�J�뚙9@��y�=�~팻ɲ߸�I�,^W�J�k�e�3�fA�A1�q����Z��T��֢�u�o�<'p_K�S��FǈmM
^^�P�����8�����2���:>1נw{��y�//H���;�x��6(([�LI�b��G��s^����M&�����1+��y���Y2󔭞ޅL��B޿U�2�*�̾�W�|�׵�>��}>��fm��#=��+�׮��R�[�u�1�x_N�y��.���7Pc��A���=�������<Ž���m�'�	׸��{����7ư[�m�N��������ڹ�K�������qmM�+T#�v������v��{;!G��ڜn^�λ��Q�4��./�yN��_Mq�řq2̊�[�c�|&.��X����[���i.F�)�T<��}e��'5�R`��Ž����.S�^��E1�w��-pm;~T��M�Nr�8�mg��Q9Gv�Tg�f��`�=�n'��V�^���
*�I����7y�k2�,[��ʕ�N�Y��sk[�kʐj]P�U��@��ېX3�-�f�-��ε\G0A�=3ogv�ީcz�1a�vk��'[�6�l9�c�&����񡤘����Ə/��&/O):ɕw#1���9
�N�7;��(Ɏ�����z/�C���Tw%��NB�F|2PobZ@�L'����뇠��k5���[|��bt�*�}9.�yi��Pugwl��R�j6=�<�j>�}䷇�A��J�d{1��nb�҄+2��8��z93{Gר��O�;�/}o�>� �r���'F��Фk�&zW��h��n��Rq�3��u��)oӪ\��^��o���Et�D��ԭ�0Y@�����S�&�Op��}u���\���3�܀��ösJM`}0��e�_�,�
����󲺮=�ˡX���m�\��c�\.'�
����

���XD�����a\.(�>�b��J���2��G�:.X�0ݮ�����?eTY���eiۄ���I���d��B���|��D��ܨ(a
K7�f�R����d�R��R٩��/�rk-'���8=oƴ��Up5Л��Fp;������v0.�:.�aL`J|mG�P��7<��\�nH�҂G�K���=�-��n{���v�mޝC��TqT�8��ȍ�G}�S6E�hi����+���O2����rڕ��B��f�$�ܲ�n�eV0Z��RM�F��Mm����k^'Y�]�H\qJ�K5�W��N~�BT��Bm,��e�N��zN;��y^"�i��� Y�o'@c!����5����Z"�[^a�����������̮t�$ͩ�@g|$�<p��ۦBc�7G����W�� ��hЋ�-S���Bo⧇�|4[���̙�˨���`#�m{^��o(��k�댟�~k��&�e�;�`��~0LTH0���0��4�[��g�㼟t�S���K8��_f�ވ�=�0,��+ɉ#Tê*��J�d*�5��Go1��J�S�S��ohZ2\�^@q�X#}JF����x���Y.�'*3�(�✍�Cբ��36Ѥc�P�\������$��n��9�<˶�csQ}7cB[Q/b���Ow�{���K/�7%VB	f�Q5�,�E[p	,�;�r�Z��	��^1�]9�Q�kg挃9Z���ץ�� �*�=�pd�Q2�)����[& ��+5�d(���{+#3��`c��47V��&

���^��pH>�׳��6c�D�<=z�ba`Wq�`�V�k�i�ģ�FX��p�L�ܹ��xƭ�4_t���p;1M��\vú�є���:�[�?Gr�]~�59R-��kC{�{�z���.]�$k5�����$��s�W���Y�8Aԩ c��t�IY����V�U2�7;4�q �̵����>�'�}x8�����Dk�W-�M:���B��ӮG��v��R�Ō�4f�\[��A��͂_�6���Į�j �~fI���U������Ȕ`�R3;,�(R�Q��1���3�&<�vP>{�)�/JT�L��b؟���ܘ�ų�Pw��=�^H�e5`?�v����r�!Wp��$���Q����>��G�t���@����Y�.��$�%�!;'�S�����zJ���c���(�׽m\α�-{�ג����;��4��#��1���(ۺ��όGtm�<m���&k�Ӂ�K��Z�\q�*���ȩ�3�������r:}��t@��ϣ���'s�?4�F�(Iȳ�n-z	��_^�v{�T>�v�i2-`��)@�=S,UI�Em�1��듍!�dL`�I�������{�t�3��i�+�㮙ɯ%_��s�_��=ŋ36bL�2�1}Q��9�p#}G���C�0U�k`��.�� ��.�֏�lr���l�Ωm�E很�BU��*sx�t\�<�7����Ks΢�Ռ�iK|��f��mK0�@���F���׺��t⌽UF
�m¡�D�wTt��)x�P�i7��U5y�F�iG����tN��
�%](���S[Ai���	2�g^�������|��zz^� ��R�XηNm��j�Y�����䅇��4��N�Ù��H8qX(����,�+�ò���1�u���>`S�vAW}8V%e,�*�|������s��G�# �~SVp-��1���y��{0b�Ϥ���{�w�T[���յ�2��wJ������c^[�^=>��Đ���\!�xHeL�Ǫ=决��t�z�N�C�t���/�*�F0��<"�}�*�=��r���j.j=�������׼ O��~. ��ݖ}���z�g�oT�ȳV�>�b+�E��U�nS��u�dt�K�V�A0y�Tj�E�6s�7���S�)}�$�D4$��P�(����Nc"|��D�ƫT�1�x0���#MP��M��:� �퉨�ڰ��(�4�:�����Q��S�;,{�<n;��y��J<-Y����I���G��9j�YXe=�qC�u�{,<ut��Wf���11��OBn8v9��ͯ@�C`��Z�8��/w��bK�E����˫N����S�\z�������+�U훑�«�n��*�&�C�Uvw{Qh�7��n�!d�P��)'���Zl�h����vs\�#aρ�����:79r7E�W�^����uv1sNH�0Hn��0���9��qqRo�,'��]l���v��D�:�]�<���ZeاhD��*�)��nT�8A�����6����F�%���j�XҢɶ���}34�Y�AE�)h���#b�^����IMP[�#�+u?ױ��6F�}�K6P��/7J���h��p���:�Er�B���pؽ��v���P�|�+[�����]/|MsW.�����U�C���93B���<[��g�[�v|�c���znl+�ads+:�gxe󵞫����E��;��x�e��a�"^L9Z�	���{��qÔ/���ӳ�����,לo�ԟ��<�+��׌}�'�DT�9��_��t���G=<��c�U�+�C�/;��9��x+G3��߼��zP<���wK�3^E�[���NBr谄;诚��x����B�r�u�t�55O��J�`܌N<���.�Z��¾'�4�jH��j�	�޳u��U�0����ā{ �^ڬco74p���$5>-˦	�q3�(H��L�O�����%v�M�/`I�pBZm���}�����Tf��Z�(Eh�7�~.����;��˜7�����sa�#�ks2u��3R�m�Ӵ>x=��BݣдyGm߫�w������E]f^�,G�$=S�[�)�]�M�Bl��v�Ai�(>�����[V����Ы�T������r�O�=4ߡK�Y*����@�E���׫om�+�`��*��s��s.гE�ڲr��u��p�-,�D[�.&]��ѭ�Tĩ��!�Z�E��bgaǝ�ԛC�w;�l�%+|�M��v�[��%�(\9}���g��vr���ʗ_r�*^s�t�ծ{#p�a\�չ���$x���NE�ԈAAȝ�B���޽��۽�^~��p*0��o�v�`��.�X�EV�g�w	r�s$��C���Zv��	R'B�7�@F8�{�ѝ�闄H�=M���W�<ԇݦ�_�%�϶
��Q�J��C�a�qV�#K�S8���`u����x��;ɸ�1��1�ԪE��ɾ�h��d���@���#M	�8xCڝ.~��BӵuDiʵ�j����0�f<!]C�և7�����(b�����q�mI�6qf�z�'˞FyV�#���Ω��J�'�#i����--[�>�%�O�(��]S=q㽞7b�Y�[�Z,�%C�QC�*�d�)�����ίO<�{C�_K��c*�˯M�"P©���a��yVH�>���U�7>����Ŧ/P�1���S�0L�y�7��f�W������<�[kT2x'_]�+b��ζ��|+F֏RWQi�t'I�kG�k%E��{�c��͋����}�p��u�6���J՘!J�>��Vp��:ۙ9��۪�wec��_��/!�^ �(����&��V�b䀷MT`����Rv���Ղ�������SG��%S�G�!h�����d���j_!�O���V���J�J�,:�Z���g
̆Ρ�D,7��nq��ŝ�/�wp콝��C�ni]J+��x_d7��]�((�����s�������?Q�tT�bڽ������-kߩ����^gh��-��{2q�{ �>=o�``���4/�C��Z�h 3+bV�;��w�A����.kâe�G�!5"u��HO�W��O��tj�-�Uv�u��"h�s+7�1�U� C0n:����)@�D{١B˘=s��;}�%6�WW`X���(MnΏWW=7�1�|'�E�#�){������L�B��VVͬ�	��HO/��?<]	���8��Dۃ��']%��* �+�ȶ���(�b�Ț�n��A���{:�;ްg�w����"Ƹ������:/,���H�����P�_"6ڪ��*���:��r�W�j]�����-DÂS9�����R�Ɵ�9���߆�wH�\����Nr��O��+�6�ӉK��Pg-I���ݧD�ZaYH\j�!1���{����ƞ��� �{͸��q��ω���X�y�(��S�p�3J����O}��B��}���v�xL�Ƣ{ ��Au��>���<���2\V�����M��k���^�:�1�����'�J��:�Y|@Zl��[!!-�ͅD�+�f͠�j[�M	��l��Nѹ�
&�5E���LJ��Ѱ�!v
'gj���ep�ilg@E���/T��~l�`7�Nq2^����-�����^rv�Y��*�nr�СBZel��BI3N���gfV\�O�b�8�3��b��h��;=�.�~�}4"""/{��U�~�ً��w���iw5�rW��UQ	E��H��d��/e�Nm�*ïo/�)�T"����`u�j�:��	ǲڂ�V'n���N��"�_�{�uNM���J�B�"NV^���9�|�k��*�'^`�&�N�h���k�I�W֮ r>��ܓM�����ό��ڧ&�zUJ=Y���諒 �nw~zj5$�oo5rB��Mճ�Y��jP(���T���q�ǭ��L/�!hyמ�h�oo>�Lê:�JY�Y(�}G^��[}��a*�����V:�0^��-�.�5v�����8q-V�S���S�M���l%Q']�����UG��+����R�aP�L�C��
8�I-)��n]]z}���'_߮�:��-���IsW�Q�����Go/����Q�뾛Gy-��f=V�>�V�W�)�7�g/�ᗘ�$���D���Y�u���ާ5�O�B����#Ǽ�������,YMp��2I	�L�,�h@B��ߖ��b�Sp�f$TB9���_��c\r�{2������
���CNsތT*��'b�h����eЫ/r�+3�H�7�V�w`[��}r}u+��K��j�g�;$�_����4J�ϩ��ޜ���z�o�t��u�X�w"�t}XzJ�j�qޛb^�Q�F�	rĹ�)�I9_�5[������޾�a(ȦD�<�VRO��#M\#O����yۚ�%�����W�b/��E��ĮfHn�#�)�� �*�\�yT��lM��D�[���IOw	,�r ��9�NՅGe��q�rL�yZk�����5�Л���	���N�����X�q������v�^JlA3��w����|н#kH�Y){�d�œ�s���f��ff����W��Y��1km�껎U�wW���G�G]�n�-<�Ưy�E�iSy��s�0s��s��℘mZ!�ѳQ���*V�Y�,!�3.�ЇxR�e���T�y"0�����`��v�j���������Dw��e�uØ8����ko������!!=A��`T9�݌$��M晚�;���0fJ�1'l�Ki-i�����;;%���W&�\N$�K+��Ff�D3;�f��%��g�#�R�ZZVU�Z��Y����w��,����]�շe�7Ý;䘎�󣝼�k����n�J��#��a3ʎ��o��U�l��� �ige�(�5i���aI�t��.���.�K�id��-]?^�Ɍ�ܸh���i�go�.���]8JV�#�,�<w!�hvL�d�6�
�ؼ՝���TY�w%�<��Vy蛋��N���<wk9�w�T�G]���2�j�Ks94�+
J��Y�%ݝ,���/{��ޭ���W�]J�I�i��̺�(���eU�Ԭ+��8�����i�bc9���8r��`�����K8� w�����V���,�2�ޫ�\��g�R���V\�ݢU�|�4I�r3�m���z���B z��)
0iVp��쥓��P��u��V�L�e�ĉ�':dʗ(��a��,���O��1gH��پP%���T-߅ ���Խ�N��?(�����V 9��i)��l[z�uT*���#2z��&�o]���GX�Q;cT�O{ȶ��ӆ���� �Wψ�7�Q��g��Lu�
�l�mV�$�C�����w���B'>�Pc��ъ+G݆�知�w�b���]R�Q�Gb�i3�^��@��j��Xū� ��5j�����l� �fٛ��7l�`���}�xk���A�E�ϳ���^E;T���3�1�a��^��B�K���l��X 3�c܌����#�ӱP����s�0{g���\�UIi /�tt���׻W�ǭw���@���iķ�p�ۚ#����
r� ��n*)
;1ޢ�˖/S�G*�|y��v�c*�gT"�A���o�c�Y�*y%�0��z��g+e���Oq�}�w.2�x�˃����{�t���xr�o�G*�������|�>Z��6��s\,vΊ�u]�:������5�4�{��t|���\����r�_��si�U�T�˿:�<a3���и7�oP��^޺6UY*'/gp�&m����]�ZEq�b�W^��r��-���X�[��bz^��&S��9�Y��J���z���3Y��#� �zR�_��g�eCÎ���0zt�P�
�+��	ɍJU�]
ߨ�z'��Ӳ��9�����~ꚶSQ��N���Ɂ\vf�M�ͮ�wt��6�o���g��WsU+�>2C
k��ò�Tk?[�;9�X�%2���ю�Fb�������}��!����g�bt/C��uZ��9��FO�ĉj���h����A��kË��u��h_L}���[r�]
�S���c�[��y�2��o>��R��w��v��aW-΁`Nu:�g�'��ub��G�!��^o����3`}j������+OZ�v4�vf&��^�Y��ғVt�{9��C�l}��$ٰ�E~o���ԗ�o��=�����^C;���E��
'�/z��g͞�a_| 1|���n�j3By[�j���E�N���3�'�N-���+&��'�f^�`K����	�_�E9cÈ�(`�2T�N�mk�� �aF?�s�>����AQ�i����3�E�Ga���yKu�#yвOir���}�zʙ�7Q8]�sI��l��|�,R3Jh<�,ա-��z{sCj�lp֛�y��qm����6]D1-�4ɀp����M�q�9�
�1K�ݲ�]������xA�]��q��7����O�nV~+ZaWٗ��n���}/�({�Q�g��'o2���*�L�^��h��g��9��������-(�sOndt���O���]��b��s
C�ۊ�������iy۾�����ΌR�rz|+�OXoA�C��y+0���p���Bzdm��@��F��&%���UġÀqF)��������(A^ݬ69Y�} �l�T�%x�Q�|���MG�6�p�x�;#q]+.y^���(p�2���Y;0lj�_1йWD�Ӥ�r4 ��8D���4pW��~C/�՞��dn�&�G=���ȵ���ԩ�ZOo��.1��r.*�U�Q�SJ-j���!�ne����;�GE��.;����P@�r\�s|�� ����LLj[���'7�>'{k�ȣZ�z3R�G�g��Dz)�Bh^���U�y�8qj�����=��9��S�#���~�v����
�jv������z(ݸ��M>�3G�~�Z�Et$�9�34�ZR�܋��6�;\HYQr�]�[��P�y�����nvFu# � o�23. ˘n�}
�5.:�v��6��K����y�.�}j�\ͅ1K���)K�9S't�FvZqr�N�'�1ی����P�ͩvRk���@���s�ͺ��/����b��=���1S��Ţ�j�u����!��q���V��`��ؔj��1ݽ���W��S�QD�:�����R��'�f�kbc��^�~%t��4��jp�v�a:�Kָ��X�V�/x�R�R��>�s1Y:m�b��67h�� ��A�Yn�o��	'	�e7�&����-h�/.F����F�ӂ��y�mH��_k���l�F�U�Z�/<��QC��J�7�-�93�
jQ���FF1��sݗ
oJ�ʒ�zWHO@�ΧJ˿E~���V,��ć�l����7'u�Ի��i�/X|w��m����&�כ�/5���V˭��r�����6s�w3lw(ֳ�&���C!Pwn��F���컜*]�!�74T�7�h��Λ)�=����u����>�ng�t3%ҭ��*}�"cٚY=E[��������O�t]]tC�W�$BZ�I;_:).��p���Y��L�Y:���q*����?]Ei7p}��������;;c)a���)�,��b�J,`�K9��`E҅��Tyws��*v�DXp.F�a�2@:��$�v;}�pǱӌ
����_X��q��2f���\�L�kc8ƯL�kؽ���}d}Q���9�:9��v��UI��uT������+���ⱺ[I��N3Eh
~�� �tb�Ò��;�5�7�Ooe��҆�+�']�+xS/"�S0tY�Y�{���_��t�6��2��R�Ɋ���3啥1\jM��`e2ܴk�n'BTC��<T#��!��@�.N�If	s}��#�f:_w�:W}�,���^����6���hk{�R���;(�q��L�/8߇u�Rs���k�B�G����thu\� +H�ݗ��Ŝ/m����;�}\�8ol[ʝ}��ϖ�!O�Qos6�kxS��2�9Uu�;:}�a$�������]Kr���W>�Q�� ���8&��Wq��L��=aJ�Sl�|�S]`�׶k���w(q�.q��ѽ�öey)��##� �ƻ�Ց^�f�2�{�6<�Z�x}���軘v������a��Ϥ�b:�[Qr�'���`�י�>� ���t�� 9���T��3x��1G�c|�fW�0�o�=Q�yQ��(�ú�&��	�L��1�����ǆ@�[�nI�p6��3��
��Lʚ㽓�b��]�ԴD��;�?ln�d�H㋯m��d��ʝxl�y>��÷B&c���6}B�:��[���� s�9�13��V������0�V��%T��MBؼc��֥l8�iפ\�D!�I�kr�|�=M�:��P&(^4��N�F����>�	�y\%��k9U��c���f�&m��a��/qt��K�ߝ�C��EC�A�ז!|��㱜�T< �����{�c)uĴ̢�n��'�o�w"�;c^j}o�M��I%�k^�V\U �n�E���I'��s�=⾿,���7�oƨ�v���ܵI�gٰ��Ry���|�SN��n䉅�J㢏C��ԣд{�Ѻ�[%��H�?U�]�s5�;��g
��*B�"����V z�_@Ǌ��ԅ]dҍ��q#`���W��G�b����?{��3�Ztgѭ�y/�7
wu���gv�����n�r���w�ʄ��ژ�{^�ϑ���k.�d�k+���gù�oB��^�ۇt?X*<2�y�i��^�r`$C�Q���=^�ȤǯP��_��ٞ�+M��'�#�=�g~Q��1�#��$�
�:@���pt�.�A��3(�dw�m�l�S_�K�I	�d�];��_��ȏh�"���2�d�4Nv��͗�Zn��7�Jo��]��3�QV~���3B+��sb�Dǂ�#I��/�=0"c�M�A��ӹ��^	�=̽��j���4�L�T;g��/����9�}k��wOŸ���r��l��W[����ϥf�q��Oލ�w�nH�b�x�)����z�2=��>9���W}ܯ�-���LNJ�x8ymo��$%~�=�X�4�s%��	�[E�̭�X�:dh�9i'�j�o6�m��!��
�iy[��+�5oa궲�W-�A���_�ʼ\/�ԑ�Es��N!�j̣2��7 �YM�R�-���̼i�:%�p؎6��"�e��7/u/�����x���w���{��1�w����}�hdvB&W�'4����P5#���y�OL!� b8�"7j��8ߝ�k��~ZPC�Dй�«oT�{�2W����G��������c������_'��w���.���}:� ը�P��Zy��t֍�0��%YgqyP���*��c�8����|Lׯ�bF���U�L�"U-���Ɍ���R�蚀��Ƙ�|�C��a�E�\�����=w���q�~���y�"�#L<�r�(��\O;��N���Q�v<�yH ��p�#&�<����3:J�2�8c�)�v2��Q�Y(�0�V�vܬ|E��6"���� 4���VW_���5N[������阺��Κ���uh���R����-�l
�97uʯ�%����Q��c�j����7�G���ɉO!���gl�`�+v���rP�'J֭}�qn�8��a��oI��qdf;2~��:�A�VfDok���G����ƫ8�bB���=<F��`U����;Ѩ+^�x:�a䑄`VE��T��R��"�~ޭN�(�o��@Ϋ���+�T|��t^�`�����D�}]A
8�-tG���"�1OWMw����xO���9(��W��ro7/;�qx6��m�46�d�]+8�NW�]�����5�;ʒ�U,�h�n���sBw)�i��xe�vb�&$��jh{
s�A�!-�OP��������+�dr��1�y�7��n�'J�[����}��V�� �����z�Tx�U��vf���D�I�˚���A?�b~"�;��**;Փl[Ⱦ1��I���=3�xxa���_�Ce�9����6�m�g}4}.z�/T���7ܕ��e����XA��Y��L^>����P��(*���$%��뜚�y��B��g��k�Z/�l��TNv���ʄ����VFEQ���]�2�l�^���ZOZ;p >x�H�ͻ��e	-��8�����!k ?J�"�5���z�V���=ciԫ�ͻK��s�D�d���<��	�m������˱�L��檕�������B�W�@���
uB�etM�1J��ِ���4�_��M�9#�C8�n:rs��ќq���x�U7�tl�Kٴm��s�P'g�Ǡ\��	x@V����fTvr�����Sfժ~������Be��B��F,>��?P�z^)��Ly0ӑV��5��:�T��U�4:�`���U,�\te�Bbx9|�]��������]�:�YO��H�J�c��HER��$U�m��1�ve�)X�\}*؀enuk��蔯�g4�9ٖ��*m��խ�gW_u��{u��Ĳn���t¸k���<�Eluڬ�9H%��f ��^ũ*v�=�"��B=o*:{��E�y��W`��E�X~!�-�2�C�Hy�c䳦��i�9u���Q��!�b�v�g����JP��͑G���_����@��a\>�p��TFk�13ѵ9<WD�˸����Y�|�5�����X�*��Θ��nB1��<fNa)hou'e�!�y��z�^n���M��WK�ڵ��<�k$f�~��`ϲE=�s��޿���9�*�!Y���Nk��>xU"���HY=���' �FD.��~��j�d��M��C����pX ���VWG,�4rֱs�9�yn�c/��E�< a3פB�]!��:~ފ���mw�.�Ѿ; ,$�3#�AF6k��S>�<Xvf=��P�M�e�X{�lM��Qn���p{$.
N�;F:�����A(��}Gr�D��Q��L�͖�"�Q�uƢZ��mN�^�����a�҆wo�������c�*4-�u��8�ˣW�Kc�|>�kl��s�RS73��&�A�FL�aqZq��5����Mh��o+2ue�z1�rv��εBoaٽ��y8Q�b@�+ں��V�:\yW�����l'�Xb'rs7V��p��&��j'��X9�hA��jФ:tt�\j����]q�����I�F���,;���u�n������Ɖv 0�w�����9�J~����|�O�m��8�����E���q~���Bc����!ᘮ�q̏�4ñ���˥��J�nT�z"�!R��]}t��3[=�@�xjK��Bk7�,ݶ�SB���/qW�$n��Ͻ|�ڼlbtl�$���o1v�D��dj�ϯi�Ԏ�'�,�%��ߌ*��s�ص�
 )�s�i��Js��U�1b��@���i�lz���~��d����%�1��y���0���gS��V��T��Uu9��9���G��F�F���ȹP22��@L������w��v~�������xO��S��Ĺ\��7�����]o��!_<�VG}�/gvFř�~^�^�v=lu�i����%��7�^EV���^yh����FO�4�/�ػ��l��6��60bR�X�@�O��3�<\�q��(��g�#�Fc��F(�>�?\P�T�P>�����'r5c���+if w�p���ŧ%P�9Sf6�D�N��AvcT5�9cȞO)��������|�IC��կV���5���:�gU^WeK�ʡ��7��۶æ��yπ]9[���T����]<�]�"�0�ZgIN���LtVoxu�깺zF-ތ��d儦�(��S׮�V�>Y���%�����.0�Ӻ���E�)��C���H�8�g�.�k��镼�^�����<D��#^-,&��:�c�N:S�vE�e%��܉Nܤ�D0U�|g1�m���. T/���1����o���0�V;��̊�r�����h�%j�W.��}���.h�<�]X�������f�l7�bôX6����F~U.c��sqK\��:�� �S�0"|���S����oT]Q��N��Vd�+a�AӼ�
����!��]�X�;ww��{U��H��vU~��6�/A�l���]�)�Y6�T>����%�⡊�*�6�%WOo4�:��LK#Q�Qj`�t�5=�2E�$�aRL����{:�1b]����~`��H�j�7M+�z�#��-�����o�o�4�N�J��
�y�(DU����Ҷ��$� �� ��� Y��NS��+M#Q3H)E�OP��[O��Z��Fv���̇	�+��iwp��Vk�V��JX��An���������f��]�W�>�.���_}�a ,e�b�;"q����E��éK��m�E����3<���j��I�sQ�������A�䯎.�n���u)&v�U���Wj�3�s.����v����-��^��*��N�z�:�_*�3��É���"���/b�^�(X�����D\�VU&�NV�AL�p�"*��̝յ����c������b����*�E��l��I�y̝*����S�2q�$�y�왲`�ܫ�j���\"���]*��A-n�����]�Y�e�+%gq��&Lc�e�wt��q�݁��ɘ�.�P�ȨK�sw��Ġ"3��L.R�ƍ�`���Uu�D{����u����������w�����j�il���M�V�Ƌɒ�)C�Xcd�t�&�Q�G	*��C5�2����[n����Jcm���:I�v�@DR�X�֯xS.$F�ƮMP4 �Ȱ���WԢy�O0��W���F�k���jn�M"EC�,^%g�˳
~�'�`_��V���G��| ��s��������'n�ע_RN��M���b����4V��1��Vc��;Yww|��X�R��mޙ��=;F��������V����ՏNu.y�z��Cl�]mE�v��v3O�b����7� ���Z�t"jU[+w)Bİ7FJ�`�&:�ƍ��r+�xQ���j��j.�lq�O�4b0̰�_^\O��nV��)bf��ۅ-p�pƄj�f⮃2�kCe<uA�Jy �YsŀAwQ�1j��[���՚+bp�Ke��5f��!o�h�ێ��V%����9�mp�l��������N$d�2#���Ywj���UwN���[�!�'N�T#��s�t[k$ג�J|p<��0ò�X���9�^���t=֬���N�O�ו&�C��)_(��B�V�D��LMg�菣�'د۞��q����8�[<��wC�2��`�=9�(ns��G<Q�u�vk/Q����CN*���ۇC��9�#����5av��(~y-�������W�ya{��Q�;�f�+�-{	���]F+�N ���eҳe�7���Hh��,��ꨔ	X��Lzw�`������=3
��BB�q��黍�9CY�+��fd��k|+���|=�~�̒wD�:�6�ڕB���5�-�G�k���(Q�ھO�QN��;�x��w�/{(Q�i�?�
(<�4l��~�p=F��K40� ޤ���� :np8�.�h+nV��Q�a˜�ϰmƛ᧚�7�
�e^?rQ��Jg�.J���C�{y��]�Y���'�{r{+l�=i�r*:;�,G=���¯�{�y�|�
�z���?`�U���1�9%�u�qֳ��?@�5�=*E��i��:XZ5��?�I�l�q�29Lp�r�'��o�//ЗU��"c-`�X\����n��-J���L��rL'}�b��<2����!��+��O=���ԙaňƩ�p���b<q_[F��o=�h���D���9�_�E�����\����}���f�ؔ�8�~�3�1K��N��V?�W��l	�&�ҖW��+ݤ����zhe��k�%����L,����!�cWN{�L#g��@I�-5Vv����̬oo�v=n�T�g8cw��ȤάRc�o��8�C|���X�<ݱ�d��u���*���Qp���������v�q����aOg����KEY�Tߩ����{2l�����>u=�ËZclLp����s"/�_�b:��p�n��;}~�qP�]�6�����y�d��ڬ,�WS���Y++"	Tٽ��k2��5���u_Lp���b�=gx{K�%k�a}>��qt�W�a���Cn#��	ʺ(J��_o�1��#5�d��c�VmU��k�,��z5� �_Ӣ	��ח����Bw'�aX#�����5q��LP�����v���ﭻsNZk�~�6��:��}��1��)H�z�f��lh.����Ny��ͩ���Uҷ5F��F&�ѵ����<Z���g��Mʎ�k�={s-~�#�p�i��rvب�5ې��+F��ˬ�O<��1Ռt���'"�}��f�)��І���8>w���Ǻv+Ӟ����1EĿ֖F��z`���(�+<�X����+���y��n�67�:8��f����-ʐ}�Μ!�2p:o�kZY,� A�lՅ�jD���G��t���e(����xu�T��E���,^7� �xY��Ì,	2���y����͋�aw��h��]Ѣ:��X�=GhU�1��8Gy;����_7u�
\2փA���k�8ٴƕ7��S2�"�M��<ə&hXFnmt}�N�J^X�pu����P�T0�E�Z�cjE���wy%%��ƆB��{��k|�ň��W��ƪzk�:��f����iY1B�L��rǻo��s��"��^���B��%�b����r�@ђ��Mz:U1~)��٦��X�wP�����P1��\��|U�ø�[隭�λ�;��Q��J���a���F��K� ��R齛�WH�fN����fp��V�ov�j�6��#±n��A�FIpIy:�za�n{��|�]��#�E,�n{;G�R
��|�x
oN�G/�i�=(""�fh4��Y�� u��E]j����Q"�4Z9�;�n$}�>LW����k�}�R�eb�r��w��w��V&f�R����2v|{��G�k$]�j�xT��BC��>������]1?&�u��`u��x���Ԑo�g�z��a{ς�
��>��w3u���Lw>Up!e�үGwA����TK��%��U��.����&3#�9%��J@>���aɨ����e&ѽ*��:���n,b�PQ�ޭ����A�������rڲ�(��۾[��2�Mb��	��=�R?^#���ܚ�e�;��ͭ��R��<���ry�l
�Rd��Ñ̫w��b$5J�=�:A�I��3v�˕�z�t��S�B�ī��A[��՛'^�l�I^s
���u��+-�����F �7}X���Ld��P�ot&20����*�	ࣴ?���O�Y��n\�P�����E$�w���c�Av�7J[ef���P��1�H*�������@���J��NV��=)Y��3���N�Q�[э��^Y�p�|0鈞V�eOu���F�B�U{r���ItMԐ��f�����Ge�9)��܊jU^���2�kc=u��4�s)Y��-	)-�e_�I��".&�Z+�|˵q�vr��}�#��yw@�x���Q�w&c{��D%������a���]�U��IS��֜8N��/(�Ul��~t�-��cgޥ�.3�����`U��c��+gn+!hK;<#�Ve��;�n�^h�Fc��)��v�bxS��dly}�lyA#NT$H��n"�Ac�o���,�ɯR���j9cy�vL cX��Q[8�QlW�mKdÂ��]�kӊtP�`z���.4�ʯ��=A�w]+J�����+���z��x��s�"���s�y,�^�/�jO4����~j����<*gA�@�"Խ�pr��|�F�����������T=��.���_�1�o���V6���j���Ꙑ�ⷋ�W������gK�:���sG,OE`��9��.�x��M�j�u��;�[6-�q��^�
��;j1B��I��^o �s���v;�a��WMA,�.`u./N��4�!�u��c�˩�+�L���s=s`��:W[��N���^q���8�����S�ў�^�26�P��w>��=���s64p)xw���L��@q�te>�v��*{n&�\��i��q;p���x��z�ɯd�>����9�V���S��]0F�r��>
���;��PS�{fs�ݟq97>!��P4�u(v�e�w%�s�7}��n.Bs1��&PWQ��Oo&dn�9�a,�|sZa�e=,̈ ��XiT6�Kr��7����(���W@[��jH�i����d��h��������s��x�'�MA���^�I�[Q|"���]1�ri���S��	�s(f�i���8����}�Vcp���"z�#R���U:�Zk=C�>y�l�\�m���j���x��Qך�h�e�}M��P�{��\�q���9��[~>�;�ҍ���Y��BN�`6�����՟?wu�̉����k��vb�v<�-M��Zc�;'���>���T�(-�`�=�8�vF\�K�n�H�ʭ�Ȋ;�D�"��H���jw�WC8�:���L��*�q��l!�J&���"o �X�R['s��:�7����Xm�d�o��3nM;�ϗA���'.n���Bk�ޅ����|і��`��Xb�Zgf
r�0�b_4�`&�����*���"z�w�5)�� ����U��r1AT�f�u���/�To���Ơ���y3���|L͗=�����ເ�,y8�1A���&�=)®+f;C�}*cR�J�9Z~�<�M�WWy˽��.Px��}mҕ�>��3K�0=�MȌ$��f;�2{�$�cO�6)� 1�.�p�'���f(w�33	�=�	̜�Yq�]�����T ��{�<�þ��Pur��Ҵ��'o��5�B�L�����f74��ġz'�&Ş�^��J�(yn���b�T�ǃ��Ư�)u�72H	i\�E���1��ݓ	�t�Y�q���c�8�TP�w��̎�E�r{�d�o����r��v,]����~��P�_/�\t�5s��|=|
2Nz� ^U�i��嫙CLʟYAi��Z5��R+O��V���ݵ�;f��WC͞�7����vT�!;�r�s�d�f���zcnp.�$ϝ�[A���`��K0�Q��	�
O��&7f�xO��]އ�4�n�����7,X�S�K�Z=�s���Y��@\��i͠��c;��>F��8ڎj3<3\w�_��};���	��[�z@Q�Y����S-�'[ٖ��,tt^U�p[��e���v���3-N!tv�Q:�($Y��q�WQ�c���w~ژ���H[:�v�n�74�i���;w�B8pK����Xq�s��\����'LD�7[q�{�p������&�j�՛���F,�8�	v+%����2�����i�/2� �{�Y.����t�w�:.���h�Lp~���%�����go�R[�=F��s���[�T9��~m]������Պ�hB&��J���P��Oh}�>�fF�3�x�`�؁T�:��x���g�:<�=���Z��}:���D,��+`���3:�B���٬r]S��U.ɾ&��΍�c���_{�����7���H��i����8P~�}�W�z�X��5J�zy;�cف���Py78�jf9�]_h���~a�I�������q�C��먨���]ʠ^�J՗��v�7�WEoF����v���cY5Z$Âb�\gJ\�ƥe�L�a	Sq�.5�m��u����rb�4��4,ddd�[ss�4Y{JW�7�Z�����N��[w.<�b9�v  ��[.?U��g�zjF��8
�^�\��]�uz�Y�N�p��n�>��G�ߜ���wk�g>���= ��O=	n"S���]f��X��|)�`���� ��ɰ�}��wO&Ub����d�����K��Ϋԗ)�W��՝����gYR��Y��)I2W*���~��{h�k�Zے���p�^��*v�-�i�^����}��	�U��Tz�.��쾊Q�N+�u��Ε�p�P�ʧI��M��Ġ��YyoŹ7���LÃ�i�� �W��uL7Ȅ�y�
h�R�q���]�{B%B��oU��ufz�{�C{:as,i��N����_]���(ܭ�]C�^m�,���c�HkW�|�_Tw���*�G �d�HZ���B'
��^� D���Μ.��q�x_]a>��G��=�����}J���]�1/gf��3ݓ�=�P��u��o)Ln��{\R����!�#K7�6��� ��0o��|���)X��[r�u窺4D�z�,z�I�����L{��f�x�Go��beC�ȕq)&)����Ϯ��L�)V�{.%/B�<�såjމ}>b�-�=�l%I-�B�����Ԏ��cV��MH��Ys��"�����ڒ�Y�C�o!@������[�}}�Y���E��yX]=���R����(_y��m:������=���x�s" ��*�&zG	�Ψ\�Jf/���"gʦ�{��)U����\�s�2�g���ܓc�f�.���Q�_ni����\Q��}|������v�]��i��}s9�v18�1���LR�	WWe��5v�9eixi3\N�r �i-����e��)i�E�=*L@�Kw�۬�X�d�1���W(�0�����SZtK��u��wR+�j������=͌]��s����gt�;��+��O��.m]����� L�v��@ŬG���6���f��eF�Po9�&=X��DT�g-Exam��>p�V_R��9<��1�h$�s��F�WLg�b܊J�y��k|␳����0�b<|Bz�nB�ҍ�12��rĢgޡ�nET.��ͨ���ـ�=N���ZY�=�]<�r4j�atA��"�2]�{#�i�<6�י�SJ�P���@�Z�p�eF�A����M�6Gx�u�͜vf��+M�sިJ��O�f>SX��t�f�P��{��{���,���q���R�������= � �z�n}�R�v�ŉQ^��Rἃb��7�"��q�jӝq\���6�$��-ߍ���I/Rq%F�p>�T����E�&�u�?(qK܋�HP�Y�o3!�3��6��o�[8����lM����� L���Ӟ�,��%�>aP�*;�q/�/�7�(�o}����U3��4E|ԣ1m���Ω���*4��5^P]�i��ʙ�/� �E7ݹ�,�۲���xV��i�Jٌ�4��s�(j*�!Hs.1��q����a᫶ٕ���}W4��	̬Ŕ���6��m�W�gn�3˦�����k���lM9��f�c��E�����q}���賴�B�;�H��|���][`�\]M�KQ�^"\&�6�{��<6��O�xM����-]�_�����uFWvS�C�8�oT�1��(��o7�F��9�J{`�����_x}+nJ�h0�mG��P����ڵo���9��U�Р�bZ?c>�&���\�odD�����whǎ� q ���id�\��UܣM��T���H��= ��*M�h�=0��t	�\\t5�l]E�'t^�8~�>���	�SFš㪅�g@'0B�D��f�lO�8�)A�l�](�jI�;���e��γ4�#�G�e�k��v\ږ��;�U�GwA���j��=XX����}<c#fT��z���:���ת�$M��ۗ�l�jVT\z-��w��\i��qS��3�����p"�Ξ�H�Z^y=�&�B��U��e��|}i�h<�_w ��YΥ���t�P���+�t��}	ג6r/�渜�.ܿb t�E�b2@�ea�~;�۶-�*}�}�\���/u�\yМ��K��������&�x��:�T�ф�T���
��K��G�P���{��zj�W㴵��cEM;B��D�ﶼ����i�r(�X��G����	n��� ��h�0�eQ׋x7ݙ�T�y�)��w$c�4_�bd`�+�̴��X���Z;�ܾ�1)��ɢ�k����C4m�ZZ�����`:̘��(���Db� S��/f���{m��&���V����֒�� D;����͙ɥf>���_���/�!eqU��lY��gO>�O>ޠj��K�i9��)��iN�����;��{9Q8�g ����ucF0�2rH/a�v���aN����uf�b ��RD*0�8 �Y��P���h�/5Ⱥ�l>O.��Mɂ��25ŬL�WVJTK�=O�d�3��AY�H�uqG\� z�P����ek������9u-���l��I�8�mv���k����.�
�������.#(�e^ �]��Wm��+�i�΁'K�����v���i��+*���Zq����dR�ݬ��u&���K>$��Sbb���x���Ueѽa�x��¬�;�+iV(�J�r:���^q�v�nC\���[G9w4���ǵe^��X�9�H�;;h���`0�Zf]���/�ܽ=C���xv���r���ۊ�mMÕf!Y']�<�e�([N�'��W�u.V�N(��,zE�5�*P�׹�z�"Ƚt�,�:�j��t�J���6AU�f�A��g��rNO{���0]�\��f�67pC��7���F3�mK���S���י���F3NСswp��yH޸��0��� �i�q�����z9G��G��KE�|�\��`O����ɔʺ��$�5@�h:���V��}7��m�q�e��CV�����\�R��{�V����15L��B��|��&��q�X�S����
�Ѩ��W��[3��R�Vʺ�w'-�K�ƛۗR�ͫv�p���[�H�S�8
צ�Ohv�o1���V7�/�4AE3��R���tYӨ���(չ�����m
�U���4Wl��zW�!�:cF��fb�trVsHs�ܴ�s1~����)z�@s�#L��M�[B
��7��o\DO�+�����>�vY��,�:.o��y�ۘ�m���n������X�C���z��pf�&Z4^"�����7��8[eOm�1���\
�;a���M��Y� *I=J��Ϋ��W���Y�:Ⱦ+6\����gm!1u�4��|?,E�y�n�̭�Ԏ��{��G��� ��U�G���dB��.���y�^�Vz�]_	#�6N�9����n�I�;v:��w�O���`{�8�q;u>�"��Y>�>�#�C䇇�����eϓ�S.�`#�:;���3f����k����kk�&(pP�B�3Ew�*��7���Bj;w�R�[nw;������Ir]����1 WA��������3�>�J��Ęx)e�0�H��+5dP��<ɦ%4˪�N�UI�����u�]��1�ݠ'F����.%��y��$�f��v��b�c$B�qURE�WJ���Mc\�.�	WvXܭ�S4Q6���N,9N����/5��,b��{D�5
�+d���(IC���S[{¸�P01�^�z��G�ex�dz�<���%��k�5�����V�G`��61�h*/�P��{@�S,ȫ�ud�X�$�jK��sN\]`*s���x�i,��^1�'��܄h̞�C6=��~����W��	C��(�O|�}��+�݊L�]��G���;y�7w�&���[g/�jZ���|�%���)�u3���*�Ɋq�^�撑o|9yWb�jd �y�ag;z.�+mc����~P0�f���|&������[�/. X�醢�ﴤ�Y�c�/v۫m^v�ڿ��c�R�u-�������1S�'�EN�����6�;,p[�vAx��Ţ���\[:w,U�uM�����ޣ��T�C�2�����w�<�}U��`�S��>9�lÅ�!b��߲�,�J�7�:=M8v���7P�%T+����z"����+5����AQgyl�Ň�5�4;��\ikux=wO3��a�^��H�<+)gBx.��J��q8��b��J��VZB�Tj� Nv�W���S�c5Kf�5��;�������q�j� S���ط@�*���yX�r ʿ\�&L�f����#�a�cƄ��ōW�N~�8�PwJ�2�vj��j��	&-�4��C�8��U3h�Cb�o���#Ԭx����8�~έ�b�pV#�߸���';��D4��a���*�A�:'xjyA*���Ŧ�~*(,���4���y�äɘ�e�]��*�,��軨�6;��>� R�����ˇ."A7��sr�w��G���s�*U)��<�ľ�q0��FպΗ�pdH���v�#�0ؘٮ��:�ˡ26`P~ccj.��JX�����j����Ƙ���Ղl�ЯA��j%`�N ��~�'��y��V�tၙ'o��+�NÍ�1�h�/=���s �2 ��6�'�B�x��m�OmS�L�nԪŜ��>(����y��{Ʒ��$X,���=}>�Jl��"�[~7��O�}y���{<���N�a�3��Mp�l��l_�<$ .�����0��^!�Wq�j;dV5���G+��ٛ��ְ@��0�'��w�Zp�f�Uʴ�-nw��>w��{О(���w]���¶�b4炻�9G 2�6V0�&lt����5Om��b�jd�uFٺp���Md8��Fm��b��k�/����PY�[$��T�f�Kڑ0(>��w�{ta�| uU�*�9M���4��
����CEZbw��%�S*�=}MÛ����VC{=#�ΡE�2����󯾊��"~+�Wv�%g�T�[YtA�G���CWy��غ�
�����nX��S��dyT�?mq��8���tX��>6/�sHv	13�U�k	��"��ۃWi_Dه�3���n�{\���$�W�籂%�N��t��碄1ލW������xv���?�f~G0��|�]6��q�V�$٘�W��z;MK+"Ю�f��3<Fp�Q{��k�G�Z�8xe%U���C(oq�&�NƏ$����p�[�5D-���9Wb+ܾw�YR����pI��s�\�yb��~���]9��Vz������6a�SK;�o�ű�Za�i�j[����P� �ޡw�o���I[��Do�|�2�~��/EQ�ښ�-����q��'#��3؈�鍋�͑��˵K=�[����դ�:~-�o@�GC���G���q�~�k��+>�y��.�_͛���ч�)]�%��������Գe���]K�i�����i�6���c���i�X�q�tdL�P��<���X7~uC��hPoO	u�u�@B����a��OtȪ�
���F�K*�]��]9o���%vX�)��-�t�%L�#��r�I3�M�8Tᔚɵ���5���U��}�}*��]�(��C��wæ�3Gi�b���B�:��W�Au��)g'����
.Ri��v�>̿Tߒ8��;�0
�C���K.�X�+?b�sV�����~��޼������q�S���.{4iD�$��˵�������>NH�߰�g�=.�\�|2^�iY�Ļ��S�Av�����t:�r�Ҽ���z��x��c����{�l��x�B�ޞ5�3��ެ��?Z@�5��;�̢.;���@��zW��P�&�o]Z8�"�wJF_�_�t$U�����dI鮌�1��S��S�ط��h��Y��]Nl��OWG��x�����g<�}�ѻ�1�c��U@����3�I�?�[�47�$u
E>�~q�M��@�=�������[�?`����� ��J���ށ��p�7�?z��1�1 ·�k�\ [	�f�`=�T�z�oA,�*b
uj�^A���7z�M�@����2�,�o^β��@��;j%څq����e��Ż�2[���%:n�S��j���/�j�=nm���c;ޚ����\�S0�γ ����q��8;�k��6�멯��L��__ݛ=y��\=e@�|S�nxų<��+5N�:�f§���K�yK��~�"qzJ�+`�G:��ڍQa��ؤ`���MP�U�m�l����Ukj7�c/j-+U�K�b�^�X�D�DB�fH�6��R�Z����!�Oy,f4C�B=��O]��h��8̅�c֕���M�RJ�I��:oJv{;����?p���K����ZKR]{;�n�e�A��m�@����E���c':�A�[�9H���B�	N|O}x�	�}S��R�5{Q��[�
���X�ߦc:b�O0n��s������4���AEݴ�pp�v�ush��zj�w����pʁ���0�P���G#ʞEK�A���5S
-`r����O��>i�}�^�)�s>���W���{�i��:��*�Z�w�'>tv��55uN=֣�{�?o(�r߯����Z�lV��5����QY�ڀz+'��"�JظxX�FŴn]��X��J]^·�n�7��vE�4�=�^�+�Җ�NU��ثT��{\�LS9e.v�o5u�R������75�32�'(b��zA*2%�5�`�%�t�]l���:���s�C��P�&"����t_o.s-X�α]qY;�}��YP��4�w�n�i��:��L�*�xIؖ+��P��Fz����4xgÀx>��K�����Ե��2��=�M��?fg��Ю��h�������(B^�8�9���UɊ��pj �wnTɓ���>�5b�u�c�� ����c�-90��Ľ3*�&�T�,�S.��	�ec��kn(�����Q�yy��K��f�nLL���*���G#غҖVr�>�>�v��~�.|6�Yv����q��L�������J2�a�����\Vw^�����{�LT,E0t�͛Vg/��v� ��Nη�Y�=`����hsA3�����-����5Fa������^#P�.�f(�H;���*͐ˤ ��^���)�
.�bwp,u�J*��'x��9��Ǩ=7�U�z��	�(fu�wqj�Xz��L���]_*u�oz�֜��ժs0��:77~�4��ވ8�c�yJ�˝�wҳO1@h��f��LQI�
���"�
c&���*RO��!����q�M�%�V;��^���_m�촮�(F�_�E, �g�<�jf��&`�-�}0�;�����X&<����M�I\�Q~��U	lUkǢ�K���w�ݿ{+�R�3N̟42�+�t�#�K�sPVe(ο1��/3����ǂb�����4)<9�qݙٓ��=S~}M�7W�O#��Ʊ���z�1���u;<�B�g������\'zNJ���Ÿ�'o NRoJ�i�jl`���UN�[�P������ԓ{=���lK[^IL�f�zώ�\'�dՅ}����,/o�܃�P�(:;I���bE���X�a�Z&�؜����z`�����E�'�܊�s�3�o4�W���J���A��:�e�*H��\��Z��������?�ف��}Jynl�l��>du�gn�x_=U٨EJ~n�d��>%��՞<نm�;E�ܔN����e��gb�O\v�NεqY�vJ=eqY\�hk~�Sc�lFr�bME���YI9����V��"j��J���t%L�n��g��]KB�ul��?
�_ZI.*w#��hw쬲���Q�}1.���$l<H�󊷧k�'�Y4MT��Uy�wY.g2��H�EԘ�q�r}�����N�n����gB�"O�*�==�˪�q\�;sz������Y~���	܅qV"E�s/A�y�:v�3�\~�%�},���#>;
Q՗��qE�*��n��Ţ���/��/{�U��%c>��� ��ѹPpPsN��^/zq�1�y�g�3wo%� �RL��i�xF�]�p�W�����~���9������1o5�[c�O#��|��_|�ub��	x	�X�=�\�08���M��Vg���t82ŭ�\s�ta��e �T=6_�,�Q`I�;���υm����K�|=J��ty~>���f���\x��A^�ikf*Q���7F8__Z׶!r�[ɋu�\��Wz=�_&<:�[	p�t�њ�������V�SÙ�г:��f�
?����Df�%�O��({+�o� ���G��}�yͺ{�w�����������>�;��l�֯0�#�eIk2��~�U	:�����,��n��7dܾo���)��i�M�P"؋��y�W^��4�iކ���gԓU���|�.Ј���A{S�g,]�e���Sy�2�2GT���o�	��o:ξ�ⓊuY���yxm)���+ڔ�%.2���	դ�!�[��m��yt�K�܉��˄�Y��k5y�rD��3�U>}��+-9ta�52��w���-7�c�]�+��Nc�~��{a��m�5��wP�v}B����dɌ���`�JH��	u+��f��p�,�7Hg��[�{[J��W4��ژY�dd�,l����y!#�<4����u�>�n_�݂㡻�D{�C�N��l���Q�Y�,�%4��]�bU�e{�xƺ�"̥�I#X�c.OWc�~�W�r�{w"}#=�r�a}Zq�\vg}�X��"�՝G��>f�΁F�޻��=����oٕv�-��ÜԽw�ǒ�Eǫb��OyE�W{��DR5y���'-MU
�F�>F^]I�XPnYB3k'��D }p=m#iC�MX�W��Fe�+*��5(x�o�Q� ��Y����c�ȿyA�b{�;���,��k�IR�%���nZ�u�愖��Џ��q�{'��8,��^hv��3K��N��#2h]��-J��Y����N.g1�9m��n��n�	]��K�s�s��w��ʊ�d����v�Ȯ�X[8ݸu�\l7���յ�\�+O\ �^`�	wE����	�Qv����������y�|M�3.�q�v~��E���JK�O�xo-ׄW��x�eԱ#�bpk:��ȰD��s���ͼX��=at��ǞSU������D<���.��)ӃaFMfٳO�=y����:����;K��^5��J���0�a�T��߳�ʅ�#�����a��㍋�Ib�=�0��d��mD�Խ�M2z�� �*����4�Y�R�-����Pl�~�S��!�C�3ل@+���j�ENK��<гkJ�o<���5e+��_w_r��Ni	�8������g�5f�NnȢ���zWr��w7�Ų�A��LB�~�&���BW��B^��b��)t18��F�קg�ʦc	�y��*Qf&Ƚ�r�����;<���vub/]��OחK�4�=�2����Fk�B�ԉ�ٜ����T-���v�)�h�n�!
ѩA�Ś44��&v4���;;r�Y3-�4���f�h���, �S,�ⷲ��\OR�K�u���b����[�j-�iʷ��2⴩������U����p�M� �m>�I]���Z�Mt�����ښ��^/M����{^j}��,���dN�i�!X�ٲ����"Ϋ��w[�9	{[�w ��6�������5��{lJj�i��ֽ��BJ��e.b���K)AW��0&�]�����B�8��ɶ��kr��81���[t	]՛�N��b��5��Sg�X�E,~��7)h�Y\8ޣ{�*I�섫(�:�H�{���k�B��`� ݉�ߴ��[d�W��^.Fm���V��;���F�aMȵ_JDr+#4q����a/��C�6W=\mv�=��h]nwQ�-�̖*��|��s�������](�u�a��LU���ܻ[�;�P�d%�"a�1��t��5�Qk<Ɓ����7��^��2v�u´M�u�4#�<+��\��
�S���Y����V��$+���M�"@�p�=���b�:>�4gm�H�{)e,B��R�����õ���?�M�Z�6-ś�"8�bm��I�Gc�|'g��˒�ns�;v�R΍ݪ[�r2a�����������k�	̓��;-��h�����3E_�]�n���\&>*��]d��F�VL4���<4���L�T�{��"���M��X���.�+a,):�{&�ģ�L�E��|���8V�Cu�t����.wa��,F��i�ޮ�U��{�)���6��^��Y�2���J-Ee��w8�%�@FsV]��^vqW���:�]��Zv��8���X��LG|���4����y�J��_3as�@k}�9��Q��1j��2��Mv[ټ5R�PCF+�|-]f��fp�$��{���r��a��;urf���I�2���F욿�D�2x������
�c����Q�lt����GS�6�,��b3tS2��Yu��.A�G6����]�aJ�Kt]֎�'��������f*�;P,t���Lơ*�����]+7D�SRY�:�2�¶sz�o]ҫĉ��.�j�)}��:}��ޅ�X�i�솗ta�<��+�.v�P`�$���"�����dGn���w��^���ꢦ�V<��/��t��9�G��\�n���#�8VWU�����Q���`;y�Nq�U��<�uN[��ף��e��2��*�ꢟ%8�D�S�2 ׈��^���@O�K$��AX�������i���=� 7��R�{�m����I����&����o�۫�MGB	5v����y�f\ �<r�ӝm_S�]�Z���ݺ�l�VQw����3V��:<?�,h��8��W�J&�s=�\Kyq׍���~/N\�c�Ŷ�k�2��XSX^�h�J��N��\����s5n��e��T6�tD;2Md ቢ��c��ӟ�DDG֮����\�1�+ �}�mb���c��哏股Zm�����?E�Q�p#�4�=u�f�\!ےuZ�l��v�,�:�5�(+���?��Z�B�W�E�i��=�z��p�P}�r��}7���3�q�}A��n�:�6yj�A�Dp�Ot��{��\R���~ ��E�������J�:�+Ѿ���n��H���?�g^|���bk�>�%���|ŕ���_m@��xGa���{a�'f��MvuȾ�+f�.�����ö3+�eb�;Q�ko�j��G;<Ϝ����~����zFX�Ve�_��0c��Z���6�<=�e=�2���pRT�j�u&���m�k����W.��[��jI�{ٟ>�~�����N�W���YJ�8S���d�[��Ogs��W���`���=����ׂ���m�M�����)ݛ5T�����J۽\ol� ���zD-����v���	�������8_i�S�j7	����=�n�S��yʸK�q'$̢:p�v��y�͒��0��LR��@�G6��Q�-p�9�82A1!��͘���T�{�VZ����r�j>ی��+%t:��6��

��s%�z��ސ`9[)�'� .,g]=I9�tWo"��eq�YA�.uvح[��Z�WN�i;U�0uf���io�>��<ӑ�x?{:�g�n|�����v�W�gr���j����cۘt�"���4��e����l��m�xY�G���5L�kY;ںwY�gl�i�g#�As��`Xo��Rv����r�^��O�ǡ��o��� ߣ����[��Օ���[n�`�-:��x�f�����R1�K��N�ry�!�����J��zP���I�b�ǹ2���ڃ�ju�{�us��O^�K^� �e+"^e�A������x���=A�()��i�ӧ�K7�_Gz*�
<r��r�|�y}�`̔�I�(_���j
�X��5frr�\.��~;�X#����V�x��B�4f(�J�@�u Y�5�ؠ�Z:��	����Y����T���}anck��IMw�}g���py_�ԍ"�����Ϻ`r��7'#�Y�s���m7��6e[<�����l��
E�,BZ�E�yM��º�n�2u,���[��w(9�/A���ոb��K���J���(8��M<7sGq`哫Z�mwY���
���<��X��;��v��M��;�9F�*��x�{�wwk�,�i�n��}3z5=�x@͌O}��t�G�Ҽ���Q]� ���1��&�;<�W?��y���0߮�3�ՀHG����V(��Ld ������s�B����Sÿ
H!Թ�{�j,ýc����K��NF��S���r�g�5��K��*Ҝ��D9VqO��p*6Cf-�z�֘ύVp+1VsC�8���0�b��K���Y͖����R*p�ut`�י����.�.7B��V�D�0����s��������hn���J�߳�WtƘ��s�O����j�J;�'g��7�$]���'�.2}U[�°�v�àtK�u�1�o��[p�)�+���*�Q�D�(n����5V;��w^S�{=���:��}����BT�%M���O�5����T׻G�g���	��󋨽}�?��Fz=|3��M���u�=�؎�d��Ml���ڭ�킧�{��w������O��x�QU�C��u��W����ӵtSMj�Q䏿n��x��W%�Nwg��P������u�mq|��_l����%�:��M�X�b���0���:�x�]v�U���{�aww��Sr��fp��v�);�gȺ��յ��u����:���\4E�ª&6��r(�P�����~|/�3W�x�q�<�������g�z��Gձ�^X���GD\X���T��~�G�t���W��Ǿج92��cW/S�v�\��8�b�;��[*��2E�/�T�aN��t��OE2����G9G��pW��z�^�Tڛ/u���֧�������>�P�0�]]A�:�wj����`@�D(���o���0�B[ɿ0bq��̊����>C��W�w�Y6~\��MVZ�7��J#�N,Jg����x��!
1{��E?7{,S?R������v�)�C ��^�/>�}E��1!�q7�e���^{�	D��k�YY�c�����\a=1�5>it�wG��h���r�t��P�t�zⁿ7c Ƥq?��\U�SM���4,��&5�
}\���]!i��˒XU*Vu��s��0?�|�ڊX{7�u�9��曢�K��v��1�Ś�֮��4���-��p������7���W�/�K��a����7�hȴnb���ܭ��ظ��S� ����Q�VD̥�k@u�-��/Os�����/=㾲�n�ͩ�p����Mtϳ���n�馐�N��&=_(����<rd\�]�V���p4.q�����Q�{��@tI�q~���Eo�r���V���^��8��xM>���3�hKA4���z����3�P�r}{��
�q�����Ru��>�r��0B})�ެ�i�Ȝ+<B�B���>�Cܜ���3�5�j.�!�)ܛ��w7�w����W�\���w�r�bY�G��L��ow
��pC����]Ӧ�'=��O���.�v7�>��L���iz���Z�k�q���NI�=	P��'=X��q<��o��y�r��׽�R�ܼ4j��16�;ߺe��@AA�f��g7���R�������K��;hM���^Ƌ�OT\�X$����Y�ǲ�nc���l��@�q�>{�8_<w���"�d�/�1}s:�E�e���HN�.۽�+\��#��%Տc��g�*�jbMLع��1�eWP�j^]�e0�	w�O�.{c_u�(_]��T�>�Z��宓�\P�Oc������۠�����ø�u�Ƥw!�$�V�ژ5aT��;}��aƱ��gA�m9�z�����{�>��ll�MΡ{$�ұ�YP{}ѹx9���C�w�@�7������&��UE@G�9N.�+� �"]fT�Ύǁɑ��x����l[����NuV�>��
&�EE_l.����p����׼�RL�b�Qκ������{Kz�fY�B�省Dхuh��J��6�|���;�8�/n���R�1��黌ڲ�X�<{��mV�!D�N�R�Sx�]Il��l�F=+������'��u������jj%C�%���������&�\��<�'�X�?,��#�]�2b��Iy��^(�α�N�zk֟����D8��/����w��I��_T�}���g���y��~w]�k�K��|R�ex���_"s��	��$�7[�"}0/gD."�p�u\LǪ�z&fM�m,# �Uk�$u��J\���W�l���[sH/q��i�IJF؈
(��H���)p��o�س�s`Vga{��]����J�״z��ڲNQ�R��W9�3�-�8c:��Mm�t;k ���e��}�F�NQ�
D��������k�+�z�7��HW��<�pb2]�v���$;g�	�]�a)2Ϳ��+	���m�|+8�׷�;�N�E[�6���ܵ�E����Wf0b�D��**��;���f��G:�����X���YBkTc�P�)����\F�D�;T0�Umz�n�-i1���٭Z�X�2��^{��o��{p�ܣ�ں�k̡�׬'�ν�^���H��P��yf�t����vs����<��\�f.��v(Hv�{7'���������Ѭ�o����Onm�]�j����!�,�zUᆍ$&������W�uJ�����G=�����z��|{C���q\������~��aa3�}���{^�a�𸮍��P�3g`��S��e�~k]��la�xi�{��h0<����'����E�BJ�9�%��oZ��,�ܽ1�����
{�u�=^��'~$6<^2�6k����[,t�xr>'É�J��S�4<�5ݿ����}�t���������wN˅=�B���_X�촫5Y2ܛ}i���8�y�Eo\y�z�s�L^��E��;��a�ۖ93yN���lKO�Ud��A�[�՛��1*�����ՐKx�nMN d���sG@�W��C{{Zቻ� ��W��LZ�ƥ��
�3^��;&�NҔ�W'da��y��w�N��-{stN�������W����ԗ�x��v�T�:�(�5빺�HIz�ۥ�Tw�.��Tw�;:������ga�0�p=k�s�[��caݕ��+�����>���y{�o5g�l�Ū�$�B�[�8)����瓡��D����<�.3up�R�c0��>�^�Z�Th9��`���T=��3ry�w>WF��;=�=��P8}��&�o�;��]p���[���#�t��%��:���Q�g���8�>��۾��l�3�f��?'-�Z�}�d�o��9���\o�?�]�[�Uf{�7����n�%F�,��'A.�gGO�ѿ_K��"�܌�5�[�4]�3���Ի�c�&Ve�L۬������� ��ا�B�ڎ�&ǣ������2���oHN�P����;b'k�6�U�¦qե�`H�CH}ڸ����+�Y�X{;�V���}8��oU�n�Ɔ�k��š]��Ժ�t0�/yY��5˱��zS��f$T�鷂��L��^�7�]��s#ˉ�tr�E\�|��0�FV��W�Z��K0�綝q�$��/icǋ;~�yIA:�=�0�M_��Q10#-���ב�f�2X�瓣�$��\�_y�K���"`�X�3գ��j��xR��������sM%ӟfU���>�h��fB^��w�ih՞�VW�M��Y�udh�q��'Oz}r�U}�x_�� �l~����ÞT�>�m'�_��o��䍓���ϟ��sZm�O�+�{ַ�J��Q�lrq0Q���e��ڛ��w8\Q�WjV���/M��`
��Ū�$B�9�����'1�d��0�����
�Bj�,��wiB�&hÍ/��Y%E�нH㯖����_1�/箊�����}�/�Ҹ��&�?G4���n�7�
=�o���]���@W
�v���ڵ�nd�y֜;�pw`�4o=��}�U+n�W��LQ=Kz�}��r���>I�N�`��+���хt�A��$A�r��������oy�4i�CCS���K˱t��r���(�c�+piޙP�S�M^�p�(�ݻ�G2a��*|#�j\k.p�ê�:��Ԏ���Kp�ҽ�cU��]�� �b�K!]��s/�m<;��wo��#��Zk�n��&٭c0O9|�
�ĥ[�O��j}٣Fd{"�M˿��Gj�)�F-�Z���ͮ��8�]D0���c	�WxPݦf������ϝ���F}'k݋�$�>�%�J{��F�j����3�A�]�U�@����PlW�5�e���+.�����I;��{徸z�02am�w��� z����+���u�ϫ�ո�R>��e�l��d�+���q���xw����{�ڔ�s��TH�Z�97���g>H�a�fɋ��}�0�ȥ7�e��I������[�I����4�;��w��>=z=�y����z�tI�Uo���p� ����G,�rb�w���Վ:S{
��GNtW�ձ�Qo�gΥ��k{�q���n�K,z�Hb:3Sl�r�hl7T��xOVS*�n��W�LB��#�׬�/ђc��de�E����%�=5���B�39���W�s�ӧ���>�ҵ,d�G��[Z��
�mA�UK��F�Ze=��,Cj^�^&��m-19�Q��Q�ؿJ�\ɭ�nr���X/:�6/�Ϳ7����l��/<w��3Ժ��s�NȺ����߀|�\��_����ߎ��
(�<h�9��
 �$
�	ΰUE
@2UQE�����"��B"�?������?���~���/�������?���z���_����""��������?DDW��AZ�������G��O�}���"+����u�<��}z/s�������?��?N7Y�~�O�NQ,���Bt��R�⥈3�W���`+�0�3H(6�M�H���h��0eJ��%B�u�SI�0ʹ^`��z��ڢ�ɼ*��LX��Tf��g�� ��)���Q%���h��,��{V1��,�1S�e��z]!�q�WQk`���\��[�؃r�p[����Ms
���5�W�g2��:�+tXh���%J�d��J3]�
��*5D��*��싙����f'����*�J�W!��r�:hc�W���c�x��$ɩVZ���z�ܭ:��[/���J'�9��X'�ϟ��w�^t��{R�㊤̋+4�M�q�j�Ǫ�jc�!���l�s2�VFAM�
���v�_F�͜p�6�/���M�N�H��wٙG�mq����ǻ��k�� ��IsIhĹP��H�iX�-(j��6M�S���ܼ������r-��[-��/ DR��b*Ѵ�c�)b�w5XIG�EJ&�e;��e�ͣ�N��D���ӹ�N)��b8�e�W6��6�6�Z��Y�K4�#ݺ�d�����J�d�ok��Z��mlMLU�Uzơ��*٫1�<1+ǟ�2Јc�z���'1f!b�[wS1Ӣ�7��NK�T+/5�j��r����.�$㱹M޾�e�j�� �r���2{z�TЇB�ٜ��)�Fe�F\��m�m��R@�d��Q�է1�V0�h�sYTڱi�6Ψ�v��ԭ�I�Y�D���n�!($F��
��,/B�*0DUc7Q�U�mj�i�w��;�4�4J�*�F����u.SV�U9��ᑠ��K[�E�UvΊ����ksjδ1�It��`�Ul�z��xv�VU����EF���`4�9*��R�6�V�܄nmen<���m�U DUfB�d�LL����1h2�ڒKa�^M*)�`�[�v�T�5b���ޅL�hf�������@�aZP���ɕv]��n��6�蕐�͐��P�El���(^��%�`Q��:e��i��^'�^Nf���2z��� ��R����XwU7y�Yr��y{12g���D�w)�Z1�`�z���V��w�!�K�t�ћ�z��JpB�4bNL�O�a9!�.�ZIC�\N��z�܄�B�L���
B-�pa	�XQ0C)58��c"��B�I}�}�gr�Y�j�֪x�M�2�tbr�uN��\���ޚ�e��+���e��t�I)��A+!i-�j�Qvt�r�m^ha���͒�Mp0v��J=3ZAy������w�u�}�؊��*�J�2
����	�?�*��* J*�B��*�B�*�@��� 2�9�ȏ���A����/�ˬ����?���������ϑ��|?{�q���}�����_>����pc�;�^O��"+���=��!DDW<��M�""���{��?��ɬ:���l�7y��f�X��3��?���""�a��ɇ����=�7������DE}��͕��|OÛ�ã|��~�ξ""��� �o���u��=|�������s��o�w�""+���|E�p���e5��)�:7e� ?�r 	 r}� ��m�;����*�Ӝ7r�mκ �P]�J!@�����X�[�����C@f4\�sn�"!k+A�TV�Q( 4ԩ�&��J���FD�ma�i[1+Y��V���Q�m��j��J�A%%D�U*B�T&T(Q�(.         ( G]�R��ET!ٰ(  @  P)J	)s��(�٢�ha�� x{��@
�ݗ��C�҈.�  ��,@:���`����^�v�$�A�J�-�ۭ��O�K]tat��B��xtA@� ���� 	�]�����h���G{۷�.�b���g��[l�ws;�j�k�/�|ͫ���E�Э��w{����{:ʵ}�m��xwWo�{j����x�{٬�n��{ֺ�����'5�U-UE#�D1�Ϸ/{��z({u�k���wt�Z���W�ų'E��8�:��}Ǽz-]�z���zy�t�gs��t�����m���;�z��۠7���=r��ٺڞO��Z25�B�(&�*�}�����m�s=ܜSJU�+9Xq�gt�;y�Wy�9�ғ�k�gj;w��ӝ��vf]������ʹ�k�y�ow:�f��:�t�Y�{���՛�S�_FZ�tiD���;Y�ٛk�V�0��}�_;n�7��m��Н�{�^���p��{;w:��w�z⻸�]=�\������gc��}��گ�*���7n���_{s�J�1ٶ�Q����_o�I�^�\cZ�]���zڝm��};ϻ[�9�}ϻ��تݹ�M���`o����dw��]��kxǞ��{e���%��ܻW_w5}�zc��TIW[X�E�����[m��;ԋ�����������v�׶o8v�t�w\�o���{���w���'�mŻ�j���:�+��}��oZ�5���]{���:�_>�KRN�)J���Q�]����^e�}�y��o{U����S�[���{��צ����eUMk�c�)����']�Q�vǡ��v�m[�[��9��s�Љ֤�F�k+g�}zu˝��z^���N��}�x����]\z�]Mܹܫ�Ӷ;�]:jmٜu�׾y�>[������>�C�ӭn����������.��� �kj�#�����^�{�]ڼ�s/C���{�'OVn��{��P��{��[Fn�+�l;�2�l+����>����ݗ������'��ΧwJP��w��5�e��S�	�T��� *~ф��H � 5=4�ET�MM=@�� ��RU@ � ��D�U*  &���de1�S������}��������M��Y~�z��r�������~G�]��Vۧ�}����!N��g�@�$$��I��P$		'�$$�!��!BI��$ HI1��$$��@��п���?���9��t��m�.���'�ZdtdƮ<���*r���m)5#B��O�T�t�ސ�ZJ�U:���E>�#)o�ח���#�nQ��0�{XA{l�UQVR4�a�cM;i�,��b�����j���V�3Va�jZl�^��d���%��ܰ�B��3I��̿�P�&�Ҳd`ȠА�U��Xtn��!8��L��Mn�_g=�cƁR��y!�����kv�'�d��i�$F5��+p0�xB�&���]aj��-f�I'K�Y�X3J:CW(Ĵ�������T7�^`Q��8D$��L3�	�7ѳPZ��a[�&��a���E���ի��{�D@X;�V!�M�RZ��$�;w��x�{Lƌb�Ƌ�(Tźo$�%wF`�Ej�h�yh�%���X��谐�@�*ţ�JC%1�G�+Yz�}������g[j�"�z���B� T�[JkY��j�j	�@�/MK�,��T0�h�I�MG��j,���������V��X���La�s^�d=���2�o�3<�̏;@x��$6�Y��v��θ_2[����������؞���Ɍ&]Ej��c(���Y���
�ē���U�6d��$ɤ��Е��A6d��u�0vCa�#Ϧ�4�̤�؟K�+�53.5F�H[#*���dii�e�x�꼬�E<q���6vcɱ�C�٢אnU�Qܭi�J�@BR�m����ф�66^�pYD��סяK0���l�LS��t=�F4�5���	��[�/�;������u����]��Hi�����n+�njUog�ǘں;)<��/n\9�%���)C���7�c��4���T1�VC̘=�(�@$�|�L�-�Ys/�B���m�T7�V]�eڪ�6��#�"Qp�B�P�x*D�Ecr���?3.t���˘�:�NXγ%e^=�3�GO,�q��	zwk5f�}j�;���8/h�a�t�Kq�sb������675�;$ũ�2��>��D:�q&��')F,b�PTGOU�i� �`���X��(��A�G����Xd��!�k59���s5�����ُn��z��F1T�� ݃v��,P��^f�n�ř���� b�(���@Q�^�n�9<׸e��n�6�*�Ř�~�#��PiJ���SrVΚ.��Ybn6�5B0 ��\4��ۨ�[����lx��f��O*6�)`˗�� UK,��F1�F�&��e���Ol�)�.匷ޣ3i`��X�K����G��FVU)0a�E!am:bz��6�Xw���-(p�ڊ-iHj�f��������u��;G�,��ex�íU��� �-ۛ�Ʃ���1�E��zva��^�Vɭ�O��@֛f�RVJβ�2��*A5�#HX��S�nL��V��No���7��i��f�s��{�C1��7@�t�bC�CEE�WT�5l
�����\d<��LRr�IĆ�C��x���4����$7�b>�X��ReI�C�10<���6�,6�',eb3vY5e��A`)$1��T=Ki!��i4&�Hu �1��A`k7�S��X²!�T���Lg�d�L�D�I���J��!�H_Rd1!R���$AHu!�R06��!�CiHy�����#�����F�J>y����hm|n�L
2��)f��7�H�N���6Ú����BNՓ�n�)���a��d�v��9Hݖja�7��k̢.(�R����VdG^@I����J�+j,	٣�T�5����6�"�eB�m�ʬ,L�"Ø�Y��`4�ܰ�ja%�;��5#5 ��Ek-��fN,�"����	L��fVlP��r��Z�	J@��)[r��I6n+�W\�5EYR�e�^f(&+$n�cT���%D�;�ER;�v�� ���� 'ěf��<��g�vsY.lVn䧖3TWv�Ј�m
��艭R�����%�/".o�Kn�/f�^�`�ь���PK�&�G=�ɶ�L�;�C�Y�HfQ��d_BdM�KT��f�����&�a��S@�#w!t�,=�w����,��ظ�f�6�K-�d7I�+te4��Gܕ� Eq�1�yZ��{TA7��&T��jAlFA[�#8�BI�dܕ�T*3YZ���p锶p����dJ���y��=7Y�ɷ���!-!ZM������'��1�Y��q�U:��`�Q`6��qe$E�h�q�ۑLI���l�yN����3��2�0�.�`������@pzbj1�҃�]`�.�;�*������-�͚]�f���n�f�n�٠.�=ۭv�R���t�:��;%2ᵏi��(M5tm��d�-�mURO%4s/\.�gs����� �Ki��A���Wwf��c�֓�v�"��V�ú�+Yf�svna	�
�GY@��JWVc�]�M�ɚi�&bu�N���FA�%��_$�˘�]�f�YaM5���ֈ�@t�Z�ͻ��d�]j"JT�:��t�k ��Û@���j��iѺ�&f�DD.�,�@m���ܻ��V�pa�m�(������ ���]�rf���k��-����j�ooS�JW������wKY�w�a�/4����˸���q���%�2L 8�đ�&�,�(�a��?n���u��S/]]��0��i�!a�m��dd�p�h,���ӡf��(�԰�mPǳ�A�t?:��40����ȁ9.�94�����^Cq �ZQT�´��m�	����b7�d����(1��Wy.Z�Pf�;���GV�8�)1�P�̎G�[!eK�����Q�񟅝 Xv(@����W�"ڎK��C!G@�m^X)�Җ
��N�4�&��&�n62��i�Ђ֩�6ˇm�ٷ��]w�9�f�!��YI���������Z"g]��\�u*�zf�2�T�����U=x�Z�p��N�t,fɍɢՇt��wX�ŕ����"�_":k1�ڊ@��TU;o�(躛K6�k�BM���;8�$���|͈���I�]�&���DwZSC9��7��.��{|�1�T��Sf:�����������)eLm��{V�YM�Ͳ����4ϖ�6fm�J�%bL �Rk�B������@h9$��f��o�X	��&��Z�<ZÑ�l.J*����hq�W��b�ڌώ+�NB�h|��LƄC0�B���9B74\�k5����n��>�4��$",8�~35�o��{�&1Ao5�VE�j!�n�H��E���2�ρG+*]��$��֨[ڱ�c
�G�L���C�RUiQ��a���� V�Xe�4)&���z�׵��QԢ,�DQ�۞ �n�uU��j� �O_�0� s41�cT%��� �V�8N%y��y)fcXN:0�e
xdHPy��BT]f��G�-�hEl$j�0�1�	[�"Zgq���F��RFH��?-�:˥GN�f�{0��<A.�d�T�Bd�U6���Uqܧ���)Qp�h��Ăш����!�-�LQ�RCN�m�v��pcV��,��`������Kr�6�1�E	�t�6�ͨ�m�{.Uܤ�` �!A�T�	:i�B۬��^h"�8���L����ń�Z�h$PN�wG+pU�m�f`�舞e���)�S�"���m�R�K&�Q��c/7H&�����5��ฬY���w���^\��v��I��I�~i�Ùdǖ
L7�~�H���oMv1У�Ǜ�#���ע���h1��ʽ����2j�6�P9,m
ِM�i!&�;Eʂ9��,��w��#�8�\z�^,��g.	-Xv�+�����d�ɔ��Í�H������3(/I4Um*/3a!4�]��F	�ڗW�2���&��e�U '̦Ɠ���D�y��@��d-�0]�౦�h;Ġ�	��21���ttc�r���g?K[P�j�2����&Z�wB�,I���^Ί&�ip�N��$�j��/�t+"V%6a�L��T�RL @���&ԊSu�CcVS9v�M&۽��al'Q2�e0t�v�q:5qad��^�%�!=���׌�u"ʐ��-|vk�v�¯,U��LMS�7�p�+1fJ��p�ݍ2�*|��Chւel{�5���i܀��3�ׯeG1-�-5`ۭ�d\"�Ĳ��Ù��{��}röޟ����r��WR�՗��U
q�[������`Ȇ��d�[��A[rU=�˴���ZUc,�)l5���e�;� 0���bS��,�.����m=gv�a�ݪ�6	V"'$Y6�@�R�u{w����k,���P3���>$�e�ed[5٠E˕e�7j�[0�G	{{Z�"Z;f�`��U��F��e�.�J��p�-���46^hkq���&�,��b7�Sܱ���F�4H�0U�[��s[����ܔ��D4&��X{)�T�cԞ�՚E�!�m����[��S�lM%Z�J���-���!��f�p*�fjR�2k
�{����:�n<fI0�n��!̅A`�bC�<�+x�(!iDY�aąc�_Y��}�Q�s�:[�h�f��)Jrt�s۷�Ă�C�]8�CBő���e C�!�s]i�op�i[2����Bכ(�K"G�mf�l��5���eBݢѦK�F��ɍSB��#��<�w�u6�j "���s�/;��b�d7��E��b�d֜�/!�*SF�[Q�QyDX�:Э" ��楖��\ay�m�"="D&�ʙ�iiq�wI��w,�G-0KEAg+�]խ�IAG%A�2m���΁��p6�I�r�ʼ�e�t��a�j
�¥�Ǖ��3A$���2$:��e"1��v"<�1d�����8֋�Z�w��(*$�j(X��U!Q�P��d:��n������ g�G�Y0;/�t��f�GTa)�y�dt�<�"��S��݌��������2(T���O]4.��m �ݿ�ᛯqH�`�[��x��hݐ����!��?�aK2�U.!�n�ҩ�(���8�F%0o`�;�{E���������&Yf�!uM��3K��orҙy��0��z5G�~p��mf&�9�NS�VP�.=E��k2S�l4b9Ң��2^D����,S��d�S��*\�!S�t�iɵ$��#Ck#Tc��T(���D��=u�l�%c�YIZ��xࡩ�f0UR)����Z��T�e��P�%�ճKת��+e-g+p\9j�nM�b�{-� 
�V�鲖���C*ر��IO�ͥ5f�Ӗ�e�����,��k�3U@%�+��xa�X"��n�7+i��^Q5X��Z��E(�j�7A��z��ZFnÆ�軦�*����ʙJ��-���т#2��gs�}�Q�5�#�[nnD�g
X���h��b-WPZ����-f�Z�t֡svjw*(V�P'�(TY�]�d�lV�nG���c*݆�1{"�����=@ނU(m�w��ޅP���]P�7[�$a�B���eJ�[��㱄��{�X�l&�j��E��Yx�#�j�@�aJ�⹹WJ�-T����KKWj:b�k'�۽���A+����r��x[��Qcn�e+Q<kF̤Q���r��[����5�bXP�nʲS��g[9�ٵE�_,�i��:Ѥ`�nRt���Q����e@R��nQȳ	��Ev%��.��A�"�\rl�ee F�F�8?fѵy�SXbh�t�f	e��d!�\�DV�m�,ܵw��Vl���U��#bT�T�vuܽP��(�U�k2=�c��D�b:ޫH�
��uu2���݆ط���IYv��F(dX�5fGx4ܽ�!�Te��'�8K�r��2=0,�͍����&<B֡7S�b��uv�4� a���6��̗m5��H����ɤ,����Kw�X ^l �b��~�D�1I�pD������cR��4A����k`���*�+�Qo��+*�4�[bb1n���P�#%���MZ[��7�m2$���,w��k��KudH����B�ո���J���]C/@�n+n��ÄƷ�@j�ZYkNSgn�(tQF�fAX[��[x�p��ރX��mC����Uܢ��6�Mj�Ê	El�]ǀJ��W�nj.$N�����{�:��$}$�����7�F�II#}$o������G�H�I�#}$�����7�F�H�I#�$o������7�H�I�#}$o����>�F�H�I�$}$��������o�H��]�����8au��)l[�>&.m��*�Kp���<<�y�Zq�E��w �:�)V��٫pY�)[��DJ�=�LoS��^oe����'����G�r�	E�@���Џ_47*+<�$깧�����YS�ê��Z;�.�h�̏{��ܑB��N��˗\c�:�u��-Uӹ�!�ߴsxhr-=��R�Z����p�����w�
��g[�
c�&{m��e�5��i2t��hJ�꽇9*X��X�G�����	�Ի�������a�f\ڦh�]�`��V3�{��sA�`0voQ� �����	� QnА�CAW�Xԛ��##+s���!f?d.�&AI�M�X֏H��rTQ�[���ܒ�J�fu��uz�L�;Z���ށ���r]}ցv�/���@�7�_fi�a���'F�V�U�0��e�>X���/��������NHR'�7g+���ה������Ӟ(�n�f�f�ՒvQ��������`�|�v�A]w�p���{��ݒ���.��D3Nv���:�	\ޅ�
��GT���Eb�L�5%9Yz�u���9�z�Kk;.�5Ta��Ζl�B�5s ��'L�2o����9OP�c�t=v#wk�]`�}�����|�vY���eVot�Y������U��s�pz0P�p����qr��ѭ;�{��?#d�@�j�L��������#|�a�}�uoI��D8ɯfe����t�j�������y��"2I�w��ό��2	UW3F�u�	�s�&9��m���3? ���o�ٝ���9�P����0C�٥�r��wgjת��o��s� C��`�֍��]I�I^��:�χ>ހ�%�3�ы�*�,q����]��U��;o��0h��7e��p��Q�s�:��]B=|��W=L-�+,��w�9�	�cm��H�{������|U���Y�:5��%qҭw�iu��1+�*��>WW��� ru##���缥������)MwI��s1��o]1Zɚ�8���<�C��d-�iX��9�����NL�9��;n*�kD�����+o9�U�/ZY`�d�ѹM�\5�"��w[���۲�ސdmH1���j��*4�[vlp�)m�+0tF��� <��n�]�m��!N�ʼy�)�C���dh�\�L{s��1��ng%�E�����&��}����%�Y׬b��L�cV���8����c�5[9��`���V8%���4�_)Ҷ�+��u̝8^#����Ǝ��[�Rgnp�N�4�+�6`y��)Υ�ƕ;�O����'��ѧ=��ӽ�!�aj�
��z��Tmi���ɫ57J���nPΫZ�-iz4�;1+1\���]!Y-Y��;��q�6H��zك7/h�)�,�H��a�r	{ĳ����T���,^�{�>����o��;(A�f������F7��tYg�[��QY*�w@G8Ǻ����I4���� �F!K�����V6A"�[?h=W&>53QWK���y����a�.���y�KK�7�H`���e���kו"ĉ�u�X/8���m�Y�V��o�dtEv�_)������<�.'3)u���d�8Ď���ˌN�������ʵa�N�����}�w^؛���hů����3���%������љ$����r�q�]\�X������O�&��X�&�K��C�OH�F�7�� �"�jRnY�auժ�Զ��s�-��+̼��;/�I�I�6�F=[��=GD��̭�$��0��Vi����թѷR���eM�k���Y.*�m�±���9dq}�����J�+�]%����H�ۅ7���V�y�5gFE�n�.E��U��f���9�]���
U�Ǚ��LBH�U�K�H�b�ݬ��
���)�6Χ����X�:D*>�S��St��*֗�c;�gqҠ�H�^T���Yvؾ�7��Lf;{
��M����Ev��"I:Cxv�ؐ%�SQ�U����<��2`����Лmk5"��)W]ŋ@�b�D���6w�7]*��ڜ��CRVڝ�H�����m��Y�i!K�,�&�K�e7�1�.��K���Tm��[�B��s����`�;�W:����\�\�p�YnX���p��ߞ>����"1֬z�ӄ"
s��;�#hg\�I�ކ��E�U�y��x�{O:����=��	]�W�t�Y�o�Y�ݦ�����]���%�O�����BqSȷ��v��DP�#����=.˦��nv!�˹`���SUu[}�������+�r�d��}{�b�[�Q2ru6��hZ���Ef<��ٳEfT���L8�u��-�x{Y���QW30^�٦����9�jq#$j�x�j=F)�n�&�����2{c�ZL��pih�;J�Oz�Yu%�L�(�iR���>�uH��w��,wp�oK�V�W�A�2���3vԣ����x�Z���p�hy;2�nA�O1򰳣���Ɇ�C����%[�v
���{��)�j�K �vβ��S��˻�Z�tf�hU�-���9n�]) �O�D:b�bQ�'P��d�b��B�cwJ���VD ����,F�1N_���1?f��6�����7�Z����BT�ghɼ���/d��{��ϴ��qs�:󐃪�D�cp��W)�U��eb�fNLB�+�a;|�]�a��Vr��	Y���6=�I��f�b�!gM�������椪�$͠��XY��<M�yg����]a��Ls���S�Ǜ/z�W]l��9�n�
n����W�)W��g�۾�GU�[+��j���T+����0u]ג&s�:��������j����o���Վ�Ep=�'l���N#XӊdЖٸ�Ӿ�w�e(BX%���ۻ�3nP�ڜ;5�����˗x-?b��d��jo7i�����yZ�.��*p#�$�.nw^�d�H� >���g��<p�w�[�X��l6�8��M4��q��Ye<�,�l�O+ �ڃ.�3�3H��[)��jƮEV�S{n�5�U.\��|�xj�)\� x&��jo>�ۼE�GH<�̲�;�N�5Q+�JۘV�h5�6�5�\�ѯE]�wǋ.ܾ�v�)p�ݷG��.��۬��,�Aȣ��G	w*f��&Ɗ�
��K��[���v� �{o]�xk���s�U�m�Fg���{m��̛6ZL��fN�d�ݴ�;٥5�u�OR�1��c��f�r�2�5Lt���
t�f�ŋ�a�E��p�HB\v�]�3[8�0E�9�on��gm8���h�[yd�Pr�놞εam�z�uu�,W�nku���<�i����L��W{��9�bV1�;�<c3S�J��ɠ��8slD�Yns�G��7�/����S����0����^9G�g�$mo<�3F��%�f:�.��w�q�PΚ��@8,������7����N0��z�woag�$�Ԃ�ъ�����v�d��tx�ri��5w#z�Vfh���0Ŵ���h�ւn�\԰��|����1�:j$�(���N�5g8�I�Ļ�i��Ig5�sy7:����wtq�S���-��M�|����2�+�gk�C�������9����*���^�{�.{�`�� �ۼ���[|�w=�3���ʣ�y�����O>��3�̣��
?")���v�q�o�.�{ε�V{]��	�ve���hP��+�w�gB�/�f�������UwqU��(2�^����n��yJ��_i�yV�wgE5E��zH�ޝv�k�b-��d��%���l�Zխ�ye�z;h������1+]W��nN̙��#`���W�9�%��Fq��Z�d�S�o)P9o���Qtkt�t,vh��I�Y�w�����ؾ�ǆ�����3���S�R���r�㙛j)d��"`vM];4�P�4t�D5���GF��%]󋒅hz�N�]$y�w���kK�>��M̨+7���˙�E��C\D'�K`�}��}҂m��^-�/~3��tۡ2u޻�/���oƚ��w7�s;�GY�Z��*�&& �l�<m�ae�wui�[���)f�b��Y�X�`�n�l@��*P|��K�����gdI���^xەY�nW'��ݶ ��˹ٸ�r[W� iI��:K
���-�'�j���*K�k^!��g1њ�v���P�1v6��q�]�^�s��4zi�\ƭ#���R���sU.�����ˎ���x;�F�*پ�Nʂ�<�X=��k��a��������c1f��F2⳺��C���J�^�ئ�bb�� �('��jٵ�|��r��R�i�B��e5L�Ꮸ�)�R�3a�3��&k�\?<�c�ov8��\��qG�z��꽙�;=�$���]��,3�Β��8����0��o�}*������& �;HX�Z��I��fk��������]�]��n�o�ӗu��%0���M��8%m<�@v7:�l��W�h���!JX]�&��r�˗;�c-t0Yn�B�j��Vy�r�]�+W�=-qM���6>��.5ڭwe���5�e�X��o9�o�h��܍��*S�5��nf���W+<��])>E��n���&{&�6凷8oAa]ٯj�]�7�pr�v�).�E����yJ�!����	��#��r�e�i�,�fj�+e;���Xc�-��������`E���]m`��e�,�w���{���B6SS7e��NM�iI��]��ǣ�G��B.L*���+�أ��F��2�Uc2	��(����(-�����{*�+�:9�,m��ӺL�C1*NM-)d�u�oj���*�2�յ��<�=K<w�#5�bpd��P��.SI��T��8��1��{-=2�څs�<	�\�ϙ��_Do���Ce���]7Єr�J�fd�������oq���,4{�����#9Ɔ�V�70�Ҕ���J�7���qr����uv����]�~u��a��#��*��<��Fr9q��2��qG
-W�I�\
�zz82�ug.c�Z̢t��dt�\�ҫR��7QmD���N�m_hw>wDNk�{������2%�f����y�`۾�T�w$q����6a��&�{9f�v�;�%�E�|��� 슻���̊�x����/z��z��&,"o���E͐mu��E;��R�'����{�fL$���ާ98+ �����^��w9�Q�g6��#gTM�^��H^�)k�$("�_h������-�Jy:n(+kAF�\�s�c�e+o��X&�KV~u{;���ڗܱY�b\��#y�O���2��ّ$���_u�p�h�AKm���,�BV��nD2K�R�v�|�v�M��%H�����G7c���!�0�.��C�t�=��m�g����e��P�o���{|s;x�m=�9E"{N�L7�&n�P�̫̜�B��d��뛾8.�۲l�iro��%�C偦3y��]�
��1������'f�`��qI�ʔ�tӄM[����v���wH�!��Ҝ�=O����w5�n�(��9mg��C��Ct�1��ur���[�E.�ޙ�&�Sy�o��Xs�V��muY�3U�2d���;3a]�uԫ�ܥ���U&�,n��Y���fp��말ZC?c���b�XY�}����p���t��w��T�3��k��m�{r�|��[0N7}�{4�S���39(�o*3���H��7��)�V��f��]���<Rt_>�v_��c���J8��0;#~�����塱q�#��u!�&�u2���Vmm�rk�����&�h4�y��Z�ζ��u]�-�ɪ�a^���w.*�ٙ���!�r��tj�I����s5�1�xn;8�f�����_r���s�w����&̍p�o`�<�C1fҖ_#]xQ]��iy�,��Q�C5v_ag"wsG�z�wv-���Íˠ���"�Ky��0�+��g�t��|�ŏ(�pE���{�g��-1ЮW�:�����82��{p��{��ZzuDJ�8��7�v-�u�/�V������vt�#O��[��q]!�| С������eh�ƶ79��!M*��<	Tʮ�S:�`%>��$o��Q�wZk�b�a2��2s����Ek�t��q��u�}�waݬ�rӾ�ҵZ�9ɍ�T�W����"XCn����)�Z�Y�f���t��Ns��8�u�Zk���vЮ6�<BwK�p���r<��"�R5���s�ܴ�0�V�枰�Et�WG��L��OZ��.��Xj�V�ZVD�kGOՖ;^W݃�A��v�2�󃋷��!���iJ�����!U��v�=����-�-%H�'M��sTt��e�q*o=�Y}��Y\I=e�%,T%*�I�Èkz��i�sl'���ヶfd�&�VA�w0�w�n.�7+o/%�+m�[B���N��z��/�o��Q�9��!-��v������F>�R�)�����q�5��ܠ�`�k3�	 i�ʻ�k�J�j�CLəb�����/A@����T��:��w�i�+e����h'�:}bv��ͼp����d�;��[�@���h�Q�wr��ƽ�f�5S!trt��4�-��4��X���q#��Yw�S �px4S'��5��ݻ�1�J��ї\v�l�D���E�V2]<ZKz���;�L��ս�Q�/4��#E["0�i%][�BĶ�u6,�!����O᧺��_�9����7t+\7��}�_-�n�i�
�v�k�o&�P�uwd�[��>�i^��1E�E�[���w~v�ߞ9�ٽ����RB�����!$�O�$$ ?	'�(�� H���H�$�2�$!Y Cl�6�I>B m	��l$� LI'I�B`Hi�Ԅ
�:�� ��, V@��)?�I>@�B��SL4���'& (u���>��@��LB�04�a���&�(N$��5��o(�@P�`m���	� M��!:��&�$�0��i��N$�@�b_X,����b@6�cI8ŒJ��}g�I�� �C\����`,9���y��`N��Y&��i
�a�Rc �d �y�E�`,��*�� ,6±ް�q	�Xq�b�G�,�>Lg���J�é\����0�4��$�->I��d�Nn�$���H@<8�$�	'��0�ҤyaF
� Q`�I&��'���u$!�Qa�)�IN;�15�`���vⰄ18'�C}�u	�� q3+h)Xd �&�l���`N&z�@�N$W~�E Cw�f��NV�HO��Mu�nڒ@�1P �b�a���r���Xu�2 ^�Y쓩
HJ.�LW��>J��מ����I'����f�b�����@'��@1��A�/�)�6�mz� ��1_��L�}I�w'�	�yP�P�ub+ q��f�+jVot$*O	$&ب�"�$�f+�r�M����$&2.���7-`LgY����i!�I$�)�!�o�x�>d'o+$���@<��1�$=�@�q*�X �� |�8�L��Mؤ'3�{�B��=믵r������I��nI3(#$+ S���k$�P�����7���-��T��v�5���_Rb>��g�P%�}��M}�f��H���1��G��I>߰�{��$�l"�|�5�N�{ԓj��Ǚx����� o�����9ok��LF��턫���|�.�����
����#}p���a5���p�^sX���x-��k��^��sr���w�n�TyBkT�5�sD4�����<�1�t��[P^��Ӵ뼓��|�{�=��}r﷽�Z遙�{a���y�w6Ge�k�J-,�&d3|֤�뻐�@�P5�|���`�0�����X��u��9x�D�X�,�,�/Mo���aS��n��c�@u��˽kZ�Z�j}@s2A��oPM�=;�~@�����;�S��ޮ��4D���A�`q��!�k&9���x�}f�h}Lp\�`�h�{F�=�L�o/�0�k�{\��r�����wԜ@��h�Ѽ��������u&fG&��L���2M=߻�;��'|��yִJ��_�k5�vj�|�rI����v�s2O��&oh�܇�Ӑ����`��l�f�0�_��	�� 4�vz��sY�:��l�fZJ{�u�	���s	�����CW��\ւwT�sN�l34�C7�j9�$�����B��7����t}Iw�: ��]I�y�ۄ�)1�i��5p14�˙>w�oUN�����}���=��|�w���{��l�ާ��!̰w�@��86{�|�[&��$罚8��Y-S7�)�rLݐ���� ״�PѼ�HcS�'w�sasC�̲{3�s�l�h��@yd>θ�C�%�&���A`w����ɘNf��lyu�r�g}����	w�f�w��ڀ]�/5&{����;p��{D���o�=�N��50�'Y�́��wRfR�r�A���3ԟr��k��i&�@����-�7A;���+��0��g�4{dy��k�âk�r�>���`�чx�"ն����@�s��l�u� �7_"��)uٙ�������}�����+��s��\9T���JN䳻�6�,�r������\��ɴqUm�j�Ѭg]y�9M��o&9�t��xJ=x�4���.�X�D���v�>�"Wc����M&-L��2!�n�y�s
V�
,��t����Gd��q�- Ҋ���Uk7~N���hB���?��� 	�߻�������H�}&]钲w_M��E��#���x˾��^o3O����L}A��۷��;��'][�(��{��|��Kۻ�y��hpWdvX��ڮ;˞U��A�jV��S.6N@�vDi�WQ�Ph��f];C��ۦ$g����l'1�0M���b�=�&h��i�{�GkRl������g4�k*�>�l�������/Vwa�z��A�]lD�Zk�ʙ �l��K���N�(�s�u;�6�ӫߜ}�Z搻/Db�$m��da�nk�Në�<�WX�	��Y�o:���a��[�?����K�u�@)���p]s�:痄�:w[rN���z���z�9�vƻ-�b�aI���f=��x1�j�l�"�YǄ��GY6(�����|GBfZ�ô�<s%���S�$Bf�C��p��{+,
U�3e���M^����e��yel�ڳ�,4ŪO�˱O:	��V��n��C���~5,6�Ic\����8��ʚ�3c�v�Gn<�,_Z�gs�m�s�(h��		�cf�riN�+*>L��R���)�[ϥf�X:�(�](L�lѴ
��K�\���s�%�CV�'k{r��X�E��U#��k��5�ԯ� u��H�utk&�ks+�b���sl7ky���,�d��V2h/F�p!5F݇Hh�չ�u��$�'~��2�T�莰��O��ٳs)"�{���O�_M�{{�BB	�s|��o����L�x�um�0]�B���-h��y�<�v��T]��e�J�O���wgv��s8��kn��r��Ko�}����緮w�>׵�T���$�� 7�&�&�:����"��$��!���@�$6����a1���,�ޤ��4�
�}� �@�m `c	�&2X��`E H {��~�ޭ�)�ÏĂAiTv�`�*�VAb�2�Ȩ�E=iD�E# ���b��@�&$U�Lj���X��D���EB*���\b���`�1`!�����?Z(�3M�5�Y1�s��TUu�c"�c(�F",
o}�����EUV2(���A��[DAAG��$X*���h��`�"��a�<���b�֊���NYA��E�j ��?B~��M�\��
�q���a`�QEEF�D@В��0ES,�F?�0��T��'s��}�z_����qUX�P�ET�Jc*�h(�s\��ս�*�ƣ-(�����
�?���J*�Y/�dƢ"
���Ň����"��Xʢ����O}���"�IU#�QUr��m7�Eb�سT�
���;��(őUF��1UE�*�eo��hA!Q"?��e?4c�.�~qP��%�ATXxO^v+���xwx+H���A$�#���fy�ѡE
'ԩ������DUWHX����V�U*PDdU�ϲiƨ�UU�A�\~q1"��b�/�ϒ�)��ȱL�(ϵ�MZ��kz�RnϜ����q1O�a��AV9aTD`����YO4���E2��1-��F�̨����w��~��L����ȱQ�̨�Tee��G��t�A��w�E��ԕ�_�V��1]Z��g�N:�DE�|ԕ�h��TE����m��h����b���#m�l�UQ���(�,b"�����z���:J�%TkDs������޿{�������ߦۖm5��+�b��L�p��*咟w0;K�SA��TW+���EG���b��EE�eFz�h�2��-��q*J2>�Eբ�W�,\ﮦ��U^�&a��dRB_t@O�C���A��\�ݷ�X��{�e��LJ���4�F������J��J���2܊9J�ľަjX���Zr��mن��+5�����_��klX���U�X.�����<����꛴Ģ�UD�����6�MN���z�.{��C��%��IR�J�0 Ƕ�M�7�X����Y�Q�/ΰ��b���5��(�$�^l�@�>-��4�@����\EVm�)W��Bڃ�����ڈ�S���*������Ş}�ګ[��/WA�����V*��W�3%=�i'��kZЦ!O���{w;�֧aET�.�Sc�"�9�A���r�*ԥ��f�F5/��Yg��Ww0ҭ��۱D��~a�+��2���A({gGt�A�4� �S���F$��l�A�d�B��$��c�փ��k1S��t�5F�����N_��wz}���i����d��,A�sj�!�I'�Usƾ&����\盾s�����4���2�\nc��V	��t����>I��Ǻ��/�^Q*���Y��d���k�I��=�I�an��\�<w��^Y�F���J�����(D�e�|˜�륌̡�Gd�v�Xm7�۩8�_�q��wY���~��ц}�hDt�P�9r
ԿkZջ˖�&wx}ʏ��_�~5+�=~M�ꙛLykNkF��6��j�7��P�6ɖ��N�%1,A[p����s�w��_w���Q|�jy�]ewlM4d�R.������-,(�x�t��K����f?<¥���
j�W�*����bn�5������1ʥ������b8��f�QLˑ�ڄ�ҽս���X�îǰ�	)2�$�!V�e�(�|�E�\t�R譼u�=�C��[}�E]R��з���\��3��֋�)�4����Gn`[�~~Q3��,��]݋�^}^|������@�)��&��]@*�H"���kT(�B���ub��9D*�%�����3+/��l���2|�aI��0e2b "Q�en���*z��V=ɷ�^��Q��0��9 g�N�o.��oE�*#��k��¾��3��Q��[�G���%YT&���}�b.���X_��6�R�9��.U���$'C4�8��i@�͐��S�Y%U?���%#bH�v���$�QAD����4��V��*,��k5�b.��4y�4K��l����y����H?;��}�s%!ݏj(�B���)�G�uG�>��$ ������	+�7G��Q�w�c-/���~?Y�R��\y���I��_I^�g{|���Y��c趨h��D?S��}}��沙1����o�Q�k=ut�̄}~p�� Q������ !-X毛B�J@�	���0~j�~�/���Y�&ǲ��V~B�b�@��aAidQ��-�,IE$�$"���DE���td�͑D/m��T���y�r�y̩Qgo�D��� �	���n�j�yt�jMO�o��߶j�����b߭A.���^?2�KL��9o(�'u��iT��k�ݫS���\�l�f���9i:�����S���=شK�ܵHQy��M#�-�Y���v���E�դ5f�T�鄚a
����4�E�wm��N�d:��mHc�٥�$gk�����<`5��ǝ|Y��i3mB�=7��;����܄�`%K������|�p����x��eL=R���,��T]�!~i!
!|I@�T�-|��^^DG�e�%��B���\� ���*}I�Dev�����O� �$N[����rݿp�zh:��)���܆�O����da\�h��+�D���\#�K9� u�>��WR����lOc��H����q�C+�|����K�� ��֨S �>i�D�����0��Z"�cZ���!9'*�Pq��U�Ѓ��Ӟ7~=������f�c%�HK��>g�0�z�8���-S�@=L�0$u[��]�0�d�F�wf�ٻ����μ).�ۇ��I���A�<��"3���O7޾q�XB��cR ��A8�%���㔐� � |�()��_ 	�Z��Ӳ�:����͐4�	$����8~e �ʎ[	��?+Ms��qO��r����y�����d�<�<s�Z¢�TW�t-]V�w�qۜ=p1fQ\G�2Jƙ����SH���p�5��E�@�#�ڻ�i�nJJ��
D����AO��o֎z�18c���P�����G�b'�Ntp��*S�P�<~F~�e�鱉1����1�R��m
4[oO�s� V����}*�i��D������p���b� �|��GH������Ά�bdGh�w �L"$���lw�G˜���VH"F��HB��E�B8��t4~>~�NL��O�Cņ�%$�l�-�#a�����?}EW��[��ǩ��rhy{*w>1��ŏ1��?��z*�y���i��1򦮭��#=}�Q��ڞ>��b��6���qk�ZkAΗ�
(�$�N�n��V�����ԳG'g
�S*E�ʨ�T��pȿ^�g��k]Ϲ�-�e2�QR�%$���9(d�L�G��a��`s[�a�$���U�̫H�1W���s#(;��S�*�R���G��r)y�ɒ��!!��2J�h�&r�������ڢe ���H����Tަ�e~��5�-��s=�_���t<�7k~�L���5�#7������2�Q2�F�l��T�N�r������J	�i�;�t~D#Arl�����*y�;w��k�l������z[W|X���$VG�<h�
$�>>��t�C.��ô8}���|ד<�
���6���x/�H�>��{x%Zzss`i��}⋶�|� ����`j��؅�1�F��oA�?b�B���[��'s�E��˹��ǹ��Wot����Nj��jyH-�|��������H�A���~g6l۩<�0:	�\j��g���SC'r�	F1n�ޠ�PЕ�>p(�6u!H$~ECI��K���B��" �L=��H�Ǻ� `!|�uS�˧���@�6�q ]*C#�K�ޟ�s헖�W��eh/;u�ӨU|���$�l�OƠTM^�4{��m�0�q�8'�4p���`l|�7
����F�D<x�B(�u��h��Nz�$��I��s˽C��?iC˫��f^���E�����'�oM�3���kx�|ۅ��җ� "@��@խ0��}f�{��!��!��-��#���m����j�Ś��?�}�t�yy��O���;�4�����.8:�US:����8�RT�i��C�ұO{��m.5:�L�|��*+�MwSW��o�,o���4���2�A˺S�mU��]��-~d�?�N"�v�QAS��yU�ESL�"��F�$���a�B���� ���{ԍr#�
�zşyZo�?2[@�	�u
�"q,��&;�X����[��Y��U��B��a��W���]/�3��o��RG�$���'F+�.���R��M�!���k>7w��N��krFl���ػ-;���X)��t�C
�=�h[����������ŐO��XbS`��,�n�S��A����G�5�'.-���ơ���r��vmڊw�M5	��_��w�p��]Ⱓ{#�%�^b��N��'35o�9f����2���T6�B����5�^:�l�/����Y=ۧ��@������BA.��Ө"�x���K��0,f�K2KL����N�E}}�U:n����ܬ��*�{}�����>�y2Bܕ �N�Aa`F�YU\�L&Qx�|��S��|oo)CǱ�*��7�d��Osk����S�+�D]4ƈ�<��`7>�k���?1�	a�Ti</�Φ��������N~��{�k����}F]���wN"JH���j2�Yr����waV\B6K
�����5�=nq����e���nӫ�|a��G�W`����eV�O�<�4�7J�$l��|��^�[+B#m����A�������!�L��v��>K�}��ֳo�p���� i�޲>�'s\�{���}�H}�d���"��Ԑ$K�fH�%EQLX�6�Ġ��(���� ����!�|��H~՞�Nw�x�{;�>�?}dv�^o��Gvul9Pؽߔ�&��!Z�j�.n�\��bp���c�ܪ�U���⠜��꣭�59�*����v�w9�ٻ��n8��0�A���`�|嶾b���t~�@�ؙ>nܣ/��I�}����-���E=;�|}s|̻���/��Vm�Վ�]Rh��EĈ({,|
�>�ǲʗ�����w�h]���tq�E!uЃ����~��}�M���EQ������L��
I�Pؖ�6�� �<�p[:S�Fy D�P@�y�טa��3ʇ#d*<s}w����hY����B���gp(�'�[�	H�+�����c"#�?�����e`E�Th��oz]Bh"��n.��Y=&w,�����*���ȑ��?��6��6��N����n�eWɥ,S�l]�<� PB#k�����g�Χ�ʯ&wH���<�z2$)%��W�*nueh���������2�	l�PK�SɐD�$�}|n��J֥ŵ��f�F�1��M�C"�Z2���~�7�e.���1�C��Sg�G�ʫ��!��� .���v����6J����G
�.�g��t
��:j�8z<?#D�cb���T�C5 	e+2�N�ws:�)^��c̖���:>}�=5�������A7��x_Đ����֜s6�o�>�cK�?�u㫽�	��fվc�#�������}T�7;z´H��;NȻ��ĤE�m2��;-�Ly](�$�YD�7�K�>�]���(̼����f���!���Hj�p$���� ~�@������#%�_��$&�L��=���ׯ߿s�g����_g"�/['7�o
���WN�G���Rk(j��q���%���vp�윝�e�<6���2�I�g�Dj;�����n��JK��J�g�GY1u��K�����#���i�<�=I�G��-�- |>꒛	�i�`�&��`'ʵC�\"�3���5�5�����z]iFx(�Ps
ea@��C5�j>�e!����* �8�r!�Ķ5��i�B��Q1�7�P��/�]V}�1cz/���">����TF�.^�a�ϴ�x�ۚ|<*eË�@	Gܷ�Dn� eRFf�k�(x��.=����"�s������?CLc"�"2:;�i^��Hq^9B|ou�1�0�oa��oҟu��8/lε�0����a��]�,y0�m�c��:a.��e�~�U&Y5oH����;/����K�6E��+�]s��J�|��I�޶�0υM�k���l��n��׻��=�ޤ$�xy����_@}�a��՗���f��U��$ނ	��"X{m�[i��i�P�h�t���.�b5{��`6L�
��_~�=�
���#v�����~�D����M�T�_���4�N{���@�M���i~r|��Q�L	�|gR���Z��f�Ww���S��?{՚�|�0�$�Z^q�w��A�΂AR�V�K�A}�BѮ5����G	�g�yw�U?mo����D�8��#�NZzA߯���ӯfq}��8	�zB����� ����Z7{�z�y����65V޵����-jޜ믾W��y��<��>HJg�y
0m��X�R90����~��O{~�t���yV�m=�mx��[������{���#6wQ}O�����~P�Xv��=�<�s��eZt䲵����7v��HU��S�������æ�xf�_ޑ7���D�ʹ�:Y�>�X���B�B�
���L�h�_+�@�|��.��|�\���8��@�徦��J��(��|z�eyT1qc gw6S(���U��PF�m4��b�u�_$.���-/U�M߻�{���9~��_�~��-�uv��s[��\K����wO@���yVڒ;XgS&�WY$n���扺�*�u�ߠ�傡6���e�i�aK���:�U��y]���L��r�ѣ-8J^Q���t���a|�N���;�M;oО��י��Q:g	L;7�>E�+Y���:�¼������A�$�����v��p������D;K$���vC��F█���=)���9U��~U#�s���z�f�>}[ �U�t}兆o�w���^B'Il|b�'(�'22�*��&ӽ;$�iFu��B�M+��l%��m=,	tH�ҺG��3�鱰4O\�|R��
��Ib}�f���n�ٷ&������P�}ѹ��+��|hZ�O$EgH�	��
��N��!��3ܵJ(�nE��_���w��j���vD��e�CP���II�|߄=�X�-ci�'�<4;��}��K��繿ˬ��p�o�ύ��sN�޷���� k�̙l����k��������o���9IK�k��(D�˷�����#'xKl�	�QL�pS[�³pp)C!�u�jlV9�,�`8y�/��+/O3�]6��*�B��d���ٱ�T��BJ���=Uk��]}��Pʘ�"y�!��{<�~��]�!�z�Q`�Ϻ<�a�̓�[vuЊn��bB���tc��մ�"*l��/�������S�4�'��$�� �:�ܾۭ�}X8��x<��c"ԡ�^�H$bPg��i���n�S`���M�`�l�~���Ȗ������|z��3��sg���}����"9$�d�8w��jZ}��B��wk�������	e����-�x��d��^8kP�S�S�hm�UFos��%�2������8���u�aw�,3��)盛�~���Nj�e��<��k�>�π�Ju&S�����x��&���Ly�şHa�*՚�����?�h{�ڸ��a�(�[���gب���KDG"�v�F��Sx�CPC1(m��hi���{s9V*/������HnC>�s�z:�,?&�Z�������K�`t��ǂ���'�-9So�=�a�u{S��E��B����C�v!�����o���
,�dE}�7fw6i�0������u�}��ӧ'U�ѯ��y�C-���R<���13�|{�U(A�y�d\���'��o��-o��PTZvQ^�Oy�o|�s8��b��:�1�  �-��?y��#wVqW�����\��֏
]��C@�:�RX�"��:�XG2�wSsD��?Kkt噵ZcݷGMJ-B��*Y4��<�xo����u+�b��%�W����x�`�hJ�D�D�9�n��˽o7��a�9$���pښ�te�p�o -�[;j�UW���Ai1�<W���o�85�p����糺cXO��;��%��u"�o�OE:�#�s�yw=YΠ��)$\k|��y�8(M��Nf��?h��HN����7����s�VA�ƙP[#��vyUQ&�:���h���o6!u�g��'Ɋ$T��I�:ֿuY��z(�{���D�ZÈ�B�g=���]�~�,nB{'
^ͲHfl�;su������w9+��~K۪�fM?9����<n�΍ �_miv���+S�pY=�Y��y5�*���B�[3�)��?�H�������7�?fk�}����jBI��������;@�'��陸K�"���I5P7A�A/tg�o���`�ͧ�"O:���g���C2�T�����X֊��p�ǵ���8��{��y�5�ϵ.�_��|��s��ن�v�-ABuϧF��A�Y/�=wuXyN5mվ��� ���}B����EQ��}m�i���6�$n1{%`l�͛w��	�>�v\�u�M���#�C3r� |��+VbG�VM��SA�Q�DSF/�|+~�Z>��.�_�=sTw(Վ1����m���yE�j��t��C�.g���dI�B�s��뻏;a��T��Vv�œ=rNJP��J�6Vv�Kl����<��1�R�c�WǷ��3�L� ��K,�o1n��*T/w���C�M�'6�1l���L��1�� ��M �sN�ff�0�V;���Gh�C�$�+v�?�/��Ec������4G��B��.j߼�Ǵ��Q_���\U�+<��]����8r۩C_���6��dl+d��{��.�]34h,q�uoi�2���{K۾d�{��cE�����A
a�ZՃ�eE�Q_��P)�ᘖ��߃�U���q|��eZ��":��E��潻����XL��������M�6�l���7��뺆���݉�w�5�K�i�[�6o]��Bp�an�̢e&!��MY���SG�P'N�$	��a���p�`�}	'��'ِ�%�m��U�4��:��z��u�,	$e���Y�z�:Kt��#��ǥ��f]gA�l�����V���;�Yu��:��b�OS"VN2U�ي�ک���gK��L��اk\�.�/)cɽ��
����ZT皎��l��<��;z�y�̲��r�cc��}���"[��oY�N���{�tnA:�I��B�򅓪��8�c�:b�XSWT[��j)�{�Io�篤�s��93F�[s�٫��;�C��kѿM��z�z�jthAq>��X�Ŷ�.�X��9����l��k�����2�U[��S'�.�j��(�}�E��v��h��'s@��Ĉ��wk��z�4�hes����ԍ�WC��̴�"�~�ΰ��!�g�|�D�ر�P�7�Q���>Z���N�M"�,w��h�]�	s�^M��F�霈O�g�N�9�Ӿ�.��U�IܞU�zi�+..������IQ�z�6�p��& 5��2i�:�(����d�:�̓�I<�#����X�T�$��'i����wf�6��mJ%��T���Wj���NVe�Kw_*�o��q77�a��f!�Z�����:�ݣDAw��Od�Nk!��A��x���w��3�֜��Su2����)c[�7�����f�t���\�n�̪�\]q��&U�Y�s����YY2}g�8�U;/<;\n��`ë�A�X;�U����V�|�lR``�����j�um���#aL���;���J,�6���	�]�p�G��._d ¤TΡجIٻ�H)���W�8,<�v	��7������vn�����ݲ���p�|�q�7�(�����z�9��^�vd�2�Y2��#�i���kb���$���rq���s��}�(��3U8��}J��z�.���bV�N����jw�s�X�~�-���唙a5�iʵ���BDss���3Т�NҜ�.cK����o��eI~����R����e�Rc+��CL�M& T1%Cz��?�}�a9�d�q5�3��LeC�?�4߷���i7ۉ�fD2��_�6�+/�連（����3}SSm��W�����']0yS��Z�����5�~�A:H������6��&�I����O�K��+9��v�2�>��M%B������8�x�4��o}w1�g��'���P��H���ە5Ǜ(3��������6�<��0N�4��()��~��>z��}G�!��0�ۤ���V(u6���,�eB��G�2i������7��C��C�w�ۤ�c�1�x_a6�~vɜ��Ӕ`8��|)�s��T����'|�ﾈ�M2�P��0�kZa��m�u�j_묲Lt!���I��|�~̚B����G���M�'�g�J�B�3��w�����A2_��䕋6�N��̼���������g�u*�C�6�T_�c��'���&���1<3hkVv��h���+�M���~�6��S��|���&�9h��i'Y\M����֘�#E"EH�3�8
i����O�b6ݯ��돲ڡ����G�>�p�#�40��(�5C��ĝq9�d���K���xg�/o\v��n���=�:��eH����1&�L0�B���bs��&%z�M~޴i �j���6�Y�K~�a�|���L�H�=#Z������{��T����¥J�E�<!��ݛf2V��࿞�~�B�&%G��G���'�m�߹���
x��a]�M��쁌u�<�f��~gڰ��g�'�q���`"0��￯���/�?s�9���٭����+�~�{vH���q�v�����v����6Ņn������T����$�}l�PӯY9��<�j޸���B��X���
N!�a^�OkYAG�,�DL"$B~s����rr�3�k�߬��Z����{�6�+<�v����
�y?I7��x~M��1ө$�]�i�U? o)14/�a�q+��yt�LLd�q'2�I���~���`�����{~v�LZR�	��>�n@��Y�-� � �`?�߿��zÌ/,�Xi�.!�c��?�t�y1���C�*�n�Q9ϰ���׉�~��}��j������i���?~�9��1��ӛ��N��E�'^���P��k��_�s�����y����h��(�a	�)yD?6���6<pm��Fn$d�/�3�b��8�i�h{�F�%��rN�Ps�ۮO7�Z��}��.�:u��y��x������<�~�A ��>��8���H	�Pr�=I�M~��Y�i?�sS�8��\p��"���LG�y���`�`)Rw����2�a��4�g��i#l�)�?��S�1�f�oh���z���￳���s�:��	��Y��|¢��'���ĜjGV�~����J��Oɶ�K���� i9�d���~�L	��WI���핇�~��¿����k�m���CL�ۭ6Mc���c
�$��4��"������w�h+0��V���&�Q&c���|��I���@�Ѕ�o���i�'�?��s}�C�@Dg

g�"��� �����۱���W�LMj���$���]����5����y�g]!즙�a��O"�I2�
0�¤� 9eG�C�㛢M�<`TNS\��!�?o{[#�Qa졂~Ok/��p�?���K��+��d ���>`�F�	�y��@�\I��LT6�jN3<���:���>C�ؒ�����Zp���g,ӯ�&�&�v��ֻ��&��c9����PƢ�2��p����>���s5�|�s�E���]`z'�����3��f�3i�0S�\O�O��`�LCt��� �����N!��g��WIf	+ĸ��Ѥ��#�B��T����P>O�c�w_D�z�֫�|�"=|ͱf3�pI���7��B� ��)���\t�N�����P�&~�����C�0���\g_�?��F-���k���)�P�m'�S���R
�?��d���]�??��1�㩉�I�bm�o�&���!�?�&�$��~`i+ɧ��*��3j�La��L~`UN��o�Ϳ%�%v�aS��o�7͆���i��i�
}}�ۑ����*ws|���r�=.�d �>w�Ç�8��}a׈n���[4 ���d4�5&!v���)��wSL�g�Ƴ����Xˊ��4������֛e��&�:�5����t�X���m��O������=��o8|H �I�z�?���~��q�~��h�'2�2fXh@RpB�j���M&j��~��d�hLEh�fz�!�LN:/��c60k�ߴC��L����}�b�IS�9���?_��?��tЅ�����wD�\��8Va�r
B�4".��)4�*|I}�<�*uҔ�更��fɵt�ѣ�V+�%*\֨+Vp�:fPT���I�͇H��)`KB�R@��=�f�S��,b�+�l�玊�v\��o��{�ݫ9�SUeW�j���@d#�;�q�3�|�_���2N��B҅s�c�m&8�Z�q�
����LC5���ݡ��r�ír��g��uM��&!�^��14���'�&}J&0�Lfe:�{?��ֿs�k�޾�q�B����M!�RGw��M "�{�1�H.r�3�~��o��q�����a����3���z��uۛ�����9�T��%�3lP��sI�J��*}������������]��� ��O�1����`������u�T��i��/��5���T���1�A`z\3p�h�,Y�Hm%~N06�͇���&�8ܠ�@�\@�~��>���e�!r{�>q��x�Z(�9(�����"�WJ�Om��$�z���c��*��0�aX�.@���|>NӾ�2���)m��y�}d]J�#ާ���ǁ�0DBB������W/{���k���˴
����E�������+��"|�DA��r�zǬEr9]��3�H+��k�5G�%�n��W7?T��_j��A�dӨ��~��p�>2�%C�� >�B���o��<+�{`���t��_yq�wJl1u:FfR��r�N�{y�ǫ�0��T�C��e�ꮑ<�����(�[���t���㙟��Gn��3,��GX�>�c���V(+����ӽ������A����~n��Z����A�s��OM�j��2¶w.g�K�p����~��1��H5>@���&7=7�H�h�!��8�0{�ɜ�ڤ*�O�����}����k���|K�8Lѐ	��/�ګ�C�,����g�?Xd~ۂj���;�������v|�|lZ�R��	P���:��f��</��*5i���l���wN�e�%fa!�|�z0�#��Ĩ��Qr�����8-�UܟN�w+4��]Ky�����\ȃ���yT{R����)hr���B#��Ҡ��f'�ԏz�Tt��8���5S<�}��.�Y��+8�!���I"f"�(�3�|>},�����U%U���)AbD�Dg9��"�M,��w⭃�G�u,��q�����������kug;U:o=4cu1.�UIRy���0�Ww�5�דCh��h��}� 	��g:/po�-�m�oi���~.���K����� +�|��uT�d��0�Ei�����3�.8��0��Y��lj��kн�J}� �]���e�9OH%#}�b��)S)��?)�v�$M���0�-��[�@T�5}�$�k�G�|a�O��9�c�KV���L<��p�l���C�L��\i�M]�N�u�8�Q��5�+��U�Mi+�JȜ�7�mO�y��~6���욧�K^�B�*�aM��癬����uk�,���I� /7�����h����r��~y�+�,8����mO�-'�Yc
�@b�s�A��T��~̛��"�ϚU�]�>1�
�&f�rQ>��Aλy\����Y��ݞ?,�^ۈެ�w�YY.X��}YQkj�Ͼ���؏��Ӓ�R��t:DX�����uU\*k�����ӏ������E��]��WX��������?T>��޺��gU}�_�(�A�W��ܠ�"HOa7hfF�k^$�9�K;G�Z�~�n�opѶ����_]�f��l���,ia.���^����=ǖs9.@���*�_f��{AxW2�Rfk�cx�pv���!�`%��٥>��IO/l+`oS��QU5���s�]�CR��N�w���̐�J|��/��~�Rx���J}���DDZD��]Y�{T�v!�<��)Mh�*:P�Ի���HG�Ot�TMR�]j�~���י�Ya����I�����A��'�Vj��ʡN��tb�_^��a!e�<���{
�S;{��!�G�W��� ��N�rUl{�]Ғ?M:h_�O_�����7�s�t�C�E]�Cݿ:4��%���\������^꧛h��8�\pS�K��⭤* �?A~�Ph�0���J�x�[����{ٯ6��5�&�f�o�����BB�]�&}:����(5v��&n�g���X�\����m�+����,��m͡D��z+]�N��m��vz�^'��(�QԸ���^�0�l:������ ī�d��+�"%�t��b131#���Nf�qmkÙ9�]�jHDv��_Dc	z�z�H�߽���un�F�,v�V��N*�fq�] F�2������92T˩-+����k�4ن��D}E�Y�n3jyȦ�|69_���`ڌ22��9Z�Bҥ77�}�cT�٠\�h�M���Ub:'x�^zI��_+a��w��,���$����Q��	���/�.�.lc�|魯��T�T��Gȫ?��:������AH��@p�7&�s��G���5t��5��R�#2Q=�e��D�ՉvD@�v�XL�5ӹ���P�c�%'!.��ξ�x�|�G3.a���Ҥ��!���{ͩ��r޾~��Y�nsѝM�\{�..�w���g�bmP��ڽ�Le�gz�7{ˏB��'���2���h��V��AY�9tA����e�뇞��׼WA�!�Z����T�71h$3��l��OŅ#������}����s((�|�E�ۑ�U["��}�����C5B�
i����ߍ��X��Q13��нB\k��S#����'M=�3a#NzߧN/��Z�x��ԤUt�YZ}a�|��%:��R�#�%�X�͚)E:A�Hz�ﺡ�h��o�p�O'Jv�'a@|I3T����ȸ"�j���z�K��6���q\|��Mg��ظ�N@?^�aʵy`L��M�jKԔ�\����:�HWW|�A�ne�
��1�t:��������o��6@㙯@��.���E���|��e~���8�ۘ9�;����^Ҁ�ڢj�R͛|��_�d�+�V$�Y��M#�xT}�,������]m��3��I_�|��j�|~|k2���w�{�F���F��[��+D��w���J�U|�9N�D�8`��2�(TT��FA�h&y��>JP1+�j\�ސ��ܝW�P|�$�M��\�b�ٗ��+�u���\��ݙ�x��49Z6
0��*=�3�=��%�m���~�_��FW���$��k&���k�]&Cu��
 MA"Ҵ�ta���W�j���_�e׽8c�s�8����ڪ���ͻ�����N�"�r���n�!�}J������'�i9�>���gD�l���T�Jiy���}�4�J	0�޾~�َ�]E�.|�}H�WEAvU\�V��4�\s|F]���a�f٘l�mae7�ܖs�^q�Ae���oJ��w�U7u~�7u쇏<^���aB ������DO�$�Ar�����r{���xr��3�2(����AU�.���b���Kg|;����i���N���잨�ER*,S����L���C�����N{?W�,��Fz�i�Q���0�tN�x�L�\���@�^V���'*B[Siu&�Lm$�g�-ܩY1�VGX�Z��q&Φ��6��#���m�Ro*0���iV��M9X����UT���a������*�]�`
7��{��Ɍ;=���;�U�N���f�ld�j�o�x��b�P�v:��'~#ʢ��KI��Ft����C����J��8qn��u�v�.`���ke�I͙p_��w�w�	NfH��_GuL��T�Q�p¯�KWYe!�!11�R��q9�j��rʟ����9AǗT�]�B�e�1LO�eݡ��~�M��ps\r��������^��Xx~���B�����fb�ju]^�=�ϬxH@`.�Š��m6�QiW��[_�j�Z�8O�}N�̓T���H���V�	�ͬ����?9<�D\����tf~(5Ld���י"�V��V~ 9.���m��f��f�nT� �e�>�n6�\By�y��#�*�HF�D�%���ޥ�>5�P����g��f�|"�m�]BS�e�j�^�s�w��V���.��[����o��͸{�7�fV�ul��.�{�H:�+���J���.��r�̚F��w���xC=�d���C��%�׫⇹�^�OoxO��o71ս�Wl��Q��%��`��g�s�����}��S��~�}�r�*OJa��;������ψ^��o|<u_D�0�Y2�Y3�)�5��1etw�쀢o;g���2N�M�R� ��f�|&��
�C�(�4`O��候��ճ��K�ܸ�i\1�J�yI6)fE�O��Φj�3�\���vI
@޽�󟵑�뻙*}O�ڻ�x���[�Q��~W閔��Y�	��ܦ�̼x)~"��1�D�F�N��==�G:����e
��"R�k�*A1�l�I��w�������M�y�VY�X��>� .{�ɔ�sc����8�A��P����s�{)t�S��֡�<&�	�K�]��{��dk&*&�}���{�%E���SBĔ���Q�t8d�K�#Ɋ��}U:=-��Tw��g�L��NM7�c���F�-����k��0{�j�ӭ�/b�AE	0W$iy�U�L��I�b��x��o§1Z>0��wn�n�e��ܹ���+��+$� >�rg�p�:edX�SS�/�-���#�^������'$l�챕�j'��"`T�(����Wg50_������BM�2��	���U���g<v�'c�����/���t|o�et"H �I��G���R����n�<C)�C����S<�dBH�1�NWGEQ�3�����g��k�}�e��}�p;�h�Wt;��^(������Ph���1�4��
�n�ؚ���mw�ʊ��.�b7��pQ��:\;2�3�ݘ�VGY��fI�_t0~sc[�t��պ��s~�x�������'4�I�젝�*�n��eN���d�}��*�%��U���EJ�*-�k��_*u�^���=��^�7�?]���G
z�_�ݼ����t*mR}�R��A�C<�v�,[��GJ6��%j��]#~��윆�Q��f(AGUUb~�Mg��$J�빊nP�Zy&0�z�@�6W�~�Y�������?Oӎ-]^�1��D�x.�A'�����U@����o)\�'�kB�tw�w�[�0�m��GUT����1&d��g@�D��YF�H!Sc&HK��Z��Pkm 7�$������|&����|�	K�}AU�>Ԯخ^�!]���~S��-x�.��xp)��� ��ؠ`�R"6�P-(쮍�.ޖ~�#��V��P��	D3�2jj���L�C:��:\��e՞�7"�(d.�SQʟ�G�G�r,�.A"�.�>")n�稫�q����g���>��%�5��]�r�x_����2�A�n��>ԡ�Ӵ`d9�&O*|}i�ИSs��<�Xv?���.[S�`��<-+mp��}���Ѫ�M�M�TP���<)U��W��G�����\d���{�=�^kch����/U�Ȩc�����T���*Bg賠����+�J+VghRA:�T�"R�^��ю���9@�.���^Gp���8Kz�~ޭ��f��h�}V%��-�����˄3U������B�T�*��2���J���kٻ��4ܓ-�ԃ�TvU1a�}y}�s�3�)��-P| ���|��X�]�k�d�&z�u7�^��h���ժf=�#��<�>���U�������WWR���}��.��l-s�bf�>�7T(�fP>��r�dm.��Y��}�yGjv�����p�]��A>쬡~�0�H�ܷ"E��H�x�:Ȼ��~�}�G�����o��[Q�F�VZk�dر߄��"�euK�UwG����c=�1�r��fF��yuڳ_zk�Lߗ�'�[ׇS�'��]��:��h�¢.��h���º�����ڦ���^g
�Ԝ��}�~�jw��X������hZ�6��G/Q2�s9��V�MR^-�?Fӎ�ҏ�f&N���đMI���F������-�5EzD��*���#ﾬ���P�J��zΏ�}��y����-��p���$��~�b��؟����I{����"�H��^8���ۿ���#G��הt���}wD�J2{yT���p!�q6�x�~WM���$�C�o-}%T(�"{�}�x��:�&�#ɯ�� ��>|9ϔ6��)nB(��>��̒�̊$�E��>ߺU�Zʒ�d�zg�}X��'��݈��0$l�f�Z'X���X�o�,O�j���D�$�+s�B���g*�˶)�ܭ�˙uqw�l8Ȯ{jK
J��oG�U7`������p&��9X?{%�&Ə����u�&�x6�)������_+���<�]wuњNzF�9K�sCx�h�L҄��f�[WOP�-�xq\_lǍo>��,Z�ɯ�����i��S@������άq�AXZ�p��#��aN���W#ʱeݓ>��	���}֔��/��7T�E�����1-�9tWS�ʝr���ȡ���'�\9������%�Uv��֨.���o�u�$�B������̺̏���_]�/�#�C
�j�u���dޕx1�f�NL����	;z]q`������;,<6��O	�b��ܭHm��;�j7�f�`�"���v�+��Z4k�]�\͞t�l0�Z�P'*cE�g;.�.7�M:���p)�wCJ˶�����y�G{Fp���d=07[� ;)̥K���1}��n�n�wZu���u�xumj�������^�nN��"��g)@c���kee�:���g�������n��N��v���$�I"�+���bU���X�5C�`�8 }�����v�M�PJ�s��Y�)
�ɗC�@�F|$WBb�>!�;{����{���Y��5����i]T�h���@$4&�%S�V�t��VF>���G]�7�V�50�ݓ���<8��i�oL�W3e��Y]ѭ�}DL=Iܶ#Ē0�7\����]V�U����0��e��f��>�ɸE�t������{�C}�nE�Q�Tus.Bڊ.��y��KdA���Cm$��腒�Aԙ�sl�;�{r*=�۲P��N�E�b�&n���Ҵ�Of��ѿ%��tm�I'wI#b{k�s�w�q��ǌ	���`PQQQ�{bW׆ˡ֩����4�7�������"�����R�0�Y�F�;�NP�-�A���E���7�����m�'+��{-u�u�ønq���S[e֒�[D�DZ�������
=��.���l�[����˙{9D1����NL�{�>�[]����=�w�1�D�|�e�Ԃ�.��HZ���R+o�.w��V�[�z� S�����/�"m���mP�kZ�^�%�M�!��1h��r��Y�GiM˺�[�xvS�,���v�om�8�_$s��P낖�h����kHL��I�c���P��W2�0{��-�w8��Gt�a
�%��.,�2X��?���?ы����v�v\x�^�Ѯ7�L+�z�����[
�`��m	��є/���ŅX6$�����ݰ�G'yXC5+x�;i��6�!&w"�]ؠӾj��G��akvm�hq��r�8j�X�����p��0�ݷ���g}2��v�z�10��3���\�_���7��_�sa'Yʅb;���JL4��,j�x�	kvS��ocb�-s���CuN���z��6l���)�Ф�K��gN5aJ
�9��qX�rQC�W>݉�[\���i���=nuZWvn��l���5sm�����Jח}c�k��� Ӭ��do�{�f�#}��z�*�Q�#�B��OF_IpAo�w�y�X����\�rgX���͝�I�qge'��jG�Y{d�����R��q����?�x��  V�g�D��i�G�DVEb�*���FWL�咕A��<�F驞�6$��1C�G��%�W�z#���H�K���6�MLD>,(�	|>����J�YӘ&�Vת�HR�E<.�+�J���%`�@���b��nH�$��OM���9��W\����>�/0JyU>sR ��J�][ÆN/<�8�@�$OEK��p�9�D�1:�'��鉹5��ڑjx��uW��p ��}Q�����<ݘh��q�u�ߏf4U�ļ�+���	�ݐ�5�cnqߴ�D���}3l~�$��<�LW!��T��qf�d��웮�%�T�975"50���~�![�>�}p������b�Y����;��Lq�S�~7���+�DH ���R������R��D��U)0���d��WfƟJ=�3���dU�;�PBeѲd�{7�]��Ĭ�S����o�\ַ����aLJw�b&WhȌ�7w��e�J��kS@%��ߥ�q�3յ���vy��U^�P5�t��}rj`��y0���f	�Zܥ[��i�ƈ~^��H�z�U��R�^_�P��ǹO ��y��~�>l--�������:���?,m����b ��hDh6(�s���ٚ(]�;�UV
Ī�T��X{#9Ck�1�)+嵰�!�(� ({�}{9��L�YV�0.��wI���	u�4�k����[1����aYЉ4k+�TCw�u���{nt8�r�^�Yg$!��GmѾ����^N8�Hy^y�4��Ѐ�U��/�s�`�(8_B�32�{]_�ʯf��\���*��������$��6�߿s�=�e�g�c3��u1o�ᤀ��qҊ�K)�r��D���7EfΙ�Б�؜)F���D��c���F�}��aՏ'��`l�h<���-�}h���K����>D�\��0gA�׷�cϚ7�*|�RkQ�{U���r�Ƅ]_]�QxFv�혆/ǆ��p�ǚfϑ>�r\T���i\teMX��u݈�Z��uS�m:��S}���r{q 8OmU���^&����4Zez�=�=IʻudU�Nצ`Fk��Myޢ]F��/#!�]yS���ywnМ�%�"�
R�L�t��NP�:��O����5�o{�Xޜb�"�He|JH=�u�d���\�ͺ�/=�m�>�Cw��MǙ��e��0�!u�T���?(�ͅB �b�eDT>_+\�+i��B��M31�g� ���8��	ӛ12��%m�.�o��W�N* �b�*�&|���K�}5�9J�mSQ�d���gj�/�*��&��B����/�KH�'�h�:M�b1�U,�X�R��Y'���،� �ۏ�33���-l�Z���;�p$A� ��ծ��,���L���(�%��t��Z�,뉚��h�3�۱�����<�b�ݕ׫D$j����iȗ"����yP�U�Ѕ�;^��^~�s�_ Yb� ������L��REBN�mQ�0��٤�z�4S�H_�P��t��bG�[<�{�)����u)6Pp�l,
RE�����IPI�s*�d��n�fP�\}�}�C N���*�r� W�PӮ8C��������K��?$��u(���J϶�)�>OD^6��3�����z4Y�(�dQ���^��V���]x�O�vN��55w�|$��ﶞZ� ��O���ߛ�.�op�$�*4f�f6z�&
sH�j[U<|��������.PL�6����L�5�=�v'n��Зڥ<�X����2!�m|"I$�դ� ���ľ��͟��U
��!�Hiȹ�&�^�`�q���t��;_L�忴e}�Q)��w�,���V��؅�זD�����F˚����H񿳮D�<�$��>�ڞ�ٸ��Ŷ��f/��~V,A�.��VZ 	�@�u�������]�;��3ڪ�S�N��9?e���tt���c�nw7KFF;=�Q������)s.�I���L����qRpeH��� }��^�z��K�aȦU���E�����&)zO=���j�$��uA5��j^��v3���^�hw�Z��]<�?�Άp�&�r
�$�É8�̐�v:1�fh�l)	F4����j��UW����v~��{8u�<�T!�6�5�:�a�hČ�&�;�z��/�f�f���'{g�s�-bY�P��e��.����P�d?��9�+�؂v�or�g�o�,e�ff�&mǝ��W�߸~�"�i�ح����Է8ƹ$�/P��> ���w���66��fmi�p��[�@��Ȉ�љ�l����p��'Up�}vWB�YWs[s�B�3��a�3Q#�ｓ�w5',�����`���_���[w8��	T������l��@��s���v*��Ҿʕ�ˊ�2�}�>���s���=��+�aOP�)�&�553s�{��s ��z���
�%�ȸ��T&��/Я;'�O�,(�]p�ͨMe�:�.��lM閳���KD�6��]w���Y^�F�^˰�dh�m����������v���MyCÚ��ٴ _o;�����r��=�@^{}Z��`dz���&��}9�r�L�;#�I��6�վ\}8N���rN"�*���U~߀户({`����M�\߰!ZB��mm���P���z�f���#Ya��)�oN�f..���h��Q��F�0X�>��(�䤔�RZ!YѫUDA�Q�W�{v�l|�QmU��0�h/����r�50�1�B�Yd*�  [I�և���v���ߌ��|`�<r�bF����K���)VY�Zs���L�z��Ϋ��\�@В����v��^g\d"z4���47]�vo9@՗�x�O;��he��y2P��h���+�א�s�c���lg�?���]k���dXۣ$82ބ��l��?2}@ϨM��%lzhP|FJ��3J,r1]c���}��M.�=�}�,D�K �Z��2���?B2_:KY�Z�����F%V)���Ӓ�1z'+	��r��Z�<�vf{!��.B��}��kf_�i3���wZ:I!�$o׏~m�k�{[������L�n5i:�r~�/V��Ydt����F@�ښ,�|�罔t�3D��Θ���Y%ыp� [�=aK���
U�/��h�w+ը\@��y4�˕��-\���v�F��R��<�g)unGv\�A�s:/�Y�0��52��fnmL�OӾΡ'ﾁ{��s�����D��"�&}+��8Sԭ$�M����D���Dl�e��	YX�H���]]ѣ������	�qd�y��t�o�{�Y�~�A+eӈY>�`���r���}�Gw	����[�-�>#�w���B��b�V��W�r0^o�[< G���%�zen]N��_A��-8�&�c}?U>P��Z��'�7H"a�H󮰜�ժ�=�����w�8k�W���s9q�i���*ەĘ�U8��]R�WN�����fB���s�Z���s�yLyq]���}v�z	��ew(yf�n�o�O"F�B�W� @��:�������u��T���yqi|��ɔ�Rzܺ׸��*(���NLѭ�M�Т�fL$����\Յ]4ĺNkÑ�����o���>j�\𳙯4S<c�l�B�~�B�R�	i��\#;��"2>IE�p�T%�@t��f��!��'ݖ���X�V�b��'J�����S����2���̟���W����@`�-_C���(�$2�դ:�ώ�<���fK/����繂tG^��9�g%�����F�p�<��p ��9�
�_|]���M����8�	���~�g�Ϸ�n^� [��~۟�fu��K�~�x��R��^�V�sW���s��=�'�A�X�s��(�/r��`��;��
�d�E��ļ7�N[ T\;�ted�g���:�/"������3���ᛝ��i��S�Y�S�����r�څ�%���C��Te)-�
a&�y1cF��>b�f{5��ή|#v��x�4 �)�����Ģp��+�O�^2<x[���G���T�-�
�ԴmX��h�5��ҹ�b���ʮ6����T��ʦ�a���#	)e��%]N�}vkC�I�s��d.X㏲����7��	�Ɓ��X(������t�朽Iq��s.Ef��bB�Mg5���r���;W�C�`�T�,�DGz�!*�:��|v�d�C�\��S���{o�%Z�WA�y�/J)Ad ����݅��QI%W�߲h�$`��K��d�y���U���;�̮��@�LL�B=������g�m�8�9����)��8Ͼ]�N�\����1�f���J�$7p�(�$�Pi5�c��u�.�IG6��i7ul]8����ܒ�f..B=W������"�h��v���q��mk�s �{���m��3T��]?G�_s%���0x�)����:��)`��?"j�$:tݯ��>�R7��pA,���Vr����m5)m�����K;�H9PW�]��ꇮ�<��c_��՘�,��c�:6����)�Y�wY�Ȩ4��zI��0�>�&n�AS����*q�����C�U{�pأ[���L��7^�^������/��mTgd��)�L�&��Wnf���������=���L:]���T͜a�7Fo.wR�
�]J>7��QYA~yk�B��>F`Y���ޓ��h�m����h����2�W\�����,�!�	��ֱ꾽�����b9���o7���堔��w�`<_L�7��u��םϛ�ߋ�����ve�I8��v��9��V�|m(�
�ѭ�<��Ż��8vf{��5�B�V�H�X�=��ao���k~N�����^X�����eۭg������}w�������5T{�ǽ?[�T.kp�<�y����*[�C=[b����D�$�fY7��[便��R���IYSE�0'�y����~^�W�r��EV���,8k޹�kf/|�]���{��{% ����FȪ{'Y~����t.���>����_^`�s�mS@��U`�[9瞱gܦW�`�>�"=3ե]��(1�B> }�Tj2�x�jU���~�C�0�lX`!s��.�pGE$��~O�j�os��}�w��6W��'�� 
�髼`��Y��}y��ǜ�#�sSd�iWO�b��umVK�z��-���3�W�W������9u�y~�Q3N��){�1��ya�?,�)�7������D"�,��5�1�GIL��N�ֹ�0����l͉�����\ ~���y$$��ޭ���?t�~�����.���3�����;5��f��%������9�+ѷ�w�����.�w���9�-�~��>��L{���]�����?}Y1o	�5
����3�H�^t���2{%5�u�nQ��%��J�G���6���{Ni����s�{���%OM����	��ޕxy^7��Q( �WBΫ��0#!�j��3�w�_�3�:�U��=k@�����u��m��Suk {t�v�a*���dUU�E1�5���h"����y�j�����7t]Ob+��)H19�U�y�Z�}X�q�\�@�H��wٿ���~�~3S�~��
�q<R;�թ�ʁ��<l�+��L>;�wl��;��w	Z�Wj�"Z�^��ŵ��RE�1��m\�V��";+��!���rP �w2	��S���"�����JD��lS���)����=46����t�φщyވ1>\h��9����5��׃mw*�g~w�1�|������2X���.T<���5"�m���N<�~4�����V4O֍gl���ڔ�g�gT�O�)-��^��9r�u ��[<�I�YZ#h��A�����>���&P�^���(}q��0��3~��:}�[�%�%D18��!�Xצ-��}J���ҮI�2j&�:9s�3�+K����g��r��.�uW�;/> C�GT"{�m��=@�Nc�I��
o��Y*�Z��ߢ�s{������}%rР2!Z3��Ȧ@Ph�0]߷s�}���e��J����ǹ�=� e�ɯ5�m�Î���pXj<�{�0��tX}<�%m��+lg:p������A�Vnow\�C��Zwgs&�)ϥ���(ލ��r��MQ�A�	��1��#���d-�CŜ��廩������+n��N^^͗q.*w���_�Y�
0V("*��]s>�˳5��E�L�z�Rk���oNͪ^���Ur]�qt�ޥ?IЂH��)���=S	䋟�>����9�~���]-/.]�ԥ��=�y6��È�*qx��:\�t'�{##��1ǋ��7�wa�߉;��v�}tQ\�y��{}S���T�D���Z�y��7�eEșU�Of�ו�x����� dp����D_�OC�j��v�*�3�8'״�f�:�=W�����A{%���:���'�o�S��\8Etև_gV���+s�c���i���9�$	�zwW����l^����f}���}�u�����}>��tn�+�������i���^9\��Z�@��ϋ�[��7�>���=��Ƿ�۠\�9�Wd��Ҹ��=�I�@��z��[I�8��R��D̸��E���ޮ�쾹pOx��h\�������'���B�߄��K0/v���@���)���X�.}7��N�\3&O�Vpv*+�Gk0N1���V������³�uHZٍ��S�����Gi�%ѕwz[��8��ܾV/X��by����^^k3�ّ;�$sЏc��V�\�j�.�k\q��R�3���5A�R�mH�f�?��Q���׌w�}gr�yuiM�5	μ���S��.+G9M����S���L�HKW.��5�t�%Cb�ۧ���uwv��:jKܶ�}U�L#lt�.�����-_���_h�=� �v��j>��#���Y�����9����t�ǽ2˞�}:#�$���a���vs�2�-.&�A��M�鴶R�1()��Z{���X��#o����4�q��[W҄�s�lg�0�F�2L�b�f.cF��h���r��<�u�w�A���d��^z��o<vQVD�}mͳ�N":X�`�'i��o�@�(�h3fd��20�L@�4��훛P�6$B��;��"�6&��I\|�ʣ��v�x^\�M#K���1�z��ƳgQ㺥f^��KO&�Iu;r�L�]jqN�͚�����ՕF��%TO�ޢqp����n(&�<;f-��{�Q_n�7�u�w�S����:b��N�y���.�c�EI<���L5������lm�kJĳ
��7#��tX�avC{K�)��
���H�#m��*�-l��]7�ת�����e^V=���욡��'����y���/�	�mJ|�1 i���F�2Us����W��Y��q����s��䫜�$���߇���c�
U�\^�pI�*Ѕ�e�O��l�W��U�`��l��0]�g�Z۪C1��1T"�K.b�������m2�T��+X��5H�Y��/��2��`�յ��T��eٱ�e�G
����/1^��Fܝ���ym�6ԙ��zF��:w<��6f���#�̸V����;�X^��sb>�c)��#���י��4;�zU��۹+vJ�3\�XNr�/�b�i�����q�Vmg^~E%�OD�rxvЛ�U΢;-�Y���Ru��2m�޲|���`αYvJ�����X���Fn
�%$��m{G-=X�R�Y5�М�E����ԃqd�4�WH��`���sc�����Vx����J�Iqܢ��b]���-�Ń-���Ս!�����;O&�͕�{l;vy���c9b�Y:�[��f�d�ųT�4q��9�������%{�q�m���P�UIjދ<Ab�mBl陼�	�ַ�T]�'��ւ�����fv8i�K2��v2���:���B��ל��y��mi)E����tl��8��p�n�]�������|�ǽ�mդO>��X���Z����Q��p�N'�p��-eo* Z�$��<��������23�9AJU�Ш��ݪ���hM�aĳ��b����Ćy!V+WĒh,�������2v]�)�0���ü�M�T�٨=/��YݜuQsٕ��c�땝'��,s}��ti�d���p�f��<������u����k������.#戟Q~����-꾋�T�z��Ó)�[>��LWL�+$��c���+k VZ׮Q��f4;�-5�q���u��t���8	�� ���G��q����vq�0�֩*�OF'��3}����
\��kV�}D�9MDt�$�Q���T�u9T�SX�]�&f@�u�׈Ab�j��\(��E��U�+�q�xTB�>_?�a���q��eQ�){
(j)e����O�Qf��{��\��deH7�n�=���"C1��W�6�U��Z�6�c`ݾ�o�k�vf��}7x|���U���-��X��pl�1�E�P5�t����(��g���e���u�������[잔�|�wv�5�B<E���t0O�2����MQ��jg�}�� &�dWY��"%�O&�3�f&g.�;��2���s�Dh� �wi.L�y��y}y�H�w#����B�e1BB���nV�����fw	���[t�lt?m!y�pEf�^C����qR�R�7��e�X8TMarC��[s,Ŕlzz��E��l�o�F.�z\�\˵���I/��+�?9�7pvW)����������9}�ޠ��3x	�]�ɱ�=:+�o-]�G-�4��>����	��B}�3%�r��
w{�px��O���(F8��i�3�q�%�i��	��3&ƒ�d^��Qx���q	��(ҧnz!Rdث�62�̠��~�~w$ѭ􅔡m�\$Y��5�c��#���48���w��Υ�m��B.�\+p+@>�}����Q�l^��U28*��T�
��f�`ǿO��/*k������HG�c��.�}��O`�/����G�z����"VH������p�<�y]� Q�;nw���,�@���'5x2Xw '�S�x�B��q!Z[����bU^��b����Z�9tԉ�&�.S޻�)^��;zSo�Ͼ�����" L��]#�W�ћ���K�g���ȝ^������w�
�C<����P�%!��=��Tb�(��>h�S�IK�H?nm�F���!��EÈ���J��w1U�n��o��brvh~xj�_�"�i���$Sm�	e��-(UowK��M��V`�s��8{l�g�kbǝY�bvw3I��7]hހ^�n^q��
bKI�w��X�ۇ	��c��-:�'N�{2%��\{f��k��EVV��*��eMzb9jۻ�$:;#��>���I��MaQ\%LB�1C5q_�| �]����N
��V�t�*���?z�oŦ>�GxX���8��Ө���Y��Ԛ�EU+�o�R���h�uoހJ��� �LV��h�����+ ����u9q���s���-9=���uX3��50�R��p|O��[on����~������C�.�E8�*@�;]�A�Z�OЇ�M�|���U��e4��-�i�¼�9QB=�ԫt���c��.�n7@7s�"����8��>�z=x�e$��=�SY �&q�
���z��|�y�u�=��+��C�m�1ɹ��1Q���ml)�";bB��� �<�N���ם��҅W���V��Y꛺7=œ�6��H�CS'�L��=s(�6o[F�t��T ��'���3�]�8�Q�rn5�4�u/��ە��1�#�mVJhfJ��0ӆo焵y1>�ᒭ�'�)���+z0�v��+~���<��*Gw��Z ��������8���;����;����w����
E��SIq�kX�kNe�"1���{�sW:s���o���J*���.�L�k��̵�yą��];5nk�[]�b�t��x�s�ͽ%۶�ҧ�h�^�J�nB]v�۰��eq�����QG��r�}Y�=P��i�?�dp���a܈����L]e��V�;_3ݶ\ox)���K��4���D��ӳcX�͸e��^(�%���9����(.��{	����>� �]��;fz�]A��pl�tU��
7^�L��6����JT}�޹O\VZ���鞁�����7�j�%�ARY�=�}�P�E/��苩����������fʰ�A����C���}�y�n�E�:;����SO��T�lMcU>���}������}�Y������J�p"��k q0<�Dd��t  ���g���s���l{4:�;�wé��\�"YJ�2��
�._��v���\�*d���|���}y�>���C�-uT�{��Ϻc�Ɋyj)#.�Ϥ| ��r�4:��$����0^��T�WΚ�(�T�eͻ��0zc$)��֮�A���hU4�&�bY��g��_����Y���5��#f��H�ɡ��7d|N�c_F�~W�*���f��m�a���i���Uv|7�iά,<ǃ��u������[��ML�&�fJ�('9��'G��mfj�yŝ���9L��e�Q�XX�m)�]-V�$��Ѭ���S.�k�Ұ_p#n?�v���o	�42៧6F�ֵ���gW�%f��h+G�vi��X�v�Q�=���b�vM��c�c��*N��ë����� ���`�r56��T3*�md�t���vNh�*pUKVm����	���xz)���}��Q�c�%U���������6(�䂯��{�v���31 ���G�U�]����v���$>�HM���EOM�iC_��.8��'�M�Lt�Q
4'>��sT3��������=-
:�\X�����*o�|=�^�4ȳ�!`�!gl��D���ʞ�vʹ~�����szP�:]Ã�pM��,�a:uu�M2�%=��t���Aj�NI��/]]�T�׷��~�s@�~K�[{���Z&r�g^�𝮸P^�1�l��u��]`S/��v���$F�A�Dao޼%<���1k_�?�/'4i�=4O`=�	�5w����Իc,c��4W ��>������qYf�Zɪ��g%��7n�:TP�Fs�����$o�BB�'7�QT��X�3�Nf΄ʞ�O�}�˝� �O�F8�P.�]	�Y&g�_�r�<��k}Ϸ�.��KǮ8X
."��ER)XJ�c�sY�]{�c��ӓr���}�ec�f2U�J'mƚ ŝ�Ḫ�E�Xru[�܈g�T�ªMY���$�鷬7��=#%�u�#��!<_!zpfϭ�UN0�.�=H=5΄��N�q=�8ɱR!��CbG\���2����{_v�؋�򞨯dɐղC��W����#=8�o.3��~�A�V�����97ʻ=3Ӈm�Y��M���M�s��^%��d��+=N�t��[;��s���Z�΍��ڝ]1�+�u����&�
�{�o>����J}��%����3��{���YoL�^Afn�t�z�G�	3�'�6�Z<��v�ڒ��@��{0��������%��1�����z��� �v�M�_����
Օ�q�R�n��5$�%�5��v9<���l�m�� q����\M�����q�K�}�媮��Aig��
p��vX���V�4�����gu۳�q��c�U.���]�9��X��f|���O��өS������=֧��KW)�a�BD��y�	�U?��8��5�@����f�8�!o��%q��[J���ɔ�U^U�Q7NC�F�l����*���z:���è�����r�-����i'B�p>�AD�i��Y���c����.�;�2�F��
#V�	��p�b�q�l0������K��+%ݙ,���+�h�E��ˏ���������}���9��h��6=NK�����婱�4����l7=��c-����s2�A:���n�5Wb�^�ד��Q�"���ߴ��\�Y����Z�y]��oF#�C����	��}��U��vNoF�xE2J��p�G�DU8&���d��;m���Y=s�M�躧lި�W= WٲG���Ly�~r�t��|s�b��Z�/��,(r�=� d��5&2��bc@?���,n��q�ꉋJ?^��R��M����^��E,ص(;K�Ofؘ�"�I��b_eD���pzi�����r\�n��j�TJ�8�_�~�zH��G��nA�b�4�Jf�2�^�Xg*�I��J����=3�;7:�T���P�jlR�p2�_�܋؁��$�z�P�ԮOq�7���6����|~�}�Nճ�(��BT�k�$�>��|�[y���ʜ������TVP 3�T��Zs⊃>� o[�ɽJ�PYucI��B�d�bۍ���Ed!\\F��0|�h����l�7Y��l�d=���4-��r$j���q}��|kH��,nK�k�1���)pj�x6���n�vb��\ǂ)t&JR�ȟRt�
���y>��M��˵@����B���-���9��$g.�3���WV\���;����a$\�,��p'c0}논C��8�ȶA[ORS���οN�?^��4���W�N�^�0�C�ܫ�LIA�t�4�v+Z۵uO��D��[t>W�q���S�Tp��"|���|��'�̸.�G��H���� �I���BM��~�K����ǘ�C�C��b2E�!]�u�Q��/�ܥ}3q7^%����NLٻc�&e�]���!0�R����}��D��|U�����v6�f�1}G�o�!�z/x��fWg�G�����R�=����W1��	��oB���,���bK~������q;���JA���#��/���#^�%�(*=��(=�(����|;����-�/�{���5qT�}��и��n&qL�ê�,���*��D5�p����x�*Ǭcqç�5QX�Gd�����t���e��N�\�k�&�ݧ$��5y'=��N��<�>��K�4���Po.�	а���#�!�&b��~�+c��m�ِ4�0���sr�æ>ȈI|	��AO� >�>���[�NJbN_B�7Ϸ?)�3bԊk������בv,�B��+L_�.�}
	84����J��c
����hKE��*��":D�����Ht(��fH�W�j���%� &Mt�P�2��q�#)�1��������j��t��7�e��(v�/B�/T黋��'\�bLxN��|�;���7���xj�Y8~}3.]K�E>�AJ�p����D�^�c����Fs��H��9�s�{�L�krb����nWr�o=�>�W6�`��L�Q������\Q�o�O$�R���1��Ɛ}������39�y�l����5���u{���sj9T��8_5��}s_}ˬc�����z�+���	f0���F�{�D�����p�u�����Q���jԄ���b:N~�#�J��z.:5Q�ކhE���� ��3�޹M�W��15}�����=}��<����2kݏ��?�����`�6m}�!�eG���6�GzJ������ү�g�tX}y�r�M^S����'}VyZ�v86'�.�Χ7٬_���l���\F�Y.�B퓪��GG�>���F�7&e�irLBc�N�>�˱��ل�g���L\�I����
�ڜ�5�uf}�T�]�Q��fν٪:s����t+�(��E�u8��5`����P�̻�Xyqn=O�#͸�߳λ�훷�ئ�٤����@�c����4>��M��_�@�s"��kw�>���S׫<�^��jP�GzWR+�u{9�Â��&�VA���G�i�������7������4#��H]md{�
ھU�L�_^p���G�aJʝ*�/��c�(�� e{�У��u�_\��.����#���q����t�y��)��WL�ߑ<uQs�#"��]�P������)������@��U�N)����k��|�G\e�]�}c�=v���ne��q!�m�	0�C�J�v3ʝ?���}�xw�����6�;��6>lC��|""�IbA9u0���i~������R�����ק�əľr{������j��h���v/aT�Z�TO���5_D�+���� �=�(���h��Z9z�s\7ËSe���]:�N�^b��E����R��-��	b2�Wj�l+�)�e��M\��3�Ղ^իX��U�����H
ߐyZ���Zx���h0�-��u\�/�lS�ʶ��4r��nZU�����tRa�TK�h�k�U	7���ui�K�Dэ�/�#��,�`;|�=Αު]�2:fX9����]��.�A�B��ܐ���[T�ϩ����t	U�D�94��}���bU��r�)��:�"q��4E@I�m���(HG*�#&ڼ����Ak_kӆ�ݛ��Mh��v�+���(�� ���*b�,j�]D��Fa�X���^o8r���᧕��X0��T������s4ܸ�V�[-�����7j����	u,یX6�$�g5�X��D�9A��X���˫B�Z�&�M��"��Y��a���<������h�-�	%�6��~���p=���������_k�����8�r��v�������m���q�{��ݑ����
���-����7����;V�Tx��45�̣U���O��ok-�S D�%�pr�v�ۚ����ٜ�k֯/u�W�q;���n"��z���O�Z;����r�nu�8{�]��e�*�au�NwM����2I;A4�i$�w[�W�Q�����i�ۦ�X�%6_U�{�EӤ��o�}���R̧;;N��8�!wӂ�g�`F���[��,���	�_ˠ	8�s=G���ޒ��%��`~�fU��
2X��ܾ͈��j��fV�ʭK�1v��.'�5X�GF����б��A�$ef��v��s�f����%��u�K���;ەkCj���Wlz������m��M���MS�33X����nDjZ�)��r-�d<��c��RJ�l��Uh����0��q��;I�;�X�e��fY���N�ڷ�.d8�wW.,�Yo;i_E*��]9@K ���N��v�ΓufM�fK��5�"���<݋j.z[�G�Q���;6��� Gb�#�V�,�iS��ggC�v�$��"�UveH�w`+��tN�O��L �+5�l��Ҝ�Sga�������X�x't΃�����8SM�c�#��J�d���w{���J��2���o4�-g�xD��F�Q4�۶(��ͨQ��q�� �m]���8�7�g#O�F�`b�s���;�I�-<��0�����N_˞�o�5����(�M��'��7+�|w	����1��D3i9�@|H��x�t��
]B������P�[��)c�d���!^ZuM����!a;�\�Xc�N7�o�'��v͚���@q|���%�e7)�K
_Gj��@�C7s�����3��WŊ���E������<���Ok��<.�תl�u��W�3|�r	�wU;��vs��)�_{*q�~��"�nئ�v7y���5��1�k����3wL����;�F��8�`���y2��*�<�p]s��0+Z�ci��s�TjLE�O���3\���sY:#��3�e���݆��J��fyJ���57�"�����k�7�]��ȏS�Cf>�v��xU#ә��E}�@ }o�\僛�u�Y�]D�d{�k4uMy*�jD�=fn|INo����\l�4�?V������]�Rz�}�����5�W,���de@���H��Ⲿ��o�ԥ��Ԝ��ȇ%=U!�w��{�dR9�w������g�6'�6�E���v"8r}�}Qb��`��#��Q��{]���ǌ��zo�-l�e2Ex��8���͹:�Ǝ*�(���#v�oӜ��>��"ť�3����u�������c�to^j�ߖ�pш�{�P(���O��s��G���&��ڹ�v�â�7l�R�#�f��z�����3;���4'��:��h/g$􈩓Nu�+�/`훩��έk*�)çt�}ܔ����m.�3�b��`=��9.�:aas��w��/gp�z����ṣ)�a ��m��� {��vv��q;B����Zـ}�[KO��k���h����'�'��ns)�\*��X�zt��o�fytv�kN#�+4�8�͓r�~���>�7}1e�<꓄�<멉��@mP� J�-�b˨ܹXH�r�8{����o�lק��|���� ;��|:���_u�.�-3�G9�ɼϲ�=�2���1�1�uOE���C��`,|���:�J�{��>+ٕX���c��qϾ��kNˁd�x;�>hf�I{�Ly��}�~�hg��ގ��p���Ƚ��v#P��������+ G����o���s�)��u���I��ݔOʥ�!�J��8n���UOO��o���)�����W����_�k= _����Q��|
�c�0<W]�����F@�C�1�����Z%*������F ��P�-{��2�
I�����۷�Z����i�ں:1uWHJ\��L��m��t�Y⣖�t�}ݔ1.��ã�w.��2�E�̄�+�Ը�̀vG�(�oWv�w3�����8s��Q5o�C�y�e�uC~�U�c]��;�ށ���|b����`5��YmJ�KF$��7��X�B�\:���,]:����!����O[><:�WS�y�"���a�$8��w�Tߣ%��H7��*�O���͘~�]Ol+�*B���5��o,��U�aZUw��\�*1i�/��X���C4�U���m����~�><'��Ɋ;�C>��8�"��Z��q@&�,!u߄?{��e��7�D���/	�l��q�z�jW\3v8j�0b�|#���֧��R;{
& �v3�{����݀V�K���x1���ГLU��5�c8qҕ�*���o��	p�{��A����z;���/���C���;q�ڶb�3cca�ϯ��^����U�(V�U�5�����c��o�Q�Jް܊��⼣i
��s��ji������X��Um�e�n��c�*�����;��/{���Μ蜮��Jy�� PKruq���9����涠�;ݙ��\D�]�ks�jc��-#vѼ{��ɔ���
��'�v"�����B��֓t��[q{�����$BY�a�=��
N��h������w`��߀�Yp�gu�!U�:3�����I߯�G|�Wy	�^��ވ�r
z� ��0�z7<���x���󵚶��ro�򁜎u���w�����,�9k�/m��3q2���xa���h��*�p
� _J�;���@־�=��W
u�]���[���ug�`�}����w��xz{>�)~*ac=���o�Oy���U�s����>�7X������W�V��o^������.�W�n]x,x��=��V5:�6o~^�PtA�	�׷��S�=���Ƨ4I���S�ޚ��sJM�8��z1Ab�������w����U~#�>����m\��*���]+�w2?NĔ��y�U�(^��S�=��c��w�g^57���>��	zR̙��s\(�����L�w���K*Odҙ�Zf.���J��{���_��{w�fk�h��7�Oks����z]-X"��3N#��d�z�1X��G��G,rs����mp���D���ei��XE)�^;%��l�C�tj��\po���؀>��N@����7�;:&ż�U#��SN��b�QZ�>�[g�ү��>yýϩ��+�J�^��EV�S�qk����R_�;�d��^�=ᙵ~������n�ɯ��j�*�;�}K��ǖLP��^���E)�O�!o�w�3G܌��{�����3Y���	�η.Y7f�;�#Bȶ��Ҕ>�Lx+A,ף�n�:���aK�!Y~W��V�M��ƿa~��44��6坴%���`=w;B	���J�ܷ,���y֞b���&� ����)lm�
/���^� D
�e�o`i����3�yT;�p�(Rb�'�t>8g��T3uK�E����f�u���k��A������OJ�pv�U]<jϣ������~��eE>y
h`�Ӿz�:�����:�{ٝ�ۃk�=��q��iDuO����'���}�#�Z{q9�����x�P�+M�⊬�z��4�Cӫ�F:kC���tU��N������s��F��I[��ݣq�)�RM˸f�::�r^��k4׆r���4m1F��,K�79���*��U�n����kk�z�ѿG��z��^V�PY���4�q�����'�E=1���q�t�d�j����oh__U�����]�gsڽ��Lz�w'Ɣ;#��儛ݖ�^˖xw)�F�V��HqV�D>䏸Hɍ�J;ِG�X�Y���X�s'*b�b��O�*�?@��ܮ1���z�h��Өflg���o]�<�8|�����C�@Y���
/�)}wSꃆ�@7{3uԅe���G��0�Md�;�R\�f�g_A��I����1�����]u��)��̹�
�h�S��>í� =�˚4ཾ��"b�el>����y����hoR�ըtUR��
jrZKz�L̻\2&�x"���Y��{
�w���~�x𛎎Hz�f�٭8�zR�%n4zU�ñz���"���]��^��l�^oC�S���my��ޭ\5c��H�=n���R�|�&�i|�VX�A.�-�c���)�;��J6Թ�Bx�^�HD⌿�ӽ���E���}3�֧�d��(�^�����R�_�sd��됨���$��e�L�?�!.��s��v#��>���}���"��8�N���c�l�`=]�1�9�%��]���'~�7�#����ɖ��5�da����K�u��}`H���̻=����y���8[[�o0�nV,�C���i�d��ѡ�v�5{+�vJ���Ňu�i�~�נ�u����|��J}:=񡶍�F��N�&j���9�[+�f-~���hN[ s�����s��x���!���� �ݕ�n���8�8����z�ʎ�c�ĆS���$�媞g���>�Y�6�D�͛���>����Hoގ�#�ƄA��)��~��7�kW�����shD��Juޱ�DN�2�9B�oش>"Yzx�o.ǃc�?u-V��Cm�ng5%w�]l��kl��C1�(Zb�t{zW�4Ǆr��j��`=P��u4�:Uf ���ze�廬�`=��N!=3���!vMh&���yO����=]�Y�X�����}ӓ0�.[����ݡS{:�o�+��#�6�s�&8}�|V�{I2�fz^�=1��9��J�B�}a�ټ&���X�b��$zι?�m���~�2�ͼպ,����J*��ȋcx؊Q�`�(t��-{�XS����]�:fEح��* ���N2_Ǎ���1�&�U�5�b�a�]�3~�Z��dns(��>1�緞e	�xiU2z{w���j�w���錏��*Ar����ظ�z�`Y�j������t�~����@G�fK�ʼ�t��	YiGO���	r�����^���[�3B�_3S������#���Y5�մ���G�x�y��i@1C��O.Ȉ(��,虌�^���8%��ʽ��O�}�1�;UÑ��P�4���y�xQ��Υ�50a���^�b����$s��ԗ�����"�W�r�v�q��gxWwa��ޓ�[�
����>�� ��`�bDT`�A#�l73�� !�.�'YW�\�N��K{*L`kJ���A�mAAK�F�(�o9��]q��^��ܱ9F�������Ee����t�&:��G��i��1s�{�]����#]����g� =�ڽ�ѥ[>����pY�`�ڲ2����+�TUV/\]1�q��������Sh��G�r��w�YI��|%[�a
G�r��zݫ�T��\�27��ݯY�o�5Q��0>��+8���|�tj��=����@�X�1�O�3[1���8�E2Ǉp#,����4)mʻӘQ�Bz}cN!�W�6;��iI�H}���������j(��*%��z2b�ko��B7V�B��v�wA�˱�ᢼǍz'��TOu8�����
����ifu9�SU�tKھ�������䫕���ܻ�k-����4=��P�n�ƶ���D�\�ן^����}1��Y�U�U�j)}�]/�������<WC���<���~���q�P�#Sq��׹��6s�����l����a���2< �!2SY
j�`�!�qu4���y��3�a�B@8�E@ B&� tug��
R�����GUҬ������&��N(/��#OP�j�l�mK �� ��im����u�/'<�X��ykA��*qH��;�)ν����#�.��5U(=�A�4f� ^n
i��P�G5|���e�C�l�1=/sRȚմލ_p�h���E��v�LD�c�?��p������T��1Us�x`�����}WNi1ʲ�t#���:���_�������}P������ڼgz.�5�xr~i�q��1��k��S�<)��iE��͍������:�>�a�۞S�ǃ���3j/ow��@-:��<v=�RA��u�v_��d-�";~.�b��ŉ)|Jԣ�������>�9���6��S�_}�v*�G�&�~T�d7A����]������K�%X�d�'[Jq^��@�OxM��R�#tc�S�QLi�uF�yN��-�mU��G0�i���೙p��f������2WL�����߹�k_��� �l|}�;�t A7b��oV{|���u=��{0l�t���Zz�W4�wtj����*��.�"pyK��Ò�Ҏ �d����}4*�.�o�#P��^v�Щ\���7�>��A���mp�B�s�� f��Z��7y
Gl�\��6龪u�x�,�n���5�m{�����{�_�x�kz��2y	�����v�~���r��e�˺eʹvF X�ve�n�%ev2��-�r@>�h�ʙK�B0�.��}��o$�j�v�G������xV�o�7g$�;�߽N�q�\�_ft!�_d� ���/va�n�I�|�4hî�Lo�㽲��4��$4�0;�a�@�� J�s﹛�M�q��Ϲ߼�g!��+�����]hgw�2!>��sg���'7m�/
"+1���I��2	E�A�T�d�\r�'P�q4C�D��V;�����Nf��1���Ȳ�镛\�{�af�6���L=���yAϹmH?�h=Ѭ�B�`�x�q�ȫ��[�lf�5�ʾ�=}��9"jsy��S`,�2�-2�H��>w�S]y0b�h�B��n8�Fk5��*����j���,�	�Yt��SX,���F�ޥgq��ϖ�7h~"�>(/�b����p�&�{�3no�s�q��pd�̒@�(�j�{��&�7R�:I]�X��x�	�d��#��VA�%� �� �=���6�; �����|[sE��aT��x��f
����G�
�=�h6geT�J�t���+�!�%�{d+�s��h�ךqv�)���
;nγ��ݱr{z)�\�ed����F�P�ļ�i��L(��T|w��r�W;ܿ�AX�rIo�}#��W�,Nmn��LGW	�[��-]I!j�����֋�����{�r�Yw=�I��atL� t�2é=��z�ܽ4F��3�(2b(�����q�z�IS�,��~a��������/MvM�\n������B�s��[�n�c-I�ٰef\�\���NA�/@xE�&���?q�  �|�\�<�j���Z8a��睵�p�1��������� ������dt��"�����4���2rc2wfe[��Н�Zg�9Z���{K��>8�F6j�>.��7ur���w-���L�L�wۘ�R���.�-r2��4w�9��g+BI;�������GO]�-�ϳ/{ ���G�r�L���]�ت�S{��v�g9�T+���]��>ʗM�Գt�Q1�TG(u�~�wx2
�U��4�)t/w�����%�k�_;� �y�_A��n�>�`��"�9�K+O�:&��rK�NV���EH�Y�T�[���7sv`�%*��w�}(�VL���z��rL��J��m��1�X��z��ے&�U��ET+J4_ ��[����J��3��n�3J�|�5pP���<'�����S�6��Ѕ�2�hP݌�p�+��ZT�n��H"p��w�z��b��H:]�n��I� �w/V��.&�=�-�<��$���&�~���w�,����k<I�3�<d�n��W_.٭��1x�O��}+Wr��i��+ã�\u�s.�vdb����r��v-=�Xq�*�%v�m�C��%��*shu�����[�^�TY��ƤA���fP��:Y����l��a�*צ��\�;g�=ҽ��/��M����t����~��0�须��dU�o܂�N.�4��S��߾�����[�^�#�M�
�^G|��f��V��U�/�q�p>�ʿcI\�N	�{�%�}�;�*�pӊOsz{l{U�	����'rE��k�o�{��=�X��w:��N,�T�n�d͝]������ �nG�g��V�p�ɕ}����Π��z��0�&�̽n�L�A�4�Ǣ��b)v�:����y� �����阻�����IvAu���w|�~��d���0�F����6�snŬθ�O�ģ�Wd�ǷVf���%Z���q����=��u���^W��L�f�|� }������bo6���5�v��r�."x�^hi&���kU����*��j2�[��<�����Kg,\y���|,����ykeu�kou�͈iE:[���Qu,=i�#4h��S�c/�S�]�G;�Z%mX�r�.(o�Z�y�����<��6>7�����l͇��ӝ��S���/#��q��]�3m�V�:4�o7���~�!�o��7���ٚ��)����}��z�y7^���3P;�rkwV��@V]Q��R���d1����F�ً��"�G�I�"��f��&�:1P������F�-Xu�f�x�x4���t����Z�ܿ߫���NԲ�[܋���>�:}&���"�onw�u�W=���{2���qt�WD��A�hK_��ה.V�!VyVZϫ�o�����5�4���B/�9d��p�h4�� �!>��j;��X����b��U�մ�p���S}:j��
�ok�w.V�n,���=��z�����]{��n���}�{��%�]���l�ؗ�$����R�za��S���G����e�)���+��kz�Y��ݘ.U���A&�D�ɗd"��5wq��=�{义�j��/�*��6�EQc"n�\�*�K�[�_ml��J79G��V�����È꡹q�e�Bw���gd4�iQ�oI�r���Lbcb��&�w�WO}Tu�����g�d���nW�.�Еk\D��}��c�>��Az���*^9��s��7�G�Vp�����{9ov����{�㓎>�F�N���'=��k�3�o���(mߺ�Z�y��s?�����5<dz�:�dz���N���>�e�ٽ5�5zo+s�7�M�(���=��1����[^��7hw�ts�i��gkn��Դ�A���f5\�fq�d=_D}�=��"e���;.�B��3�Y�Ԟz��&(pR����l���9��Q��Љ�p�&_��@��]D��=͟qC�>S@b�a�ԝ��3DvLeUn��C}�@���骜���w����zOK�杭�՜1#���a��9[PI�4BF+���}�U�}�O���I���`��<�(��}����Yga����V����+��f?;b"~f fP�K���W)�Vc(0o��ww��W�v�/���7q�9i�}�����\�#1�Y4_YS{��n7��.�� ŇK�Uׄ��N<�<��17��O���wj���� ���u��y}G��{��(�O{u������	��*���Y���1ð���e�~uC��o'�gĕ�.y7�uĹ�vH�٣~�5��eG	�>y&ϛX>������h��}�>��K(�w�J[N���ñ�.D�\�wG-����}�|�rĺ�����yTZ������p�Y�۰����� w�s\ӗXO�bqmx|`Y��5���7W��<4��!��cf���V?u�;�P�C�}ݒ?-���JkѶmm���=ojg/��`��2ҡ��w��ڨJ˾wjo%�K'U��Tf�|�ٹ۔���h��#���㨮������݃s�M���D?�*�'���tuے�+~-=�M!NJ�_h��YQ��l��zM���Q���Q>����o71\���L�8\�W�d���O�Z�1N�ԹC�X��3Ծ2���2�
���,����ط��Z�����+�3}ˬ�ݾ��d��1���Ǝ뼛V�����1+=��8xG�.���eu�Tݺ7�������`��^�Ņ�c���ۛ�g��&`��v]�"߿�R��ݿ��"��@�k{�т�S��i�뗺<���|=�f[���6�mburW%�l[D��mb��]�Y������U��M�يQ+�w\��̽�)�s��]c�6G_<Mt��;�,b���G�V��`["n��JX߹ꫳ_�����ou�g�V�߆G��;E@ u�;�i=���u�Z��C��g菣BN��C� �-��i�1{{2{r�R��.�(H����eVpjE�i���=tm����ʈ�}����+26��>`eĪ�r ��O����!�#�*{~���lN=o+���^��jq͜s����A�lKgcg"�����-���je���������J�j�;��zm�R�Ȏ��$��k(���M:������iۣN�ꭙ
_ �hEl:<�!X���@��79������5����.��{��m�q�����`��b1�J�C|e�g:&�ce�L5,�pf�X��Qn\�d���Q�����Zz76Q��$Fek�,|G�����?�E��}N�TDJɎu|�{7�3-Y�g^�K���9pڤ2�֪�S�Պ#�lY�?U('*���bFW�����N~;�^�V�-��C��⯗9�a6�r60�&��]�.�}�t\#�Z�N����~� �g&�����C�#���,͉��W�^�����x�Vr|ϗ��uw�W��/��
؃��j5��Tt;���'�C�:u��i���k���W�S{ć�۔:���x���A��?��5�A�FEn͎��Ps�E,��<��_�u���G��N�X�W�~l�^|>�競s..����:�Ц���n�R�H���m+.༁��݌�b���T�6iu�=�B5XVt_1s����M�����bwQ�9ȼ�7������r�ך�E�Q�%+�.��7��?��1��Y2*$Y��t\S#V*��0r�"\]n�/���[X?Z��u�v3r��_،d����V�.��%{�Q}LOײqY�Ʊ��Bm�j"��^�ז���5v�2��Α�9�4���\�K$/Q�@H�@��N���nܩ>N,L�Y�ӧD�>���;[5�^F��UN]>d9�ַ;��1��{Ut91�`n��jm+u|�O�	���Bk������f��w�&f���L�C�.���]���!��c��M�n]|>��lW�{7��Fp�c�^�)��[�i��>/;�V��@�k�W�]z��>��)�iDF���������k7�s����{�E��wo�4�w�]�۵�QLWE-~���������z�]L�|#1g��%��]Y����U�;�ߡ-�}��'�Ze�v�1�B7���=��Ն�E��_�n�}go��.�WU�~�n���8���� /��G�P;������aP�" G4�s[�I������5��T�~�g��i�r�����8,�f�����U���uW��b�.��V��E��)Y�=��L��N}ǧ��;.
8&!�R��Da}�g�9������������ێ&-U�=񫥝x�70��nq�RK����_��Q����2S�R�lJ�ٓ�̐CpP�X�o�1��Y���u�+2�����/b La"m-T�w5�o,^�{C�}��Q����U���_�}a��:���U'U������ M�}���Sμ�r��w�+�^]8SG:/�׶#)ڰ�=��;^j�(��^�6�]�m5�<<��^���=�gi<���?wu��><w
*�w*��X~=/��}q9�����I=�UI�z>�@I� �͖��D��k�Ç�w����� �M�h�ެz�M�I=x#Ѿ���S�@0	���^٪���R�q~�_{��� �e( wU�}j&f!na��f*�G2>��0*����Y�v�.�mþ;����f��n����p�}"6�އ��vEWS�/XSy�)<b�:��D�oê�{�Å����ܱ�5'��w�������_J�S�ճ�уr��F9��S���k�q0��Ha�kM�.�.J���1�w[�y��s����90�v�9�U�*��VT.���Y\��I�	��:�DT�)��,I��k%�;i>y���eg1%�Sa��/:mt����/&�9��vf��-�Z�Yo��<�+��c���ʏ�=u��ܗ���> k g�V{�; 5Mb�S�ѱ'��E��x���7�H~�<�"p,��wB[�:V�^۽��h"�b�05�Ø�{��>�*z��/���|K������k{�O_��:]�d��^���R�%���[I���ꪣ�љ����� ���7�y�7����5�i��^�m��7~��Х��V)�x���|I܋Y�K��Zo�Z�aU�r��p+�#כ�.�y|���#y��xC[ou�b���>���ή�C#'��m{��I��I�EF+�}1� �=&�o��B�}��X҆��ۓ�߫����6V_����ҡ%c+}�}�za�R�e�^�鱕��z�3/m��ˡ}}��]��Mě������y���-ev�@�p3.�/z���r�^��˵�Ѧe��t:�ov�Y#73��/�$&���]gm�"����X��dgQ\��[8]K��%��l�:�F�v�OE��N�G`<V<9�.�c]]P��%��y�W�𻺺㫬��ht���Nɽ�aUs'a7��jG����%��pe�[6�t �Ǎ��E�r����'Ve��/J�we8������n���8G�g73� �B�U�yR'�+�N��gus�OeCM���	Y�G��__oE:�o�Y'n���_�g�'�����>�۝����0p�^t:A�K���\�y�Ҭ�V��[q�=$�ʦ�^������R��&�\�}�f?w�߷��/�v�&iVMvx�4nkn��&����C��,��힎����y�B����O�<b�W��7C�1E�}��R��D2�r C�9y��^�Ī��L�?z�a����+�ϛqFK��ݙ�8s�tcr�>������B�>,{Xi�J�{��1i�P��{c�>}�p\��^^RP�]���Y�iy��3�Q�gNɟS�/�t�5���Ԭ�JD�~�wQ��K7i���2L��N���wy{��-s��ɹ81"�"��}-�bs�"��.Y/��F�y�����^�-�zm�{�Q�G(�u7م�}H�|s���5^��2���1l{ �Y,;CK�ז�����	�-�Z�X������>��UP��^l"�,�o�xl�z
�P��Q�[��|�ث������ӄ��i�v��6孬Y9,�ԫ�F��=��u��Y�q�Y@{ǘH|�J�1�}��:}�ߍ�{�}�l�˷��'�����ݖڕ"�
>�fӾi6�� �H� �AM�@�
j�8��ݜ�r�٦����E>��iy�!�l�o��:��0����&6��'��Օy4^��y�	�ޜ��/6�'h����*��SwN��l]�9���7��[z��B�C��u0�
ϤHt����!N�f��.^�yo뛛{�u��4kY�Y��s��K��!�ef�U�HQZ��Ѯ�fS���`��!����B�!6�@/"6�(C��m K(a\�P�`̥��f3�0|�u��xJ#%_r��z�W����@�H!8w�43�������cH$}^_��
;�%�b��}�$E���
��R&�Y�����J�F�c�K�ښ3�[��["ė:��v�a�H6v$Ma��ee�J��$_-?Lp��:�z�ep�6��K�rˬ�!\��	{��u�Ң���<��b��#4,��.s�F+.b�(� �_1�f�����ǈ�s��N�F��o%�U;f=�kh��qoCq�1}�I�3���2��Hr'�J�{qr�G���c�Zq}]*�	^����z���7�r,xq9�&9���C�B�h`T�	�-��S��wU��Te`hj'{n�Wma
�ԬN�<+*D�<�]��q�9D��[���׽�q��޲M�,�+b.�!�4M�ND'B�����ډ���U��b$o9���A�G5-����L��.����1��5o����FU7���<�:���>͜���)�ӗ��j�]V���E��K����b�xZ2ޡKZ�^�\��R�Gtdѹ��q8��@�9}�f��Vt�Y9}CPp]��x�̀�(O�f<�[��U)`F(��w5W��͌�/�����~GC��Ұߜ�W�:T��	\��>I�-�r��#��2q��v����ăӈ�̷�S��#�q[���)W8i�.�G�mZ�Nì��3	ޔ�ҏ��=�ޢ��V鞍�ݠ�68>���/^Q�P5#�ΘN�qT�f�;�Je0L{�c�k�����'7lQ8�v��q����Kճe�z@F�|L��%e�y�iy�:0��*�����Va���d8e�lM�٢���������Iۏ-����Ѩ�DU�f�3n\�@���e��4RZk1k� ��û��tME�R�=�Y�s�v%���@�P����Q�s�Υ�����`��T���t?=���5�J|�mJ��Ÿ�Ie�2�d��;P�5�W������;��E's};����0>�|���5����|��Yߪ����'�q��<3{�Y"ҷ�/tIՔoCs}Ss'|�j�ܮ�Wn[��͠�0v�d����@�;n��R=M�����SycrwT�@,�w��Z���	���Ѷ�X�z���k������������u��@d��6�9�}�D�v�^v����"�o��������>�����/���*�97��%���x�U���,��/.��7�Y�~Y�nt}�>���:�u��S���#E�UƵ�>�����@���ר����<��>�1��-"R�S�<��ۋwz�Ly��o\b������U���m�̫ߏP3�߱)����i��~Q�f�KT���ٮ�~���}�,��W�{N�f�so��։���_<���A�|�ֽኟ��\W�fK�o]v�4�TCb��1��xJk���K%��$p71��1���/-eY��׫��7���g�G.��%�ç.J$�-=}ڵr�\76�S�̧�vt����F��)t���3���5�u�'�Z�)�s'�ls=y~��C��}�<9����[ZC���Y;tbkݫǍܪ@��']��c�1����A��vUK���D�r�ռ� }�����蟵!�0}w.3Y��1���rP��&*#���Z�8y���A�����?\ѭ��9���cit�I��vt������"��3~���*�eRM�������<�{X$
��EGE]g�9�qG��ף�
��elʜ�\6�>8w'����ޘ�U�?t�<�]���O�����9�1��\�O�r�PRr�X<m^�1�ETfΞu�4��.<���~9g����ʺ	�1V���x������'vOF���<�Ë�R�f#@y�cט��',��og-|���
��\z�	�̀��Ƙ���|\���9��������m�N^�va2���&K��x�}��|{���%e������QdA�}�v��f	����D;q�ۚ�m��ɬ^��7Y��d�
J�f�;�mbD^�9q�V5�$״���Pv�h�:ӻ�F�8p�7p�r��.v��˱�F����}\�����NY^/켣 u-���ǥvb߯7�ܠ���t�:���W߮�G� {����x7��1M�d}���f�Dڝ3�ܻZ����:��x�;��T�?]�,hAw����Џ��{�pS�-�#��J�\הR��)�}�ڐ��䩠*nr19��� ����z�=/���/(8�������e9k* �^TbJ�3���W!Y3�}B��f�WmUB��D��?}�.�U�8��nU���U���Q�>8+�8�'>�y�#�E���1 D^v־�N�p�*�Xc�|=!ۛ"'�ЛXQ�%���Q}-�}��x���te_1��eg�T!&�}Y��\��X�z@
l}]�o�f�uLӨ>�mO���"���Yp�S�T��΃Z^��[	�q��<ݟbk��5���K���]�Hi�M� ��+�W@/  ���5�������r��p>}���E�E�v�3vbߴX��5�S�܃&�zCMS�Uy$p{Dh�)���7�tW�[ڬ9k�Tو1x��8`��v��h���Ul� Z�+/�FC�'��m0�w���}��S/5����u��[�����s��Țu�ҿw��u
��V�	���o�m��M�h��&}��w`s�v�^�����������}���Ψ��On��%��8���:�D�G;޹歉u'+��| @ �x�86>�hl��۲H���]_.G��k�w����gXȤ"�9U��p;����l��M�GB��߹�,h_�߇3�J���{��C��hV�{�h^�eԢK���=��=���#g-����޸������*�Cp��:6!ᎈ��Ջ3�,�����<p�݋��^���{"Pr�园�/��9
L��0�]��,�=��Vs���].�ӓ�5#36ʘߜ} }�}>�%���{��N>��N��ج>��������}���;��E4~Aȁ�%W_k8��C-�%��J�e��F��hd��]mi��J�gd��i�4к�Cf�������ݖ���Ǻ�S�GJ=͜x��Y-<��c�p
.w����+mV7#����R<.3�_�z�!���~�����~�؎\���n����șu�Wx�5ײ
�����e۬bdI�ҧ�k��+A���e?f��sVo|��K}������>����[7��J�����LFs�HB
��DΌ ��0'��8 m��'8d����_a\�E�:����Mg��.��,����͛�rn�Q:��B�o}@b�{�R@������/��D{(d�Y|�u:�8~97�-vT8;����0��:��딍x�A�6��PP V)�������Y�D���ҍu+�7�bE�\=y:re�s0 �~=�LQ�}�2i콡w�����,赝zb����k�ly��dL���(�F�nZ����w���~}hn��P�_IdqNdj�^��_��ǩ�}��^K����or�	ٹ:v)h �alm\�cVňT���YB��l���|$ì�47�MS�ȶ�1sE���-Ґ�p�R�6�ɒ�x3w�؝���]�6�j�R
.�d��N��+�B'`}���9SC�.@��[�w�]}�8�]�7�w���Su�����^���,ʄ�ڻ=uG��6�h��~���h�=����.{M�}��X�u9�}�o�,yS[["�w5Ll�������
��[E�"�g��N�S"�o(�X���Ygd�>��-���q0��W��E�;޵��ƛ� 
ݚ�I���"�nwҤDvf��#���.�;ʙ^��H?};�w$���ȯ/R�����[4`�%��F��
��~�ɮ�L��d�
���
��-h��fGpuy�9��͗�����s�">� ��5�����|^��og��H(}����@�ݘ�X��D���P�ω���fq�ۡ[>E)YBq��_c�
k��Kl��t�<��V���|k��㉬ʣ�H��#��6z��NW�4�x��z3(���!���!��^ss~����uU&��)lC.�"e�-��PT!�:�0�#Y��jv��7gf�ͮ�(����Ï���r���A��F~��S��wc.av}��c1�=Mu���Uݺ�3��u��Vᮇ'�ؐ|���ގ���9,h��Z�!_��C�A�޿�����w��خĸ�� vA����j��_.��wq��t}�"ޯ^��똜:<h�V��e/\�f�x��ndMY	GPg��C�����]J��5Xeu:�cgFZ����:3��?���z�=�{��mb�l��/�}yJf�F�SJ,�=k�=w���B���@�A�DE�M��[���6~�#{��[�{�|����Ԉ�g�b̃���[��`����l���R������/��_E��R�c�f#nWD^.�$�xŜ�/����M}��>��E�\�ª`,��T�L}�P��B ;�i`�Ӣ�}�펬v1���6|:G��xa�j��J�1�T��b�rw�����w��5g���M��Dw��kܶzc�	��+����񭘱���L�p���l����Д�!�5e5����L��0D@�
��%�iK#�,Q9�g�������y�!��[Zn�lؤU�-���
c3A�X�vӒ0w��DN�1ok�t�@�5����q�� G*���:�<t����"�R�|mnv�3�tR>̼���hs�W�p�U޸���V��Y��>����8>o+���>����N��o+Τb��������:�q�~#�}ag7��7���"�+ޛ"���7ok��;��)����j��uv���E�~��~�2N�V�P֍4�?�ߤ�I/G�:����C��/ˮ��~�����d]v�����Aq�x杳UH���<��ٿ��� �>�"ǲ"zq'33���/�a?j��O�p����z����w(Fz!��)_���=���>\Lw�8�)��Zѷ��<��e��9@�x?�f�0�����D��G��<�I/GE���JM��+�O}�8��5��aPԚ���O���0��t�64k�Ofz+�����"Ռ>����g���&׻��p�[����9�7����!���j9�v��\校wL	�z��H������n�3��[�i��H�����2��UѤ�*����S�w�����U���=N1����{�#Vl��/mJUΛ������u5sg�T�pؗY�fW��X�8�T:��a=g���¦���{�]��n:�uuk����BS>���z���=C/{#�k�[�c|Տ]B��M���W;�ڣӧ=wG�t��A��/�9���y�^��j��}��s�|"��+f���R��'�6=��b�{h��"b�������Ε��o=�;E��ҟ���a�`}�J0@�Gtf@Yo޵�&k�F���6Eڃ���y��uWlvu��G<=���{�5�����ۮ��{���1U}i��<�8Fׯr��\YI|͏������O��u(G�'c���1Ɵ۸�T��5���ͼ����k�c��ﾭ~ӭ��߶x��}�I$�yϾO���\"�vB�ETt�r<�V�］x����R���+�w#�l�5~���|�XU��g舱[���fi�_f�������4�;,{��r>�V͇o�I��=5�N�p&?�:$��
��cs���� {/�D�z!;�Ve�؞�Hã2�N��������^.=��j���YE�фf5ut�M�J�m�`܈J}Š��O�}O��Lޱ*qf-̫1]r��d�%��������*F��w��z���b�穈h;��m&��.����BI��|�q�z����~���/b�f\bsM�����/Q�����ǻM3S���5'g�$�J�-K������G�>@Okw����\���W=�'�`�u x*#|Py�6��@��
�^�:ۺ ��A���&*�ed�fnqǕ�wb-�nd{�?��e1y�Q��s��M��"ߋ_YB��[�X�*
Fr��Xz.��r�a8+}��{6���ebn�c�'�'��D�������nZb��j��y��v�O:�aQ;�}�CpB��Z�=��}V}�,�I�wx��+@��
h�M�ʵ\>�Y�.��n�ʳ�S�<<���qy�{�"=�޲o�P�55z2������e^�r>�NEp�|}�1rs3�5�G⽫1;�<�,����\��NX���,a���fwj�C�.M�Z���fӦ*n��f[��A���F�[վz&9U.34u�闕|�i��,��O2�{e̲6Jj*�Y�EW-&�3�(����J]�7b���v���t����<��Bsi�ga�9��K�..��ounYivC��7�s��CK���)�m	����a�cʌ�NU`:E��n�T��{GmM��� t+��Bkm�7�j�NS�����~D�π��r��n̣�{E�[�ʷ����x��̦A������x�׹�G��2kM��������]	΂8�rt6�sN���Rr�A_qŻ8�tOͪ�!0��C�8��@B���ݵŸ�kI4x�FXlj�4g��4v��*��Z;JU����pW�Ս
�Qp��8�\)����J�v���qYss�k��$x��R4�ȰcL��Z��� VV�(���ŗVp�4i���c\O����+��s冷�̅�沺�n��h�˧����A�9:�lPKD͏��s���>�>�UM�;U, H_�	úr�x�D՝ĮaX�����i�mΏo��S�X:�
R�e�Q����'1w:S{��ZT��6��xM�yʖ����M�X�S�5>�˹PN��_9�Vd��&������=�tY�d�RY���7&�˧Y§gݻ��'mT��6�]�@���.�GO("�M��BZ��轡9��y�iɻԉ�gA�/s�V�4f���:��'{�ޑ�F�m�!vVX�ݹ��f�C�0��z�=��u�	ȱm���˝��wQ�'����{�+r���˳��ys(�o��Tׂ�J4FJ�Q���Q�e.��;'f
|q�2�Wxqb��>L����=�|q��wa����A��A�"lV����r�W�Eϑ<�ۏQ<�Z���u,:2�0��j��ґ�w14�L̡{��T��]�7�)�q��ˬ;ܭ�o���爳���6�\�Eqn�B���n�,���|Fj �W���K�	����;uK�[0gj%���n(E.�!у��\o�2�J���z������5���f�����4r.����t�D�:�۴�-h$r�\�����O1�+������q	�	��2��v�H��҃��J].�����;�7a�A��'p�G�y�����T�5�)M�Cu�wb�� ����|���C�\1i7o&ʂmd0*l�4�͹uj�d�\Ar[@^q�Owj���1���,�w
�m��W/�*��ҧsX�����N�\%i;�Z�3s�Z��t��^��v'��M�霃�=E��f ykt�؆;�sa�f5۩��2��"i�톝��Ced� �P��F㧷ٴ�oPٹ�Ȃ�Y��l�f���ӌ�9dvDS��<�8���Y(v�4��+9��;�km�q�m��[9�Ǻ��³��iy�aX�T��/l�x5�=_��| ��/��:(0,gE��X�[�,eY7M�؉�V�ʀʝ�{q0����AObp�7�{bV����-��'4]宬�h��uد��E�^+����g��Z�a{{��-�<kV�<N��F�����*����� ߷ /f������Q�ny.���X$;���B/GvXm��-^�X��r�c"�٢������imrV}�c�<>���2��2��|%j�&��6f�4G�����OE����yz����څY�A� �3��֗�$k�b��_G��.�o�{�YO����n
Tﲻ@Y�1�g�+�7��jΫ<�o&�x�c	�NTx���g�P�To�T<��*�lF�B�x{@��ë���^w^��*5p�JsZ�*i��ʾ}��k�d�=Z�ފ-��~ݾ��G���+BXؚ����uF̷k���)%�>�CZ�V����U��!�Y��Y�%��8����F�=�h�IH��}��ﾻ���}^�xS�vޙt�gur���oF��a����0A���L]�����N�}38]j��!��úK�ɱ��wPY8X�Tn��Lc*^\���� �����Y��-y���cl������!;�����=��F���W��u&� �n�����N���P�:׷/������c<=�]����q��h���m��U��4�*s�����8����^3�Az�羋b�=	}[��.�W��f�\�/�X��~�}�|5�o���^:�sSw��6�R�9ˮ{3��7Iw�+_ m'w[�~R�������Ȉ�ވ��&�b�}���ڭ.M�#U�֠���� ?8�Gsp#ߴ���:��
~�}|)�#>
g>��y��0W�-�M؄��nPC&mٽJ
�s�ksj������%�Y�y��*�(DA�U�o��{ޭZE  �W������b��z�uV[����}���"��h�Z��\u�'x.�M��1Ky�S�˔��$�HW����5+0�
��AaX G�O����jK���m�C��vnb6j��|�b��E,We���,����WS���NdC�F2�6Y�1��\����n�2�#Sw'l����jS�;���ݵc{��1Q��;ѣ��}�;��D��c{v�]�|����~�w�S2�^&> ����.����]z���&s�n=={��3^2���y�y������_\�L������9$����������hrBE��Λx�W��kr����,�U�����Q�ľ��ۊxQ�S��uY��<�\��k�*��H�_zx�sk?U�ղ��J��Ʀ�䩲����sӴ����_k�Ұt�g��~��=Q׼�C�]����)9�&v_*�'���s����������P]vM��'�ۼѤL���Ń2z�N�d���Ub�L��M���N_e�ת@�ܾ����md�T��Լ���� � � ��g^�.j�贈S2��>��:��)f@^ޖ��aQ���ү��g��$-��Λ�W7~����5>Ws��ւ�ye�#j�����4�['�N�p�7.�޷�߽w�es/�Yg�gU�I�4��V���4Ɏ�F�nT�6u�ֻU��.q�+�v����uX���b2Fa&f�f���ān/s�qİ�.���>�~+�5H�tx]c��bC�c�ꚉ�7A����Tu�{�zc$�����^~r6Q�o��b}�n�]���Ȋ�KM*oފ��p47��u�vϳd�Re���g�c��o:�4����F�F�ѫ��������m/���Ҵ.�G\V�4���wR��Q��[�.����]�g�=�2��sj�����_?Z�� ����h{�v��,�����G}�
E�<0��|7n.̚��}��K�����9wퟵ�jK����y���:f�iI�(s9c+�h�_}��n/�\�dog�uY[WI�|�o�v��^	����Np�����'��b��!?1/����:W��>:6���fr�7�k�b���MŰz���=�\ܫ�ޟh	��7����=Q�CtՌ�J*o5�M�Ұ^(ܵ ��L�j��Q8�Euy�ޚ��o7ǆ��ڸD�\�8��ؗM�Y+8��_+�Q�U�/BZ�;�s.��#�.r	ŊjR���v`�Y�˭��<��}���ЬgtśW�T����U�W���n '>���ˑ^�O,}-�xg*�\�jv� �rLJ��0_D����G*�>�^%�qG��\u�T�h9�Fzt�qS�W���n�O ��yB��?]�}�=���Ω	��)Y('�����f�\��^�k��I\6���^�u_*Q�o�:�s�G�϶"}�l����֟�^�u���X�f��k��۽L�|3�`�����.��_x�����R�?	"�?��m�Ϯ�Ҕ�$�tB�����H�f��c�<�L>��aym�y0�mτ�.�܋������cܳ�a�ŋ߇�d}�9Q�7<7~�����+w7%�V#�9��bk�;�B�(�7/"���pwkחU��p�� ������:�}����R�3�F)��P_F�v������KK���/���m����@e�L�+HQ��n�;y�p�7��`����ol�&�3{E$�HS�66�]�{��w4��a�����Co�6�I�IX�Sx����g���a��D_s4+F�9��c+�6{������l�ؼ"������ъ�6�?%�-���r�,1̴��ᨏ���>��yDC�^Ǳ����ԑ��W�g���欎�G`�%ӆW�S���O�;Yq���Ev��
E�N�QZ�D��[��G����Z���Ի�lB�v��?����zo��("��wS�y��&ԍҸ���j��F(ou<{��~�,�H�n�U>�Y
���@s9��,������>�q�sð80.�ĬsLs���&��5z���,�.�p_�<�!� �/ơO��O�1�����Q��r7W�#Ź��Vb�����8Rf��œ/#{~�s��U�]ǵ��r<��н���펊c�#O�ocuMS���ʇHzq��[>�u�����|"2������p���_+@���k�9�s��������z�:���7(]�k�J��Y)�|G�[/�b9��|.=�O{��/��T�7[72��L�.��Z�)��v���9��1�1/��C�+�Z5X�G�C��û��P�|�-��t���A�{�֯��9��UQ��siv_����=/�[4w�K��zl��9��
���zd���U�;�?~��=���o�6-�W���yw��"�\tEܬι�2�pj9T$����^q��#a�� �չ6���ҫ�/�c�����0�^�����}4�[=�A=ˮ�������;�P&m��I}ҹs/}��ę?����#�]l��K��T�X���#w��|��L��ʡ���s�Ν��V@^�����z���w�z
���!�E�e��/vA���F?�Y�'u�������c�g���z��O}W���#�K-!Y�۸p���J��1��߽OΗޛ�r��?S��M���Xj[�zN��hUք�˼L�H��GK���#�{����-�z��z3ڃ�B�z Uȋ�.���	Kr�|&-fD+
�u*E�q����F�H�P|"'�(��5k5��U`(��%�h�kWں���{����l.�'8(f�O{MR8��t���qɜk�MA��,�yR��bW��>�ͺw.��fE͎��7�v���^��;������f�vk��xM0l��Dx�Lc�㮾��~����z
�ʴ�|+�6I��R�Cu÷�B�	|���>�=�C�מ��ws������ZZ��Ͻܤ@EOx��y��-�5v�.�_Y�r^k�����t���P]}ܪ�u�W�
=�;ύ�����6�QŰ~��+�1��|S�^��]���犑V�������~v��R��~gd�w39�0m���/�§��ߦa�$64t:����P�]*��{�?5�V���V����� ����˭��UMB����F�8�ݞ˫��q=�o���E��$z'Pa]�MuJ�g/-��{JZ1]}��ttuQ7��TO���~��_�;�Z��3��w΃G����ژ�'��NK|i͏a�o+7�W�0���d��_6M{MA�{��w��Í!{u��9��+��[�����v|0�ّ3+nIPӧ.���<��� �a����$�mM���Y��5���}W�wj��n5��H�w��L��:F�V8������O[��t<Xg��i�y҆gm�}\�1����{�a�'�x�z���gp�1����h9���n��.�~9���{��N�0��O�x}�}��Y��_��~�ފD}��zrM;�r���MW+9�_��[�t�$��p�O�T,r���PX��*>�����Cr�$ǧ�Wٙ�tz��r��;��@˻�ѱ� �Z��1���i犅ڙ�j����D@��;Xo�#@��#밼S��5O�G�Y�h�ؽl e��Y��1V��ڠ�&X�[��4�������>A��S]�?�?�޲}��%#.�6�Ry��i�r^���cv�_f	�jf���=���
�@�s�@���u���X�e�*>�����zr�oQ^���+WoA�Y������O0{Ü�������y.��{4��f��ۄ�o�,�ηq]c�c��g�p��O��7B�4
��㋶����5�h*�3<�,�T:�r����8���{�<�+vGs&q�7:6�5���.ML�������2h�y�$b{ԏG:�p}ڟ�4z*������w�!O-
��/a��C�a�ٝ��k��q{w\糺Ɵ���
����ry�*�����nqd֥OUB�^԰��P�t��=}��/
���K�^xM֡���NQ�߷L����W8m��\p�g!d:�k�}��?{�%;�Tf'!Gz�٠v�iult�ٳ͘���j3+ۻ[��쇙w6|�l���G7��7Z����/a����C�N *�~?���͙�5����`�	]ﷵt���p���s�R�k���^(�l�_k]�+To�>�9�M�V9UL���)f�_l�c�˅���v���[ S��9q#����n��=�j��/��n2���\�� $}�J��I+�L(�)�s����S���uGx�ul��|~����|/�'Q �� }���G�\S��ܪ9}�d+'t=�ڒ�dV�:x֥�i�J�Ԟc6n��U(Dĝr���D��gmvs&f^.�i֮"��[�dc{��y�ic�����o"�}�5�q�r�CY���eT7X��{�@[y����u�z�~ó�BV�� �e�_�6�<]�hA?��W5�T_T�X��Ѓ!�w�ƻB�� o9Ӷ5=�ƽ��H>��-E���@�޼f�.�`x�4h�2(�����+���pˆ|a%H��Md�F㉇����8x	Ś�/0^�X5�邕jN�00ٻ�p$����#�^���Q!�EK�qP$���:+��1	���ZpvtJP�^:n��$��#8bh��|d!$ �f�N�졼&$�ư�=�b��gi�wب���s��\h
��OwKm��9G���X�z��x�9��=�ܫ_fZ�y�Ulۆ��kSg'j���Zf��d�A5��_ PZTP��0��]�Ww7�X7�M	���ょ\:��(<Aڇ9�$�|���ވ*K���e�H�G�;�K�י��=��#�E{��=���F�煊b�w;�$��Sy���o���{.�{�qg rħ�5�V\���['��S��a�w�9ʐA�B��ǶGNo'o�����]��u:��ܼ/������X4����' W\��{�vbŜ�ا�+^D^U�����;;��o������Vw�n=5�t�3����߶��2fR-Q��a�yx�zo�!o`b�T4�_Y��5���/t>n���lm=�w3��z�.��%�{�in�	����:ڃ�9(ZWq���Ba�*���.�wU�%����f�=\��U�̃ �j=��ʱ�����ή�׮�	$Lm�yd;R��z�hz����O{�K[����êT�n\;�jG"�fڬ�v��򶸊h�S�WMy�GLqf˾����s��ol	e�[�.f�ӫx�KI \���u�2Ů�t�;Mw6sJ�+�Ej"/:��F$�$�tn>D�1=����oI�o��th����h����s.V�$�Y%�ģn�6���q��+����@��mQ:��<Z���frx�wN��J�A%H��O�*�7U[���*f�o���-2�c�O3Ll;+��D�>]�jGH�v.��4�k7�j<��8)�3�,Ӏ䲍-���ʔ����v-6n�R�u�n1�n�}�wic|������F.��x�>؍̲M��kMm.�����JݤS���V��8U��ce�J�U��!m�|W}��oc��P��Tc��,İk�b&'WU��:�jQΜ��l-��-'Cѽc��Ŕk�ؾ�IVd}�M��7I=3����ic�ۗ����@`�����9�͚0虧z����pT�#��q��� mK��)����+cs9�ؙ�N2���ScY��$�t0s�T⃊��s�T��Xz����s��`�c��f�;4��X�\3���D++%\z~��o<�{��glZ��}QC�L�EE�>�8*��߶��)�U������>]��D����=�������j�"�s��˷3b�����p���4.�O�Pb�_l ���Tk����7�ٻJ�&��S3��;�J��F��B�)�t>;'EA��J:!���ݷT`h6"I�84��e�Z�>~��lU�{Q���u!�Z�Q�䠾��ezUC�q���#�`�'��2b_��"��ʝ�"LZ�2�r�M���}������țuݲ[��5mh�F��䃎�*"�VTt�j�p��G������j��^whL�q���q�����������\]�ă�QfTNp����	>�?  �[�̞�C���6v9	*��Ni*�슁n�៮��I�5��9��^��xu��z�r�]/Va�k��)��b���~�~�[	��A�S�7N�Nd��:P y�,����ҷhf'�?TH�EPG�V���Esn����`��X(�¶k5ߝ���K���0cGE��t�E��#`\��;�k6=|�N�(�G7���y�q���mF��}�ﯴ�Ūqq��9g���Ӹ�N�R�F�mw	{�v��׼<����٤=>h�۠DYY/U�{��V1�:jO�1��=Y�-�:��h�B��C"��B}��g?���k�A��DÑ�4��wA����۽���!lHL�z��l����r����x��D�ˇ�PĿ�]!�a[^�M���'����~g#~�t���\1öQ�ML�)��A͘�Z��錬뾈�P�D-Gt�ڊ"�cw�˪W3P�ʜ��U9�M�4�9[���r��G�yw�0�	Q�f"Dgo@��a)�����Ouw0��@_��}��{'c��"ݜfZ[U8����I�����*:-��#������7FC@8��O��_`<��<hSOyWn����A,9Wْ��fh/Y �Y��v�ĺ�s�n$�����u(�w��AA(���ED�!� t�g�H�̡[Su=��z���0*�1�����L�1�p��x!�,sD��[�u��Pڗ8%��w}��ܟ{���||2�t��21!f6ͳO��3��cau3d���ħ���"���tN�n��wi�]�5B���V�d��8N��2=ѝ��=���-��Hk��{����:ɾ�Q��u8�yv�"�Tت��2�u�w"����ί�~YvŠ1V]!�U@3�VM��k�{j����+��+��8�=˥7�_{>�uH��+������0�n+X�= ���{2�/`(�%-Ӹ|2�����xTf3�S�d��n۶I;/�i�y�Ճe���c!@����zfB���碷`���2���y����!y��=_3Y��h�9j�E�"nxΟ"s~����ثT�	�;O�5͝WT����k�"9�9SәY�[��C��s����z����FK�R
�����T�6F��q�B�X���i��Ȇ�gy>����c�+#g;���t��iyѪC�ۂ�V��,���P�U5���sX��"`�nVAެf'{%��셼�K��5S��~�m`<��N�|�.�t_M��;�v�A+�/Dyˑ]��tw`}��ʨ����7u{�}M������e5�fe]b�K/E"�h��b����.��1�d+�N���s.���h�CJ�u�حZ$3xs�+��e''_
GBz�{p���t��v&.������Fj_WV�+�6qk8��(gU`[�{���U��;�����&����W�N~�K\�ܠi�~�Ρ�w��5䃾��`�8b�H���}0Fֽ�#5a�gִ�tg���Z�����D�!P�g�6d����dqc�hf�{����.�A��B�W9O����xҀU	��}��Vv��O�=u���}^0��W�`��q2�vUS$t�aM�Ni�t���W��>x���)�vW����)<�|O������� ��b��@�"� }�ɣf�Q.�/�W{m��q��Khu�K�I�A*4L�IU�!N�E�_M�?!=������ܚ�{�ˋ&Q����v��7ƭ�*�	Ŗ~���E�&Z7�9ױ'c{4�<bp��G3ب� T�yN^hC�B�_�����B��b�@�ܸǮ�f�+�5+�
�~�aط���(<� G���v�\��hQ��u[����]C�ԽNl�n��1����c�������iq�LK�Sq���w�oټ���w>�>���pTd:��HcLfӦK�����0 �h"�0~?���R�m�ٽ���9�����.{�h��K:0bSe�N�7,;�0�ɚt�����K���*��^j��������wE��c�c�V��W]�mŃ5��ҽ�謘e�xz���ِE1���n�`�J��ǯf��ǂ��%�)z�e�/�~3�:-fcO�A^H5�{��,W��Zn}և^��]�b*�Bva��|X����u������.%҂_�T�Cz.�D���X��i���g�F��~�����8�YӏoÙh\"������~���os1�݉G��G��~�%����B���!ͭ�	��)g�
u��+� 
��%>ꛖ�=�'+�L��[��!��2����c.'o��s_C���G3G���en�~�LS�b�&R�v5�a��6��~���p����][��p�m2~��T�k�)�Íeԑ�%E��B)^U�H�o���:��s*�ǧG/�Q��sim|�խ�"N��yWr��3֟��[al}���׎b<*/��a�@/����L�����"��N�#�>ͪ��rO��b�X[3��TI�
�*%�z�:fl&�"bI�$/��)�Z�k/�����cu��l,W`��XL�����ہZ!5��s�+1���sU�"{�����k�[7�9#�,�S�Hp�v�p�.�0v�)z�]B�!w�Z��P3��F�AG�y���I��t�5p���~�y����4�fTxxr���D��cp����/=��b�4#�#�/ft�{umv����g�ƣ�9�/��������,g��&`j[ILЀ�q ✧�(8�~�g�-�w���,���L�����7g������k�\���O�}��Χ��W�Ux^H۞�<4ؓ�����B"��%�|��ǽn+{~�NF�uz�߈���j�l����L!�?1�9�}������WE�<d8�G����ʒ�om�=O�A��Y�5��а���e̍��`�c�F�P�˗�s3Z��.�os�����-���*��z�6z�`L�!�D�`/�'k����#�i*���!;q�-��L�r˫�W0*dx���)!�ӻ=�؄ב{6l�wU�:�	-���i����_]��O�5�f<ռ�s�s�����]WD�Y&���������nd�
�ͽ��:��K�O���!F�Q��֝J�CX0�T
�
1�-���6�:>8Q�u�1a�qU���i~�ڻ���F�^����Cq�p5�7�X���58�ytw(W�����N.��(�F����M	ʓ�:��8�����g�(�����Z:]���Vz�֒1sq$�W.:�F{�V�e3���M�$���|�</���^��IO���_\Ue!��N�Ž4�v�5��ڤ��8�6 �v��9����4�K*b-L����]=�M�Ӈ�$���i�kq�_�󶷀�}��׽�� b/g��{[M�^�Ϥ��^x���]�l%��Yy!m���-��/	��}��Ë���:�QL+2]����(�Y.N&����������gD3r���L�k�3��4r ���p;&�ec;Y�|8��I�D�l���XW��p��p��x�wC��32��]0�BE���ʘy�� Z�R�UfL�P���J-M%C��=�8�B��΃ϔt?\�7<�����v�d�N�&�����gp�x��dg�df�S��l�5�D��
�_�y���ї�J{��M]���X\]�`�<1q����>-��\t�tW"���W���w��ֵ�mJ`�W5��g�
 �H
�I���7-�r54pR�� ��ܶ��Ի�s	�2��Ÿ�'��*��{*�v�W�ȳ�(:�/�%��{���d|>D��+w��{�Řb�=��w2���gb���pd�^�Rs�u���P�
)��Ը��xqЏ��[��B�g�>"���ν�c�-�٢0��{��x��������eeӿ��#E~{3���û'?a����aiǺ�D3s�0\uUwZ�l�*�N ��D�B�ﾚ��'W��9�������׍��in�r60�ځki �-�h��Z�z�M�ة�iTnI�֬����E���oŝ��/g�<�^���[���^���}�	Վ�^��Fy�J��w.�/#�}��(��8q�����}�����G�=����m��#o�%�B��t�_�}7%���R������Cw&Ft��o_/C�T�LnNX�e��o�গ� w���Lo����ijrn��">�y��]P����f+&���F��g��C螣��J���Z�/���aG���F��T�
����{����|�v=��af�.���z�v� �S������Źض�l������Z=��v�����u��k6%�¸N3.��	�OG�j��.ޚ��<Z��[O����>b�"<	�Է����c0��)M/Օ�L5����_���{g�^���������8�eG�\�/�!�ˣ��!~-�}��;�Y��g_�N���v��H{w&$��	yVKTԈ�a�>�6��d�Ot=�O�\�Չ�����R�.o�	�pA��+ڍb5��rD��XɊ��&���:}�x���~�[n�q�Ѡ��%f��H�uHjv��5J��^�.�X�͜���2��D���OV�����P�,�ܭ��|hEɀ��*�$�:&r1���Z�O=y�zN�t���s�޹���t�w?e��WAR�u����2Ku��k�����G�ș�q�a���XVt]j�)u���2?y��=��ŉ�i6}�?��>v�j�Jz�+�q�9�==j��үͬ�}��_
��G�������S�0,��?m�;��c����W=8��]E{8W�������Q�e�M;��Lܱ"<._l�f�ª��G�����"%�#���XB�CN&���k|�%���ͻv�,��|�yn�G:>5���'���e��*N�zj��Sv7nˏD���K��â�˻�ز`��3dr��U�Z�{9�/d����:���ZUi��������hk]�R�d䪨�Q�^EHr�\<�/=���qp�'׾-X��#%^�91*���	��Y�b�`\o1��P5{>ý�G�A,Mg�+ߒ���8	�t��~{���YV�Gm��2�[es}�,��v�S��\ۈ��C����ݟ�Ȏ_��2Uq���V~VƊ��aTV��x�(�;��i��t+���<����ʌ?c��D���n�.HzB<�/O�`�����)�er��W+�UT��_ݖ0urI�s9*b���)�ϴ����������Q��z��*�7�Rh���������6+)AZ�9��
3�'�[�z$6��6қ}Y>"�T��&".�	�Td��[4��9�-��Q=�{q�������V4�L�Hޭ��+�G{��QU���w[��R��ֽ�����}J>��3��쥵�r�r -n&I�ǆ�I����g�`[}<OG���$R�_ZׯW�������oY �,PJ��se���5)��&���H�ɫ�CYD ����h�}YPX�}R���oq,�.>�"�|-X]ٰ1kD�=��H��c���K�º����)#����U:���!�^�Cl1�	��Q�ٕ��]u�*�,}-cfv@`�X8��{k:�0�&J�㠮����v�ӨMJƋ�i���t-�ЇC۹��$E��eb9�c�����x.��}:�5����7;x������k���G"�R�s���PA6b5jn^�rr���뭌�ƌ�ٵT�_��X�T���&u�9��͹�Y@�d�o!P@�j�0k���o���5�e�+f�V4��h~��;>?Zy���`ʗ�f.��JLU컠��C�>��b�����dѶ,f.��� H�JU�%E_���ݺg��lIS墒��_[=\��iV7e~љK�|����s�ky�����3̅@Q��m��RѺL��f���%)R�E��,c%j8��f\]�f�S��7�t��,�^�p�c��A���\�M8b��+��e�0�Ӱ*�B��I9x-ng�L��*Gw�%��4fc0�lc�E�Pŏ{yf���ݎ��t�U�l
�ٽp���7���4v�t�e���[�5깅m��}v	�n\&]���.��<�=�� �)CV���s2�f�������We�šX�K*�Eb�Sjԋu\SK;Xd������]�Iu�M��j��;ήj��ɧ�Ee�O�B�oE�f]�K�6�H�F��X
�uh���.�.��8^o<݃\���h%ÜŐ�o ]y�Zĸ�n�j��9�1��A�Nw͗��v]��рh���	Gtb{݈�Yk��=ѧ�[�1���e�&����� ��:�v�3f�醅/�F��v��|�n��m�6M���+7�B��m�N��oY���F�����ޖ��B�i�ٮ��+ga'G�"{�N���<+����Y��A �ZlJ1*89G����\�3�����(�bG,�q�
�Y��6����zsy��4����{t�R�i���[q��8��n�C���{ύ[�v3OF�d���
�pi����#������c�����u�ʳ;Eܽ�f�̨�t��v�;������e<�M�`��m�y�qܧ�8+E۵{5*=w�ն�RreIl!�\ӳ�׍�TsڟT}�
Su1���͂m}}4e<x���p>]`��7�)��|-��"9]2��+PA?�L��V�2�й/w�1U�)s�z�����Kc��WYMjj�y�ِgm��	����x�W[�bua�]tto�LkWl�����-�� o�*JWY��?+��#����q�$���Y���qV3;qC��[��Lg1�E��*�;f���c�6P�j8�����V���V�ٸ��h�٨���\D*��|\[��sƍ��E�)赼gW:Ӯ�Oo���U��7P�=��Bє`a�7b�aV��A8]1W��t�^�qu-�p��Rì�Q���e����c'l�}���/MJu�Q�����*�}�i�}���^i����q~-t�9�}�}�����[ȧ�RI���<o4�׫z3�U���%�O=U�f�{�.KU��b8���6G�1��QG-@9�sG�]>�m_}����lzY)=y�s<��e�N�=�*������+y}��X2&ɺ�8�s�ɣ���
Cܙ��;ub����ڐ*�ci�N��v<�WD:IoD���;��{=J�Y�̑�����uf�FJ�R�^��*�W	��KK^g�n�s
��0#_�lך`�U�UA��GjN�j�~�;%�!�g�o�}F�X�;6�>]˰xj��ѐ�����Wb��L'}jU�.jOY�~�MǍg� }M�{�޶�ɏh;���v�I.q��\`�7����������U3��rj.Nx��u.�H"��BQ��'�	��z���F��w��o�6�AL��w��>��;���_PF^O���
��3�Q�����qְɸ̚K	�)k�T��Xfjjn3d$*BIm�'7��Z����}�����ټ����rS�M�p���N��Q�e���4۶xi�S���w�SR���hּ�l��@�/9�qQ%0a��hr�"ub��!:Ny���X\���
���jC�eE�����򓞗e�`^�������������T��B;��qd�-����ܥ�v�b�l?{�G�Boێ�/�?`����fw=9��� '
���9��n��:k�˿�Y�D}K�)�ب���YayN�?Jg�.�<���ъR�n����;��K

m1��9;Bh9�C�D��2�2(;[���b+����e���h��}��}�������	�t��T����6��<4j5o����>*.ew�hG��fQ 8�<��<Mmm�\��$��D�zeGX��m�G��ƕ2��A'͊�>�M�F:*�R��!4$�4���ên3�|N��~c����=ٮ_{N_?i��§8�b����y�.��>�����ӷ�!q�<�9ˑ�����O��٭Ձ����"��YZk�C�>����
�LS���8F���;)Pt�7�mw��Tt&��e����<�[�p�5y�I2m��.�~�V-�UL�M�N19��ܨ��p-�9�i�v	Ҵn��*AUPb�+�ՙ��
�!��˾h�J� wZ�$�yuk�oq�ׯ��V�h�����U�Y���'l��]�t+��T>-��9���'�z��H�J��}�ķݸVG����zș;�d\�3�)]�6�hI���O{p�/�.�����p�����1����֊�겠m�^c��mҢN��׼�99�� ��a�]t<�K�Nɳ�b�������|>C���kXD�u)}�������;U��7f�??�>��Ó���<��LM�]7���k��Q�����{�P;��~�<Lx�.e[��ԡ���˩ի_^6�)|N%��j�
����z�����C�WK�H��{���@����]���3!�ׅuN+ ���ìu�;؟���~�9{v=@}D�/�%�b��Ay$v�h�?�D�����-ʍ��|d��6!���+\l-���o�P�a[�z2&Bw�H����I�ȷW�I�]�WȎ�5���M*
x�X�w:����]:+<��]��H���w/�X��e߱�S�ÿ_�˔��&�%P��m�>ڶ蜽3�y`[9����ڰ�;u/���Gj��H��x2�ƻ���b�R��Q�da�|9,�vR]*pf!�e)��Ò.��>�cF��=.���l�dW��9�z~wv���"k��D-�Y^������ݾ�>%Xc�]2�Qq
���ʹ'I��w}7/�a�Q
��u��Ȝt��8�LW�3�)�n��1��Q��O����hGg��`�!���Db�߀��=R��f�Up��W���i���r�A����=#0-�"޼�,H��WYyuo�E\[����{����FW�@�Mv\A	�[��Pi�����Җ�Z�~�t�b�}2�I�zvC�H��|<SF���^	����̇�θ��c5|p��}p���Y�A�.D:�W��]��y�h��?R6e	�|����}��=@h��$��]�����
�]�����N�\5)(g�{k��ě��u���:�9iO37e�&�eӨ�^�q�C�Ò{��ƹ���Y[^�bc��l�0fە�$�܉����XG=C��iŤ��K����ǵ��*�:B�S)�
���y���� W^pw���Z�u�']yE��f�$�&>Qg(�AG��[�ƻ9��s�U8���ي�<�Se)َ*�ę�#�g'�O\q�o;�mb�͚�	K�����l⮆�b
��cl���,zf����#���偆^����㒖��x��	���4|�`����9֫���?���)�H�� <���m�s�bX{��������.��
Ś��\E�6=���L���*���>Q��7���S.oK��F3��$#�h�d�9�n���_[�:�3|���?>�������ص��~)�Bb�1�߫�d��]3���A �:�t:��ދ�}�=�ٷ�~�rv�sT'?��452bܦ��+K�Y�7U�a�*��d&���u�a��#�������i��K��ru�)h�7 �}��4En�L'YI]�{5�������I�u��Ey|�j��ߨP6�s�W�uFZ�3�(	�U4�O{n�:w����F�Ç�z�\�.�Ia�]�ye�豻Q���w:^�MO�����ׄߏ|b�Ӯ�����Ld�y�.����Q�z���;�0]n� �͋N�ӽ����d�"�7�� x�m���_�,�Q+AD,FA��b�2�n>�Dj"�{��/)����g_��g/2�Ϲ��&
���yO��9]��t�ܳ ��A�  ��6��a{tN�y�e�	sV�;������T{��1��lZ&����6���}�lv}䧯F�0�{r��li�9���t͆]p����/G[�t'9���KO��Tٕ��V�ɘ��ޓY�;6
����E�)�t��(�YY+1X��Lrw��{���VG�h uOn��]���������U����p��ߒ�[L�����L�)�}���Uy���Q/��#|^w��O�.Qh2)`Ev�oW3>�>^D���*K�*"1J����q�r#��R���I���`����ϒdT�G�}���Ԗ�=B�#Ы�b�;�a�r�d����ɪ���t� g��5��ջ7]~&*6/N�1;�0
�l-zV���M~V��cNl�p��Ͻ�=[�v+�e[��I5���\ŝ.�Y�O�+�A�}@ly�L������������F'�)�K�h��y�'~j\E,'�k�Q���o[�g0���7b@l�n�x�U����;�Π���2�c,�AT�����t4Fx�Y�:sR���3��<h��`W�],c��7�h�&���ByB67ɒ�A:�_wCi��w6��0嘆q�-����w(��`�ޠ�P߭�ξ� ��x��{���9��x6wB��IM�%:�6����{d�.g����}k��ϭ����rtB�B��#��%��h���s�p:��A�R�ma�_
��S�����Y����u�ޱ�I�hz�
�t��R��f�|�@��ċZ�a��^��Pê��~�&]�ʄRR?���c>��.�=~h�5����h(f�OE�tONIG5��޿B{�C�G3�H�iz���k�-	�xu�E��N�ؚ �yta��eY����ֵ��j��9���H�Z�X��	<�J��$K~�'+�u @W����0���鸣%�zOm�㼥I�[90����!��ZZ��?z�$�eyK3W�gs�m��ȝ�Ќm�K)W�}hUm������B���L�=����9
�(wK�y�󼻪����iH��ֿ��WK�J�r�����><Kº��>%����n����-Q/�:Yr��Q!gy��n���W����v���tz�[9zrڵeG�Z�v�wc�����ꕏT��Z�� �9����L��i:��<�:�ـ��.Q�t�ܺ|d�:I�c�Y;qk�.tw+Ǝu76����T8�=+��$�R�&N�Zj�yDw��]��VF�~���])�L��N_��Xɞ ��m����&3T�{�x ��菾�=�[7�aN:DςdE�ߖi����?s�yG̨[�.tM��2h=��+��~U�-�S��S�SI�}���G~�Os���%�����[��%�-��Z�r��\Z�
^�� I��G(vr�`vt��NF�]�ב�J$����G�i�̽@櫯��?3ǐ�r��N�l��h�M��2�+M^�ٚ������S5���{���=������w��x 4

���dĨ{j�X�܆e��=�*��k�����37E�BۓK�p{� �!SSw�(�5p81J�ףOMW�V�����EM-̴�2���i���#�y��!œ�t�H�>����D�(�t	Vס�h��������A;ZZ�<�Ћ�~�7�����7���ǉ��*�i�����On3�Y�p�hg2��.�� p��G�p���i�4�{�u۫T�\�>������
�9����a�8Қ�Oε{��š�	�h�\��w,=�ǩ��j�\�T
�[�['�vʺ9�r���uK��.t�L��0Y���S�f���LT�x�HP�ٖǇ�ނzY��ݡȽ�NL����qEl�{Hwv��C��̌���>{1 p?���1��J��*~tw����}�͝ꬴe���aW�����??!&��9�� p�]�_��F��c=�ȍHyo ��M�a�{��J�kP���7�<����h�U���[��׾�7�n�6�|��y"닸��z��=��][�k��r����魱5�U81��R�3KM97�蔍2%�"bn�K�h��*�����nmf�}�[~f���v�Fl�Y,҈.��[�g�s��^��8�6]ȟGqՈ���[�c��c�Gdڥ������ECrø~�� 9Ȃ��5���ލT�9^�+�1�Pݳ���\�v�[�8�%2�wj腝Fy��I���1� ��\����f��
��նs��`'T��W���1.����E���f,�5uz��� ��=��ˈ���{�jV�|M�i2/��Ȁ W���Y�٭	�`xf`��֩�VwJ8.���+�,I\އ��{��D"oc:���"��(.I�^�n����BV�k�4�ַYx���j�(���ì	�d�kI�X9U.}1��3�=wxr@F�nj�"LxU-E���� ̉S����1�^ᣇBQ�ǛT�tFY��5<H����f�VEFq���X��_:��Yys�T���ŭN9rؽI�鲽>�����5g��=�������mE�my}��$fa3�hx�"ozb{�.����򡣌7"(��FM�b�|�&,�Wl��+{�� |���"��&xV�*X�}�VMS4;F�S&E�����:���E�ڥ�;y�*�-�a(���h�ƜE��Y�{AC0��1�d	�>^�"�]V��'�Uã�\	�Xd]�}%z}G�~{)7�z��n�zmo9��Ԟ@�F����L�4���}:���W�Ə/��:�f�_�]�93��|�m������Ҿ:X'�������u�F��D@W2")��ݨ&�;��T���F�����b�S���PH�ࣴ��
�ە���n��C�uT�d��)��u۱�ӈ�>�7#��
9�m�A���8�>��2)�ԧ��kr.�z�	{,S��E:i�(4&Yf`p��Qr����e�(�Y�%p�G�[������{��>�������?��!$��!BI���I ��B	�kB��$ ����C�l #��
HI!��$�ń�	]���� HI?���B���B$$���|������������?������!����?����p~f
"ٱ���[��Y_:�p[�&���k-R�(�'�I�;��R�)z��U�S�.�h���Z�T�ƥk�ѭ�,�s�Gv'��J�lۇ+;�Dҹ�R�oQ砜#�	������7�)i�a�oL0Z�D�ݻ��3)-�.�c,2�ly��9��Vv!��9��&���"�'�형�Ĳ����n�P�zvΪ������l���1b��ibyH�������J7�-^��ٌ�4SƎ���̺�U;܌��ʭ8�rcyW��G\�f���,R�����ٵ��e��MV��(�s �[+(�,(&VAL�NQ�e�G��yz�jQ�Ke\q`*�\Y��#/&֖�"�T��u�+^��������6�MS,�X+3Z��U�L'
l�B�xK:��VFP��
P7���]�u��n����qk�T)��b2��P�ʬ�nYX�6E�d^Z��w`D2���4�F��:�7I@�ǌS;�0ukÛ�~v�LreˋW����$v`���9/ T^��G��k9����n���]��E��#l�� -��R�^fYQ^3!ٝ�i�;��.멌���-0�]��������ɗj�v���	��CڑKc͡���Sɛ�SIV�s �@y�f�+(�F%(ۄ[�A*��o0C�ښk\���)��Hr�,��N<ثQ�Tm�]E3h;�o�
��A�(+Gi�ׇ,�n�1+"�c�x��٣X��Ea&��f"oq[I�B�-T���$vCT�oU�Oo!9�S�D)��.�R��P-É��M�m�7�e��Yu�TN�$��4�H����)����\6���r�&�b��p+ъa�Z�f��Q�D3����R/Q�7WO�{kd�[.��n̬���v]x�K`�֑�U�sl��j�P���<�$�d�� F� $$� H�HF���$��		����0$# $� !	$ ������@����_�O���!$����?����� HI7���$$�� HI?����		'��$$���o�����4j�!$�>� HI?�_�o�� HI?�@��~�C�|g�ṣ�?�̄ HI3i�p?����߂$$��Z� HO{>�_�b��L���DY��س � ���fO� �`7Ǐ%+l) Kf�	EE�D�Ջcl�"�͍"�0)���I�mL��m���L�
k`T��@�͔�ɪ�P��)��@�AOY*�� PPE
$)�����P��
U Q"��@�Q*
�YUT
��*�	fT���v⢄� %%H��CV�D]�uu��
eN���Ү�Ӷ�l�c��{Wk{2t��;+.�u�ډm֋���]���w��m�Ӯt��Pi�إQ*T($qР (�A�   �L+��l�v�ڛwn����{v�n�6ش���s.ػ뫭ׯOMowuV�I+�Ǽ�����k�Y0��"��QE:�.�^���OJ:�w�ޚ�x`t�׼����l���9�ug�:5L;����ԯ ڐu�*�
@ۦ�{�o9�
�:�ݒ��vt�;�:U �'J���C��ݦ�[eM��w������ ���� R�w�i�����zPj��z�攽iY�=M�+�o�캛���	�y�s��ՃG�gJSU����Mm�os�z�mn��f�Tm��D�T��'=.�uf��^r� ��w�]��x9�yIR���Z�ٝ)�
y�Nzm5�p� x�^��e=�{Ļkf��@ �B�(����ކw�u,�;Ǽ������(k%{�=�)[e�^<=;�y�y�Zz���E/;�ޖְ�s:S��g��H�^�JB�
�qWl�ku��XǹEQ��9v�U{����IK���PAy�N����U�ݴn�������oO4�[A��	W��QUR*���mW�v�RWw��k)��̇{J��{x*��qnl3V�ü��2=�z)*^���x����;Ӟ���y
 ��P��D)/=i���;Oz�IR�y{{.��z�g���^sv����x�9�RO;��Tح/w��������͵���y��Bx��)PA��C
��� �S�$H  "����@@S�*�SM4�I��$�OP i��׭�n+� )(�@�Y" b�8�pf;�ϛ����_��� I��?� �	$ԁ�� I���I'��H�2BH�@���I��8f��s��ٮ�%�`=X�쵻���������D)���� -�����2���}}]v�����i ����j�--�Z�4+uxu�u c(��G�D�����$-8��^�WQ��z��Y�)ⰾ�j���e[�FS��d4:�wú�A������@bԵ8�]w��a'�D��}H��̻���c�7h��^h�@U�}��x֎ ^�v�M�۷���Ǝ���)��沬+�x��Ҷ�u"�+o�ݴ�`eӽ��wZ�B�ڮ�b�
�>
1����X"ӛ����y��w��﫻��[��YawfXs�f����E��v�sƏY�ye�]�-��Ӣ��vUe�Z3(S(�����藔M];�K��EA�1�-f�t�o�#iY�=���"�;�	�tB��.�1w���"���Z� �V<g����c;Y�׊� )��?ZvUw#I^���J�Li�
�Yyטj�w��w�`����evn�*��;�
�1gf�ٷU�w�w��F�^u%u���˯
G][F��k�o *˳���/n=��r�e;�!�.�ˆ���ku�L-�ڰoquG7�	qA�դbc��@ݑ|�j��6���|o��*�~ά���)���6;R���9���;v�|�9��o��g3|s�X�Y��ѡ k.���8��F��OI�mwp�O�E����en�e�d�u��>{@nn�vq`��j�zt$��/oڮ�"���A��b-cT<jho�{Q7�*kO4s\�/��ױ}ڏQ˭�K�S.�ev��y�@�T�R#��	�Q����Q��`e��M�� �<�]��<ݽ��9�g�����luYB�)��
f@a^���X���,[- "�7�xu��(�����x[l��[����F����u���0� t[řŴ�Wax�s�j�V{��!�V�:5���.֪$j䴪�ί���ֵ���}�t��D�֞�ZV-��u�ej|����������>ެ[w�p�c`�]��`�	PI|V��]����/��n��������Z%�ǚ㛺[wv-�`��;H���Er�ԗcC�: �ĕs���B���F�
��g)Q��Ǐ�f�u�Q�\,Q�:�^[X�YW�6�HݾǉP�Lf1v���Y��kfM�ޢ�x��.��o+�N�Q@Vn���VXЙ�pi-�B��v�X*��)�o�q5Hb�ʛ�{��]����믬���\q�U��FZ�=�9ͬ�VVmƱ��;͝}�Ⱦ�@n�|]f�T(�*�Q������y{�䴫�o��t.�Z�m��LK��%���A��b�Gm��I��7]ݎ9��q�5�Ւj�V�1G������;I+�]f���-�wf�v���x���r<�5�h*o�h|Y�B�>��+z�V��a롙���H��Kաm��Z9�I0Ч�+�w7xx`�֨_Q��H!Ʋ�f�h��\��t/m	���U�wI���.�.Ne$RC�Y��*8�*�y�O:�V��J���̚h]�'F��\��A�t��hԆ�V����[Y|sY5�u�����.���`�����6�:�� ��raڽ7�z�F�n�m���0P�+r�z�kk��&�k#X��t�j�D��Z��6��1��>��iݠ,wp��P�Y�V�l`���n���}�z���軆�߯E�=1�QZIչul�껫�õƮ��k����ވhw�s|�K��7��2V���O��D>��L{��i�|k����A�O�^Rx��t��U���V0���8U����Nؤ�sU[4Oqw|;gWj)jA�j�ִ�]�]�>o��������Ul��w�*�*��QES�z��[m��S�Ԫ����(��F���M-t73��Ճ�QvU!�@��_
m�:���J���Y��H�b�sUZ�mo:�l��� �p�b��ⷖ�X�i�}w��^7/�5����o��{���St7uض@������4hn�K�R�M*�z��!�ۻ�F��޺�X�әuû�l�o�X��Xc}��`<�	p�^�'���w���2u�ګ�r"�5�T2��ʴ��(]�Xܶ��i`�]Z�|�ӊ�e��\9����V�CsU��1��-6�5J�x�޶Er�Z��W�,��h�V��E�[Ț;��{��[W�ʻ:-�\OxPƴ�{ֱ��wF������t�Hݼ�HZ�̣A�� ��d���|P����Ho*�7=�����k��;�N�v�׹�/�]�ګ�`[�֞�+��X������g�s����.���U���U�A�'_x��Z(b������w!K���{otD�V�F�
��ѧ���X�L�����J��@n���]j�5�i^o6YM�c.kz��yOo��t�f��EwIU�:�!Lv�{�B ��|� hM��h�{�X��oQҕ���vQ�u�2���m�t�Gm!mp�ޤ��;�M��H-� �zpv��t�w��OF��xY�i��GP�C8xo��vR���@�9nnR|4���m�F�붨vziv�<�3�P�W��M��LU��+tQm�1�ی��F���jn��5Ν-ku��f�N�y��	<�6O�q[�ov��mYР���P�b�q�3�O�CB�h��qU��v�اk����xp"��uX�x:��D�S/�5�I�^�,����'kJ5��)�� �>�C \�:��o[��7_r��P�%��C�mv1U��@v0F#�WǜEQDE}[�Qy�\�k]���Ƭn�y���a�{�N�0��˜����=�����5՜m4a�w�|���L�/�y毵�AJ[��������3�����{��y��,DdDpl��pù�$��:��n����/Q�lYYu�m��`�����]�b�3[&��N{9�܊tIy�o{Go���9Nw����o^k����\�8j$Q�g}�xGz9����4����ؽ䒠��+W��l
��)VS��ްD��y�xu��壮j���{�Syɻ��&wo���&�%9뼷zw�5v]%f���]��Ջ3�,�6�F�+��Q\P���~��]���ꥷ�]��]�靻3+�҈����1�)z�}��&�3�(�훥tpw%F�����'Ĭ/z���@�:��7w�֩�g;:]
(����w�<h�֛���.��e�P�w֎�m�t+�]���9���\�X9֍��!!�9�'�M((��k�7����޹t�|��'G�7G�� C�h�85g�jL�S$ڪ�][|ָ׼��_]9�j��Q�[�{E+�KˤQ��*k��My�hY�~\/�?�ؼL�Չx�f]1ηhU
��:�S�_=A�����V�����֑ζ�FV�۽�fӺ:N��]d�լ�R�k��������5�]ֻ)�e%ݦ�2���X�):y�[z�kݼ��	u�������nݗ��㵭�p�^�����0ؚ7�=�|o�����Y��a��n��˴��g�`۫��N��%�]^��[J�b�X�n���M,A��૳X?X)��*�N�����X�4���c^�l�{����hu֢���w�G\�=��˫ۿ4�3v�QQQAEPQAEQEQEQAEQEAEPF"�oyw���k��u)�sA�8�m�s5��|o�_SZ�=��� �g}ӋQ(��*Q���iڔ�.=��oeް��E;�-L��F�/�IRS9���O6k��=��yu�Jɲ��1I�Ԁ��-�<$�o:�~��ant�[��¾�\��3~��Eop���S
aǔv�ksN�h�T>�F�H>�7�J�gY�f��p8��3p�Kss��GQWo�=:^�x��u=�=��ׯ(8m�S�6�A�������58YYS�i��{�mL��o,\E���ѳ��9�z�А�JA_��y�籽�T�1�0D���fp���e�]�^���v����	ለ��.��;�]k��	��@DZ�t7qg��b8YT���3�'�O��N����rh�1��Ȍ�b�DR",�P�R�P�Y�����]D��]_� P/�,�x:�f��������]^�G��Vկv^�w����]�`�#������ˏ3�9��u���*�ʶ�����fAmcY��-]��U��ǧ-�֭����h*�]��/��뀦2��L�[o�������k�gq�!�U}�n�
젊�C�R幾��w��5y�aވ��o~ᮍH�hymL�� �}YJ����b�e�O����.h��s.��z1(i��׼7�k���G�a�̵c�i�Xf�TT}��9�����f���^0��$�cyD=姭|���P���Z^]�����oi�%"]��35�5��L�L׷b:�p�)ļ��Ou�7��.�R�9�E�{A�ڻȮ{�k+��r(�U�`ZC�����;z4��5��rb�b�DQ�k�}�����gM��p^)�g�n�@b7�w�9�y�S�G9˻y�9X�V]�5��vqv�?R�j׋2�t�G�f�f�s\'s��[����N���%���6(�D�)K㇊�������z]�{N���;����^����u�k�2��J�%.<��^���f�����k�4t�W^�o�ե�4�j��:)ev�̰o��s��7�f9�Ǟ�|�La�w�ɭ�-���ox��X=�*���,�5b�.���8+m�i�� *�KJ\֍	y�hD��ü�z���t
�{�������x�������Q�Wj���k!�*d��ƹV�c(V7���÷u�˃�u����q��m�>
�hZ@�d�7;*�Ӯ)5�,.ڵ�MvwV��m���]�![�-�޻�j� ��QŭފT��)�"����=�����Y���WDv�MR-ݗ�A�H��]_����<�S���]�����u�����v�*�5� 4<Z�W_���خ���gZM*�z]�D僡R��6wU��T��^��%��>8V��zv5W@z�"��4%��٣����<����՞��N�w]���-j9F�]����uv:�k4��u���`?��=;j����]��Ҭ���R=��Ǵ��C0�,��,�y*�� �d:Cw�n�o�H��m�d�΅Z�75�:�k)f��yGo����$��[yw� �2�͔z�V�Uٻ[F�{�����v�����݂[[����B\,'�}�A0��e�Z��j��wF��Z�_Z|��e�\�P쳖�4;��س��]fַ[`�=��E.t�rݭ��qe��M��Y΍rcI�y���{�j����t.�tgs-�6pVk�vR����E�Y��L�����BƢM����*�Ӊ�^��kowpr���|��赧W����ќw���������ҳ����]�W�ѬF���Y���3I-�DY��j�O	[�׹�~��j�n�_k��Çx�{�\�;����h�1<k���U����� �o��C�uy����9j��al�?)���Qz��:���[i���a����t��l|3��ٷ�wK����;�B+I�C�AߍZ�P{`�<���v�uV���/�� ��>Ն��SW\��s9���ݷE��+�,�Z��Ձ��9��N���Y��5�^��Xf�6�d:VS3���N���G=�u����.Cm���8�W"�-<��yJ�X}���Z�{ü�,���Go8�QE��"�4����Ím�ͯw�a�N��kttW��>W��}O�R�@|�Y�k�e���>�#�'uP�V�WWuuWu�[��h�m%�_[�`�;DZͭ�4�k)�hk]�{�m�+i����;H�L�9G5mat�մ�ֵ]�4SԺ�6�u�0�����
�z0�t�=4mǕ����=���B�5���o'�W���N�ϛJ�m�\z���l�����v��!v��(q=��@]�gUX��W�XŸ��x� �@���}�w�F:қ����ɶ-��%�V/AB��{J�8�ؤ:���%7��,-@[id��9�<8�G>��h�W��;\�o!w���W��	�j�^�%����x��Oj��q�������c��
���2�&q����!t����Ř����@�#v���ѷ���oh�����2��t�mq�����=u���V�.��4��4�˼��OFޑ��v=z�zFp'�v��ZWV}׬*��?Ql�<��+ou:á<�[��X��G�b�U��+IlV��/=���N���ܾ�םl�w�>}ػ�`6�
H���w��.�����|Y¯�ds]\:����ֽ����*�^��Y`rgo��l[�����T
(��v�SE4iQ%�:U׭��Xk��O��k9s˺<��e�
�uo���$w	w�e���˩�s5��=��`Ӷ��uun�
.���.�ӫ��,zVr��9:z77��
�1B��@W'n�����o�+�oTɺ����Z�}��ˢ�E��[�D^�������n�ാ�Q���'s����p��W}D������,�c��߻�-����l��h��n�[��m���챽�)*A����m�����n�U��+s�oR�EY}��wh�W��4��B�a�kv���C��I^���Zw��*"1˾���f�޽�;�?e�27���FPH�99�+�ok}wͷ�wo7س!�:�uwNFw8y��o��g�:��"g8vw>Fs�y�����wr�оg[:�����<'3��鸧9�b�,��H�a1(�l�Im(�.�v��]�Z���Ñ�N�c���[f2��9�F$�'��=��9:�2Ȗ�ho�������y��R;G�؂d��	%�Q��'��7{��m���Ib�w��(�SiZ����n��'�S{�������\_`YCG�;�&	̬=��q>�2�������W	/�<"���-(��{��g�ur=�-��L$���J�_A��{�<A+�szl���C�l�k���3�=̾d�Kp�d`�x�!P�۽���˖���jKV�.��p�����m�iF�Q�n��g��Ot}�uw"w��,����w]����)����$F�}���۱��]\����vwsdn9��AE��A8v�-�Fq�����x�|3���{��I�I*MaIo@õΦ*㷽�R��b��@��Sq'�:X����QK c�yM]V�.�3:d��<ɉ��{����u�`ec��ݔ3|�</Nq��w~�Ӵ�o��f'�Nw�[ed=����I\���̱W\%<����s�Π�Z�J�]�k����yՈ�ݰon��蹎�n��KE�D�n6Cxm�V&�ͥyzp͙LI��SU�[�K�փ;u��࣭V�]�[ۨ�C����E��i�JN;}�7D�����k��JH��X��3v���d�����n�X�Sظ\��̭ܬ��M��q�+�Ղq�Q�
Z�i��z�
��Ir�f�t*�6U�CF�R��U�)Î����j�k�f�ƭdD2f[���[.��fJ�����y��U��	W-AnوG$�w�ˠ�OGpz$��,š�[Χ�/Ge�h�oo'ju�㛸;zW�B.����Q���
�ں�����8���j��\tA��Ɯ���о<ZfH@�-+��j(M�J�%J%C�,CɃ��\����#G4 JX�G'ψ�غ�)��:���O^[�%Ť|{{%_�h�/�c���V �G�e��ׇ3���H�+�"���1G��M�[��u�l�3/&�J6�G�D�| ��0�$�^A�ɑ�������JRh��ws�f�j)P���޻���%��� �w��l�\#���<{r����ak�M{3D��r&��sY��1���wG0\%Q叆����SU�$���0��w�kZ��G$SB�lBy�:eE���c�C�q�)`X;]�-��.�7R�$���=�Pf�ݦz�ILG�ޱ���V�y�ӧ�mo+@�=:ݲȓȓ�(ݘ����6��u1h�t�k���H�#�I�����y/x��E6܍���'I޻�]�.:�5.�MWk�����nۛw%�;0��(�+���^p�ok��v뜌��]{��jUp�2��,��}��'��ZmD�&;������ތ=��|G� ��Γ��m�n��GS1Jz�w12��8I�=��Id�׻���jv�=��b������H��M�u~=�����vs��&'�t�d��̛����n_e��/RY/���
�+���M��]�[!�rm�}t�[+3K���U9���;��e���e���R�A�i�����KbW���
�c�����*��[���g���.���8�L�0�m!W�<�d��g�A���t��UÒR�������݊n�t����Z�/6�$�7�������I��U���'*�;�;��$�7��g1�cm��zҚ����V�ui�wQ�(�H�H����82��,&igb��ث�0%��fwP����Gq�B�<{�tz�V���U�ƭp�r�����xݨEp<�Hݝ�˷"o1�=�6�x�ܽ�4���#N���M8ہ�/���i��GՒ�nM��	 ��ae̻���-�د�ݶq�傸f�I)�A�^ǆ,�L�%�=�sd��탙ۧ
x�7)!�M����'�a�N�<����.��d�k&����θ�/�����8u]��veX(� R��U��3�YK<�]]�a�f�]`ӯ��ۺ"紱']�p��kk,��\k��x��mཽk������4#߲b�[�
���w�����(���#��u�T'�_[�����E;�g����*��A��3 ��b��.� ��qe- n>�n��C��a��q�ٵ{�_!P)$�R��	��MD����뼲��-־3���^B�Xt���ҹ���균'2��aCe����^b'/iOO���ޮ�մ��*���Ifd칵z�fkZJ�%�\t+M�Œ�W#8��۝��9(!Cgd��NQo`��y���k8���!m�������*��
Ny�m�܃��{h��ݬ��hn��N\4v5�hN��F�0S���l^#Y��L���w����IR���9�`j�t��mul!]$��fq�\:����wItu����Q��&��xre��=&�bD�d�8�wu�iQ��G��I��K���ё�|�Ư�9��pr�o)�B1lf��bW\$* 7kC�ʫ�!����T'��#��ln{)w�	ӕ�̥��N����(����7�ٷιJP�|�`
��u���|�Â�u4tf���Յ 2��:���#{V�fjx��&)�:Ԭ\j��i����}j3��28��jԚ¬�h<ͦ:�vl�<�ݻ=�8��d+S�V��5�5�$V9I��oc��2n��+��#"ymA�Q�}{g	f����s�*���72��,��S&*�eJ��L���6n���Nu�-A-���ܻ��90뭚b�Εu��K&%;���T��2&�O��!��R����v�&�{0<�byIӓ��ÏU�A~v�Y��Y�&�=���n�Բ!v7��((�x���}[|�v�=P�k\M��w��\P�dP�e�v4e�w��.kWjd"#���*i[�i�2u+���d�Y�AN�������x��Z�۬HR����?��ʮ�W���Zj��ѷ��Qu[�d���"�M�7���pi�8����8v����\���M�m���\8[�"���vV}֍�Hޒd��Yd�;;\@�8�+[�]YF޻cb)�Y��B�կf�0(-V䳩_"`&:�8��u�*uvr��H=Ԝ˾���(]h�t�Pp�YW۩�sM��kˁ�&��U|����<�[J�eu�b�@%Mt��(��AP�Y��Ȇ�M�[��f����J-�X��b�,[�1��-�㬭6�QI�*�u}}���A�A=[���]ŭ��[F.Yj�5�W);]v�k6`�C�Fp��ieh���ed��#a<!��������b܏l��o[��s\ui�k��(Ihs6���'gQ�S���9��u��t����_^1js9���Z
	T�)��]���L+�����f�zye&f�Z� �l(T�e��jw;�єP��8ԏ�Lm��7]8V!\�ޗ�m�M�s��ᮡy@0�UB�U�f�����u�޼oQ��7���}����½�5jd��=�;:�?]=+�s�J<�v�q[kqyM��<Et���t}�,	}N�1O�����l�ܬ6�=�b�1L�
����3�u�i8�]�Z��O}��e�~��ږ�,G�9k]U�7K����W���x�#�T���H�9 o5G�qÒ���p՞|��l�
=��-�_ܩ�6!�%d�m�Vj˗�nJz�j�\p�-9���S��I�M�T����9R�Ä#� �����U!�i��<�Y�F8��oq+W���vֱ�a����Тbȓ��zt.�x�
vj� ��n���}�䰜}5Խ�A���(nQ��+��!76)��P3F�n�H����m0/V��6�#ƧI�����M�%Mū��X�����{�d��y®���2��;9�����/�ӵ�ݻ)�Χqy���ǥ�����#LVpN�4	�[�80ڇ34qb����Q�;��lW�ᶖ	t��b�Έ@�֔s�\��C_!����	��J�l��{o�Vw���db �w�i6[���]u�Bq�a���r=A%��U�sp�TEiw�%��Z�ƻ��{ݜ�{�7e�;�"�v�}Ԧ����3y�2©`��R��R{w�,���JK���{v�r���=�4��E2�U;0�f=lTLjܾ�۔V�O��a� ��<��=޽��]3���-�_!֥�he���������[�0Ɩ�`�G�c�x3j�rT�A�k.�.�}�s �0��趇m��O�@��ŝ:ue����wk5]��rk�	���许���Rk���> hm�/�9�c6u�M��89;��:������z�cq�#�6�x9��Q�xV��g	5�	EB��B�H�e�%*�s�WKb��o�B8��j�d��\O^�%,<�\{��HP�z�fP�ݧ*��sMN�]n]�]�w�qM��Xy ��`U��km؅P�;V��.�]��vCkܗ�f���mZ�w͵�+ n�*�F^�t��+=1>�3z�f��g;���(��c ��[���1�J�U����=v�n��N]�c��Ch�l"�5�VfvJ9,�]ʸ�v.���
W����h7.�ԖEa���[hf,0A�g�0��Mz�4�.���ʙv�eLu�Ɓ�a�NwMZ+��0W,����r��ZO�m���ۋw�.��g1P����]v&=���.v�eul`�=ɲԮ�ܞ�!5�#k�+3p�/�s��V�U�u��:]"�-LԨ�n�ٰ�	�h��8�zk7�)� 7̊oMӌ^���Put2�뾻,��wr{�nG�M<`лٺ�#���c ۉ�g �ej��z�`��ΥXp �L��t��'-"^���i,U�3u�̸K����A�q�e�f� �H��Ɲ�Z��۬��2�㸊[]x�̈�|�Lr���Q;���Pes]g]�T�⮆�a�{���3��ǒ�6����q��Y��80��4.�-\�f卭Wf�%���&[��.T��ײ�-��`	+�]�Tf�f�L�F�]�ӹ]�T����ħԐm�����Z��ݼ�@l�t���w.��b��"�ka�4n�s7��w;oI�$g�X<p�;|�6t���ܞޥ����Ɲ}:�T���3��_+evM���ZUÈ7�x;gX��$��yk�n7x���m���M�:�gu :�V%@머�+Ӡejg�*ʳX�Q�G/�	�
�y{�uohJU���-�E�я�V�M�y�%:���F�����-��_%�"����Z�Vk��z�6}vW3Od�Yy��E�����/�pYbt��>�2�nժ��}͔�d9Y�fB�/,��u)��.E�������}5V��e=�kf"�mJ,����{y�x0e�'��,� k�Ӷ�@�N;t(2��<<(1�Z��T��-���<��́�v�]�7��-�+:�tShv��u��ƭ��mPÙ�N��$��EYz4_��k{U+i�v��T�K��N�ǉ��ہ�ցe@���Ixy�Geܙu�HxN�!��S�N�}N�Sj��@��<����V�	��d���hiHK�=��u܃�@GwN]G����>��W��J�݌�kB��4�d�_C'��u��Ww�e�=�
�T㩗Wev����q	n��L3��dd#�;Gzik�����j�$�9\L⫺Z���"�,P�p�z�5 �fsYܕ͒���#Un�����*t+Su��eñ
�vQ�2Ň�B�ܯ�]b{�l(;vٌ����*.�xc��٭WU۷*�}%��J����(���j��vĽ���Y�2��X���J���K�v�D��ڝn]��}5���yeF�����l
�*�[�͝���w]�#��	8�+%
��C���x��۳��[�qa
nd��T�S�^s��D{�����Y�C��FC����1y4������M�H�;m*�]�F&i����kQp�g#\�&jJsN]�a鰎̫j���hi�3���Ɩ���@���A;.�邞M�)oB-ð�I0�����n�K���clrA�뷨F��+;=��]���6r��t���-mX�vgikvfjb<���&z�ܽ���qE�[Y��#���wu�-�@�$��c�q���qּgx�/��6��;��o4l�\J�V�g�����T�'O���T����%�=yr���vD���Yy���a�:�k�U���X=��f�;��ꇘ�Y��.;z_�NĎ5���$ǹ���(�y1�eɯd��sԺ^;���e5�Gsd'��K[b��\;�X9g�'�Th�@�W��D����6�\L^#�_KkWsdo�2�oK��{E�*����H�km�Y �.K��{1��d��2�A_�_�u�q�����T/���'&W^V��}�/���E78�ӽ���©�Gg��*��aJ��G���r�R˭��У�@�$x8߰�ݒ���)��ufu�
�S-a�,��K��hR��ॾ��,�{d-f5DG���N���}W������vxW]����[fѲ+t�pt����!�_v!�����o`ނ�:�4e�92���}&�B[j�:8�,�)T���CY��:	i��;�Z;i!�6q`����Ի]�sQV�.Ei�t���7���Wwj�,wa2��(qD5��v����E+��u�2�s�)����'βnV����y͹J�@�a\�W���n��aN���0��*��;�#\��R����,Y�1��u�Ë"�L�� Kr`Mܕ�������ue�5y�>L�pn�����\6���qWj9N�³�nRJ��ڱ՛o��r��-z������ay�:}6T턛5+u)rwF���]B�y��<�JW���b6at��/�5ڍD�����ly�w�Ё� �	$�|��#�����0�;�{���n�����Ec�X���d��F��8I�u�i���5�9-�'��[�����r@q�=���՛#l�R�k��/�+�-��q�m�Ju���ۼJ�ܖ������!��\���;\9�m�go���)��c��L���hx�B�V�q�xb��㫙8�zHđ�-��s묳���or����w8�u'6�PV4��Mٙ���J]���L�n�i���6��cNp�-7��V� Z�44(,Z����)RX����q�d�黷s��Ҷ�**�e^`r�bYؗ����d"��5�}X�!���q����l�����c��t�Ξ�٨,ۍ�h�{5K�bk����a9֨e���FݤPk�T�������l�u�-Յe�d����}�$��d�
�l;�zȵ���Vn�KP}�W.�;9I�#��tC\x#�r����QRL��L%���̷��X�%���g5�U�P�KՅf�+�a������09n T����t9��xn��>�.�ZڟbS{�si\H�T.�<�.Q�>�O�*p�#��9Y$6>�9b�kLM
�n���еف���=�J�h�)�FM{J�<�ï���6X˻��+�J�����f�o��<<Pm�겺�#���9 %�hU��,��W��+M9��8,�k\U���w�:�x- -�;y��cՇ�B��->���'��������}Gw~*�tN�8��� ��9�ե�+ˁ.@��.��=����|$���*��Y��tVl��x�GS�tc��[����$�C�C��p��k�!_a�-u�v9���u���(
�`T�hs�F�%ʻ����Sn�{ޫp�#j��Io��Js��e�1hR*����01PPX��Kɵ,_�,n�&f�+FB�]���e�V�5��_.��р@L�+�wz��%�� 45(o_?�Z�^q�;�[[.�WRt��׫�CYzjsdG��V��E3���Ρu-�)NS���\�9l(	� ���H�h�;xeب;�hY'ӎ*d3.rx{�Q���70/UW�X�k W#L�FN��01�P�zJ�J�����"�㬼ʹ�=t�D�P��W�ڮ���n�g��|܂�Q�6�$����p��E�U|}�~������﮳��FADH�1�L�*,"�,��2�6����"�3)������������l�K�ޔ8���o��j^�{�	���mZ�Dh-��"�#:��{V �Lx���Upu�ii�6q�� �8�'V��A�B��ggP
�8ܢNu���j�9��q��᛫�J��tx`�δZ�79�[B�<L=���U��Ș�������h���z��^��;��}��u�nU��h_-p��>�FZ��*a�^r�SFު"�C�U�J��h��~Z��feLn{e�7�7�sE�G6@ޭ���m��x �r������Rne�/��]��<�􆇻^Z,��,}��ȸ��������j�'>PL�F�3��Ku����d$9�
|Bİ�Z��m36�AGH��+%g] {B퍁���k���G����z���I��������whwdLE��wS��B�-G��v\��e��O1A4�U^ZH�������ȞS$���;��a���=�0�����`�0VHi�*A���$Y*Q"�+
�Y��I���].f
�Ø�po6r��f���۩�)��F�R(�
T ��(!�=�q���;
j�-�l����{�6�:���Qθ��o���RIg�kD@�:��p]Q\[2�7�B�z^K��@�|���U�:a�H�d�Z.��s�D�dnmoev�um��Yy�E�q�+�>0V�i���������=v�7��7a�%D���U	��`��	����}�8>܋��;؝�#j��t� �:���x1�7��^h�Ԉ�}U�z�w�=g�����wS�}*(+[��kqh�8�4&�Dn���i.���!����o ���oE	M�n]�ҷ��=_U|X�3�`�*C�P��Zz=�{7et@m8p9��m3��U0��rV�Q=MD_]gC�C{�+��D�z1U�X_�#��0�-�~�Lݚ�x�uǗ�4sv���������Ff�ǃ��*(0!\%Y��>���rs�G���nP�)*���wc3v��D��bd�x˽��D�d�nW�WcMs���΅.ndx�`�*��D��y<Ӗk@#�z���W��{��0
�|�ͺQ�ԣ����D���2���Gb���8
׸+���{}��>7����$$��@$��L��y	���஼]	4�uZ a��tkp�O:�ij�O5�Z@�;��I��2���/���0�.��]׽^�_j��Q}�ّ�,S�x���D��t��+��&��M̕he�\;��ۚtR#9��}UU^f5�Q!��G���~�Q�����RҦ��e�Zwb��Q�b�c��	���'��oiw\�$�iBt)~�B�$��B�n�����}��,SÚl+5��i�v]�xs���UR%��\��f׮�(��N�*j�[�}���u����$�a �@=��ȘH�������o��b֘��	_^<��ܤ3,�KJ,�,�L���Xu�5$|�f�KІ�;�sf�p�nܶ��H�5�����9��L
��VI*�{	� [���V'�'����X�$�89� B��3<��)\Р\{�������9��������Hl�� ���)�G���X2�V��"�^���Ї�O�ul����}�}���}�����2!2���I4]��V�z���i5v�$�~�:R���Du�2�Ru��:g���n3	��]A4Z=��ʹ�|��DQ�B��P��@N��d�!���$K����媛�C��%Bjnn� ���lS�9�`Ԝ�&�7� ����Uz�����E�,���Z��:��v��]� U��z� �N��B��x�:,� �c�N.y5U��=��L�q�"=�Dz��p�b�Hm�Pq���VP��NdCm�lp2b��ߛ�V�LD�B��d̻Vҙ<��p�Q��ٳ���ˏD{���Fq�-de�"��S"����Q(�JE*�,���Ȉ�+ eDm������rT=K������ͮlUiy#�V,VK�@�y_%��N[�e;ѧ��瓋�� �E5:�����s�q��=iڥ�iu쎥6��&>����uӴ�Ռ�skd���(	Z�ޜ�nG��#�<�jdEb�@��P
�U��F3�DhWh���B�	���U���Tc�)bU���Y�w��#�_1B��L`m/��Tѥ}��x���=�l�W�U}U�UM26fB�V���A3�B��Cs�����<�2w-A�7��	��Թ�w��يx&���lǒ��'"�.=����肽�c��..�ΐ����\ܖb����u��iVt꾣[���`�Pp�m���+ޠ�0�P�������Z�"G�[�^wk\�l�CD�M�KLj�<�]�VVdi���a�r�8�ʵt���y-�GS��r��~���^���f���s/0���="��J Cp��%؜i�U��l�a����s^��R8'�`	U���u@�=*=o<-u������D�3"�K;���c�Yt(=�.n� �o8C(+�ڪ�ܘ�0Z��\V��.�tC.s�I4:�U�N���Q��7��=�Eǽ�ů&[�(��ƈ�bƽJ{sf���h���!��MTF���|��wv� 1�ª�՜�1>,��κ���z���=�a��봚�P[7�Wr��
�A�G����B q��y.���j����ә�[�f>���ס���� y�A\�΋���0� 3I�48TʀS����z�����i̷�/��R�f;� V�[�)3�bՊ�{ި���G�苨��f���yO�A5�[�f³L�V'D�yj�B����*��ge�
,�
����U80A�i�ޏG�}�8�wJnT��ԥҡ{��-fU�H���c�]��) �������<�]�j}w��Ӱ.e5+dc���so>��U�QϾ5Kf�{ʧ!��?gA��4��f���FIR`�E����� 
�/�jF�fv�-�+%Վ�y�6��U֝�]�m������؋�Gr�p.��;[nTٹEa�N�X1�V��{ʛK�2�[�V᷵b�顩t��.;��Ţ	�xXV.�D{e*�T�h#_�#ނ����J��b<7��@��B�;�a�ҷ}O�}��֛����tv���S��o�p���{��{����L��n)ӎ���ЬwŖ1Ww%M]M�G7��;.]+� }�)u�inP���GL'�z#�"�[ꘪ+�����D�ɉ�=v����t�f_S�0JB
a���ro��!�v��UEL\̭�jv��ޏG�) ,F� @�� 3�K���ԭ.!�:	u�=H0
�Y�&��	��]�B��/W��������e�U�W�:{��N��/�df�z�ep���#ڕ3:�U��&�o��	ܘ@C�̜���ܕ��}UUUR��S[���$��LIU+!YX9�L�ﳗӞ��W�[:Dͥ��N^e9�oL����qU����+�Â�����</+�G�g�L�Ȗ�EPV���M�ݻ��N�¦r���C�5]��k��v���rkbLd/�Iż51]q ��ؚB7O��{֖pzP̃Q�v�-T�ܬId���L|�$1G��5�	��@�}u� �*r;�@w:��������$�9�~ް���w|��x��m".Q�0A�K�(UCh!ܫΉ�9q=�/�XB�^+�E�[�`��
+�
+�í�����"=n��9�솼�LV	3���Y�d�O���}��Ci�i�L���'nO$ڿ,+B��4׫t�e�����{���:0!�i�����t��S�vc�Ʋ���5�9�9�݋;H��:F�6(4���+\M%��`{����/ �^�UQ�߼;\�Ӓ��b��L3IV��+��sM��,`� �R P4z"
��R�����>���Zʞ���%5�_(���Ncm2pՌ����^��p��h��-�O�]6��%��]�zv�co@[�:���J�5t㹢����zc�B��ު���U(��:9�A�^����m^L�P���4.��@�<�h�Uj�8~�ΟJ�7�g2Β�_[�n�ٰ6gDA��DE��r��v�1��Z$`���H�z���#;Dq݌����}���N�n�EfX�E;PW:Q�"��w���ab��dȾ�q�x���� gv�g��^��i���3/��qeS���F�t+L����=����в=��ޏDV	�.If�!�ʄm������z�foIv(�F�Q�Z��y�뫙jjr���*,����8�'p��Lg�^�W�����Q&s�Kי��}߻�vs�W|��bE����c�}�]7�퉅��1�R�Ù �ܮo+�7N
6��Օ�{�腵����fFK��7���!�z��.�l��َ�SB���R�y:s�:��MʖF�b�f
E�t{��wt(mNv{����A��WG��T�P.�$�E5�^r���Os�b�{���������uY��(P��� (9��6��)�]Ab�c�v�F�7���U���9�<�/�۽)�:�<�#�֬Nx�N�8k��wA��TS�f�̘��2�\8��2��U�#����#U
�Ɗ�g9�q�,�fXH�q�s���٢a�G2�%6����v���b���M��]���W��5n7�\��s٤ЈT�j����}�k5ۏ���&}�ѷ-y�LM��f�
�2���.4�;r��#�3k{H"����tHÆV��Z�}�f�b�Nׅ���ra��zst���\���Q��u�ĭ�Ѣ�s��ie��`�YV>��F�s���5�h������"����j����Q����кJT�Do��DE����yE_�:,��2�\�׮�{��5�n�O}t!�I*>����(���.ur�CA�O������r�I7n�����U!�Mh����.hq�0R1S.��I��j�q_	�P�BR��mF7T���}�vg�����kf�.�����^+���UcN�t�ﾃV�؀�A SP�l�~�6��W�[�n[����Y�;\�W
�ޚ7�\n�C����ezh�	 �մ�U�>YѾ29A�����R�!�[\#�O\U?oKUV�f�$��#^}�	w��#�4�z��iͷ0�⻓��$LQ����`��=׈������.v��C_5\�at�J��1�r�Ҿ-O\�F,v��[m�c=�����̀��NP�!�py��Q�!Ye�*)WX�32�&fM����2Ξ��doG�c9�4n֛�MdIR���NG�_��W(��g��6iv�M�v8�麝.D���>�{���%>v�o:�i�V>�S���t�EqK��k��w��V�2��k�[�\Ⳑ⿸w���Q��1��*�Aɱi��]��(��!�9�����B$��wL�U�t��e����V�Yg� w��e��8����8�vXY�By�dx����;7�����:���ػA��u�a����/f���rQ��m�R'�j��T���L�q���b�+�0w�[��\���5�T���W6W`1�r��=�
��'N���ubX��
���F��2h��]�ke@�#�5o�����Kz,v�y��,�vu��qSA�e'dg]<�<������w.�ݽ����d��D�����vss�Q�nŭ)�|$׈�C5=',,�4M0�Z�30��j��1�o��5Â$]�2�v�ׯ*.�'W��\�Ƅ����'c	#It���s�1Q�`�F�ubU�G�o��'5�r@&��q�Л�!�υ��7�G�S�a�} �8��)k�AU�z�\!�"��b�4(;�C39�M<ƣ��[�.:��9���P4;���k�3n���E�*坎3��H��x�8]��4��Ң�.B����z]��y6�����~I̲}���
�O��!�m1a^0�,��QC����T?�W~��]X?7T�I���B��" �c�zc���<^]v>́������߾�g�x� ��i�BC���
���0O��Z��?�m�aXm
�'���~ͰY��W�E+��P�SLӌD��e)qʐ$z��<G����M!��.���4��Ͽ��I����H�~�@S�Xc�*'濓��C�I���N��
�n'c���!��=������wן��H@I�X��T?&&0�y�~q�Mz�	��5��P�ĕ&�Y��%��k!P���q�16���逳�YS�W�V,������{�_�w�3Hbbf3��Ϭ��<���6���c���L�+Ҙ�0�1��>f�[�5���6��3�X|���*x�b*�2��A��@TX�@RE�+ Ā�Ȳ,�)*$b 
 �"#��M��X!_��°�g��W;�ڞ�q��8{�{�#bLE��$D
~Vm�4�C�;hcPP���'r逿�P��??0�1�����0~i��ę��6èV���X��"*�OkO�=�8C���#�>f0P�S﬛M0-�!�c�
�~��0�����bV
|�Đ���������'��;A����i6����z���/>׋ｙ���c��{���0.��:����U���+�
�`��_2T���LLx��\CL*Oϙ���i*ˏ�|»a�������~����|Þ���s+ |�3>��2i��|I��*c+�	 %d����y%C�4��=@���ͦ V���Şf bW�&$̾a�cm2��d�Jжr~��M+=cމ��BB�k�L���]��a�6Ȣ�~�C4ϙ�}�G4��S�?&!�Az�	Y�����;�ԕo�&2cVHw��ത���d���H�-�g߷�o�����P�,��$�2� �71�YZ·�F,ՠ�n�S�]����d(���:���J�iY�di�WȐ�)Op��.R{��g}���'�����k!SI5�Y��I��a��������c<��n�o��0�3�o!�.�6� �é��y>C�)P�,����>���}��@��J͠C�La��:�� ���d�N�Hq9�!��Nk�4��~	r��y��{[w�������i�d�T:³T�O�ڳ��b|�YP��;���!Ry+�
�'X���`)��Ci�����e�O�y>�Hm����;�~����;��!���wZ�i^��1'ߩ4����:�!P;o�}���?$���;I�P��={��
�$Xv���+䨣�~a�H}�a�l�e����=������O�Vu�yh�&�}����jk2i��T߮$�+<����L?�+��~���2��+���t������Ry1/���i��r]���럷��]~>E��]��i�?̛Aj����PR��aR@�&�|�Èi
�2Wڠc?[�i�v�u�f;@�1&���u3���������߀�Ɍ:���8��M:LIP3�a�}q��1�
ԟ�t����f�T���!�?$�?��~IuO�Ri���1������vBM����ۻ��|i<�ix�0�+4o�_�H��Oɴ��d���A�]!�~Ld�k��m��1�f3��c4����J�l�}�Z�?2G� �f<��b=�aM�ˮ��/!zi�?&��̘��U�z��yY����a��3���/�N&8�[����lϩ�4Ͱ�3�?:AAO�0��� Q	w~��s]��?��! Χ|�fz��I�i�g��
��u��+H����'�"0G�&��" R�Gvj(T��C0(i�
���d,�X�%kBXZP5a��4T.vt8�bB �Do]LC.������޵�v��	��g���l�P-DT���gg{�y|Mdk
�i�ueb�����G+���k��>~M+��@ڐ�f���~N��/�ASױ^R9J�X�-L�؀�0A�Or�����}kf��%)2�e�B��Z4gQEꪪ��U{�z��C�,1 F{���B�(�jfB���[\<v)�~1-I�]�V+���dN�����/��݇�f(6�Y��}U_W��ǅK4��o�<�Y���fڻ�6�۶��>�s��rp�c�*>̡j�3�(�(r7�T|�@ڐfA1VTz!�G�#L+lUns� �Ϭ4��ļ��rU�"c���<���z���M�Ch�I�CЪ�����m���{ު�u/e�� 1t��������qp���!��m�8�PT�ѱM#�v�]w0r�]�����TB�x�1���z<H�:�Ц�����rq��LVI�X$Td12���B� 
�!� ��G��b�����R�l�dSV�J�r�ݞ���Hj��P��/�֌���ǹ9�7z�ʺ{���hќ�����󽻼j3mWejD��k���ud��|��eH�NK����Y���n�v?W��I����Nc��L陆̹�H1�H�'f�̫����Ww&l
�
��j��N�q!�]`���VjND$�*%@HGN�D�8��芶�a�����e�ך�Ar�Q^n�w)t� 1n��\�+��3gQ@Y�1]�\\D{�^�or��S7O�$q�f�t�B[j�*�0T�u!��Z��	N$�V�������4 r���:�w&v����@䄁��S�cޏd���.��p���w���������PD�����b���5�{_J1\Ԥ�nѢAC.G��A]k �O�U���T֑�*�C:p}QN*��<�SNp}S���m�YK[��k�x���Y�P��-�o�����@X#r����}���}79�{�놬u�j9MA>��).��嗢 ╔Ѷ�*W��D�6�mgQ����K����~����u���zP��Z�'J:rW�����谄$�D�s01}�.�By��VqmѨ�_n<ۣ*Ovr�0����1�γ���Z.>v��=�I��b$s��W����`����7fz�If��j�������d��g�}s�
H��ua���y<8S�/�ٗ�_�B~���{�Uԏ{�e6��؂�l:8;J��(�VQ�A�Z  _t���wj�u���ث�`Z��+��g
�*��u�#�����x����vj1��K`	dE
�6�ӡdL_@�S�}�����֎gA�ڞb\��J<���g�k�G3��D{�"E�N�,�Ad{Y4�\��4dĮ�`b�c� 1Q�����f	"�-p������{��w}���~�k��YF*��DX�UD`
�(��H�澳��S���lE��U�<γ�o��]�(uġ��"

�c$��cƑ� �PQ`�,��P̦BT��
/�4�g�H���k�c*	�>��Dn��2�e]���j���Ά\Y�*�6���bojoc�[�Ww.��9��*��A��S[��f�2u9�� �2P	Gp@ár��c����D{��{�
��4^�C�p��]7������`����0[�	�cz�-���<�//�B�E��PA����+(Bd���2_��<�q1���{����
Qkw�<W��zlA/4r�y.�,���� �Wt��㶸�ۺl��p�PiJk��z�O���ޣ��v�6b��uB��E��B�±����2�h!c���kq�LX�ȷb��w����m#�8�cΙ;�Bqt{�_��Gf�/��Cӧ2�d�V	d��;�8cTS1���u<`�1[�����3�iYB
�p�������q{�ވ�W��,p�z�p-d�S�#EM�}s�9��o4`ꕗ{B�\a��T��!�����"0�XmW���w�a�ٷy�"��m��
D  �B=<6��������c�+�����f�i��Ua+G��iIu�x,�gs�-[)�c��M�ֻ�c�9v4m���]�� ��U�_73)3f'�\�(�<j
&�����Pp��u�Ӱ.���SmQI�hZ&k�1�[��DLXB
2�gY����<^���2��`�8 a���T���@q�P\�j���T_U}Tw���s�^��Z����W������?I	n�"�	# � <� r�ɮ�I(K�r��z(��J(�}.k�h_k=!L}��N޾��3P�,�U}T�μ<�n�X�7��b�{��ghœ}}�	�q�4�jH!q��ZX�B���M�e����bY���U���UM����zG�@�TJ��8�_����U����6/�H{_�u�鱆U�FC�;U�8PR<eYb�1��Qݧ��1�
{u�G��Wo5��+���6%qp��q�m,
b�%�F��9��]�t$"�)u�V(�ky�[.�Z�O����ӟ5[�C9�ݕb�G�9�(D�Bk��c9:�-�w|�㰙��E4ǵ}�Dt�(�r\*�c
���� �/0�����{���25���`i�mA�b3��6`�ݙc����v�إ�+Bm��BP�u1�o[=��k-��3����?�@ f{�>[�Pz�i��#M4��vqrI���i_R��%D"�#��;a�R��`�L>�y�ѷ|k�g=� ��z�����:3j}u�6P�1�L-�L�
L���:d��&0/"�;)%�;f�
<JG��7^������U9�5����k6�E�})g���|`�$-�������$�k�O��6�k&�YPE)1R+
�W����}+ABĳº�2r9L���85�%
,��N���Z�h��w|$�ez��b�ˏ�|�*|�O�$X`"����� Y�8 O9ބT���LvW4� #� �"�
�@R�
^�Rԍ�O"]�҆u�B���+n�jf�b����Ɯ\9��;Sr2p}�v.�뛚��ݥ�JI���Z��tvN��Ȑ���MC�HШ2
9X�����z���Ml���ͫѤ��������@�3!��&C`�U����l=�a�0m^�2*_�u�2�${�"���Å�^���?����JW�T^Sc�r�<kl�0v���z�k��>L�+ɭ�.���'����ׇ;�D�z-Lfj�@�-�*N�<��.�D{US�z<�L�ّ�Kh���)���,5�mVQŀ��,}�ǽ`fb���%.Յn���k�m��B��4@ݸ�.~�z�����oD
��E9�{�ӜF��]�.l��)���(T;��~>���Ht��Q����$�åUW=g1�����Ӽ`*y?G���hhc�iVr�lx< |��6V�����(�%³���ox=�W9DR��H%��ռ��c��/�a�β%R�)`�)r#�(�B�FB�*E�`eR�lċlVS,�2��R���"BL�Q��
b
����ҵR�F�2Z$̥-����Ff`(Nwi�~5�;����^I!�攧!1"E�R�*à�K1e�F��u�sf8�l���f�����yܛ2Y����c{˃��:��j�h�~��B���{�WRw��ۢ��_@�+<+�Hw*�&�Wm�^��rҥ(���a*��.k�B����b��DD2�wL����o�P��E�ᄞr�q��b�\���yx7�Y�R�I�"�]�@�Ř���o����v �0�͹Cٵ�PJU���Z����t:�mh��X�n��!�^��v�,>C�FM���D�XD{D{�=\��`Ⱦ�č�.�&��V��؆Q���9�I[�k��%���^(��+�
)Q�_��B=���F$�%5��f($�27r�ꡄ�%1����ij�v�.��Վq��X�����k�|�Ϸ��օ7#�Lov�HD��wW����J�ԄV�V/]n�H^��[��6��WZ|�ʥK+z���*a}F����wC�1:���]J�n��4S=V��Hv+�Ȇ��L�{�/2�Ҕo���h�S0������[��SZ���P����¹뼵F��v��ʠ ��Zjf�L(9]����ww�m;�v&R�V�<lR�~v�D�V���{{���sL�o*m]�Z���,X.�7Yql���GsP�w{�٭��§����r�h�>#��<*�7������խ�BK��B��I�����ƒH�釞e��aW9�J����f��=������>����&�AQ	"2{y�Ք��Ȣ1B\��{�Y͛(s�H�ls��i �y��֛�%a�`9@~n�c�7�����]�Z8��kY��'���7�$�T��6���Qd$b.wF�}�k��ʼu�v ���f�߻���*��fwz�Lrڥ��F�綬�$�>��@X��g4S��ɭkE���Wr��f5�e���*����o��T��T-�tGiW�n��;
s��kk3HU����c~��tРE�+��Ӎ8�z��=�Y͗��k}��w]��Ϸ�=z�`����;ٳ�`�®����H���4Gb�M���0ؔUڗq�s;Fd
U�d|��=�����9u'��G�k6�Z/T�B��a��Jz �q�zW��v�ROkTN���ͼ{����]K7������D�P��\Bt�Q˛H--��7�-�Ųk��l���.�2��8����{Gok�Kg���¹��`�t��R���X݌���7O̼�T�9zi�	�Um���Y��n�5�Krc��$:��&���5]'.휗3�	o��7�3�����\qT��>L���v�l�h�}O.��)���S�s���:t7��8��:�ܢ�1s)�h"�#��gbyEo�>s��Ovj���T��r��Qi���=��G�(8#��-�����O�AR���nƞ[�ge��`�`�Õ��m�P�h'R$⁘q��r���l[�V�ox����{�׽��D��^ʙ6�PO���@w������:�V>�rU�x��PێN4+n��TA3(v>r�I��+�Z�ws]�mV���u��ذ��;�h-���qv�e+ah�c�5}��a�� %�H�� ��l�Ki�ݳR�H����)
̢�&�ǰ����������N	�y�#�>v[��+�p��8f�Z-���i��:[�D3�&a-��O��s�zC�����i���`/^�bz�Ǣ�.H�%� ���%+7�4��Ɩ|&�xX�b�U����6�P�4���څ�ucpU��l=y�>}0��K)��H�^���:	+�tj�A-�Udht(5��Õd�}�&̨y��o,$�:�.o���aaݻ0�塪Kݽ,�jl�m�����x�}y�\Ld:�n��j���ǭя���=!��������}q�Ĉ���~���r��6��T��՘�9�Q������Ù�U^��s���d���p����[���v���f����joKT�ǏǞ�B�aTkm���#�)��qZ5n(�0������#є�
sq���ъk�F�;���C��+{Y�+�e�!{�B���{�5ֽ>��&�M��W��|k�:�v��L&4V��kk�Vj��z�c���|��R����vT{���|�ާ_	(��z��s�h�o�2_d��#��*G��jt�YX���Pv�hM�q����	^&���bI��CX�����E�R� �UAb����T������%�(�E���f:0�`���-�1W[eY"����E�֫��hn�f���	n晚p+��Zݼ�4�5�� .oaB�6��Ȥv�EՆ3��C^� ��4Y�d�O�s��eJ�MU�ꋪwX��4s���o\2�i�]h&�\����,��g5�v��z����5�e�]�W$�/�pq�Q��g]Ɏ�m'-�.�s��u;������c��4�_{ޣ��_�Ԥd���:W�U�U�k7�n�����w� K��鑔d)Gt��F]q���"��N���շ����6$���c��w.t�#��]9���<�b��)@pu&�u����'���O�uw`�"a �AV(]z��{L	�퍠4rj�$�{1l�����%��^H̬�e�TnG��rqe��8�<^��ު�\���:����Ԫl2LFuY�3e+� �tM��y�Ja�lX��E�~󽻻������FtYE.�n��ʔVq�h��SD�����x�N-q.$��t���wM�
�z_X��3�.��V��H�*X��
m���{�]�;-���S{��ޣ>���m�X4�[����Q5{q?B:JAk;Ŵ��v-�دeW�#�V�*:7_UW���nʪ�R�le���K�����}s�Y�$mo�r���ǻjly�������o��F���@� �Fz��B�]�z�s��EBﰬ��r� 
�+ຣ�����
""#�䥌��R}�~/f��S"���d;��"BL�S|�ݪf���=���ȶ�Kqbf+����U�	R����X�"sz�u.b��Q��ݾy E͒�۩�^�R62C)��]u[]�z��qQO`݁���V���]�:�<#ٓ�Q��e�Đ �)���\�
���hK�2�Ff��*�,4«���+XH��{jf�UN�կ�%���&����4f�n����Y}-Sᜎ���D9q�g�a4�L
j����PrI�.S�vkw�Ҏ�}�q�ѣ�ݷ�t��<߿��!OM��s�]P�ۿhoŋ��f�QV�iz?|�k��><�߭+[�-6%i�Y+�z=��mOSy�w���8&�-dp����}+.E)&r���q��D*��G@|6��H��d:x���Dzs��&x�]ط�b�W�����TvmL��v0��-��:d�9�Z�:/%VG��8��{��Ÿ�]�e����
,�xj��+�i��F��Ŧo�[�f<���Uy�\����W���%�e�>�M�)Үg�+ʹV���He��V��JN_(U��o��eY��zϫ�~��~�̧��H
6��L������R����$,�R�PPE�#*%���)H���U�"�aXT*KFX��j��l""�����0cZ6���Y��|�;�i�,�-	f;׈N{n!���C1�u��W��\C�� >��f�;$dג����;�^�<uyМ����5�oM����b�moC)�Aw9�����#��nzB�;3��꧗]�?8|M���SV���:w�!�L�-f���Μ��Ra3���Nip�����	�t�UW�}^�Q�	��ф��n��5��n�ֈ�<����8��ld��ܮ�o��e��������a��_S�gF�ż�[����)"�����법����Is1%��{���uE�W�ہ�m�SjG"��q���\7o9[��](F�e���ve�N�-�w�G�G���7�+H#>��V���{��9����ؗe[f!% O`�V�{��#5�aX�,̑K߾�y���mn.��!���j�(��Gtڒ�+E������1�욶Elp]H΂��S��\{Ԕ鱆av��c���ޭ�mw:z�W���(��՘|g�g��)V��"I�T��˖�,�r��Y7��Ʋ���UB�|�VyH�}l�9t����	�˻-y6�ms����r���Cu}6�R(w��������_'�Q`�U�x�(P��;W�egP�do�3V��q��q6��m�e��Ӗ_0�u6w3�,�|�}^�O{ޭN}��ꪪ�w��㹬ˀ�D��U�m5��;��y8Q�t��V�^yO��n�|��k�����x�P�����{��d.]=�N�]��"�>���c�`�v�Y��˰G:++�K��Ts�G�3��]��u��������Y~��W�h�`�� ��nA7�RS.u6�Tŕ5�����I���n-0��+tUs�@�b�+s.��G�ۚȆզ�v�G�����-Ruu)H��u��p��V�6�Ts���ۯk��|��k�
�B��P�*"�DAc�}�~�\���*T�BsU׼����F����lj�B�r�mW��W�^����@��u��xV��/eI�>�K���V��/I��2�-�Օx�p@IP2��ˇ"���{��j|�����uQx��L��5D���T�9�e���Ιu7L��3��:nv6�	�MQ��D�@�G�̷���[f>��Hh�l�d���={~�~�e����zy�K���gZ����Hj�z��z��}&���
�i�M6��R�0)�-U���"�v�ͦd�������'��9Aki�Lc��Z�����Qz;k�U,�@���ǎ�:v
�g��\���N���P�b��p҃s�j�����Xl�-^Z�#��2A��.�*\d�X��n�F���&U��l�U�����$�O{T6d��HIp��R�W��%)�W���{�e��.jS��F��\�Pp��^�w�d�j�qO1�����[��Yͷ/6��y�^�V��ޯ[����������\[/�o8R���5�̚j�u=�����z�֣�j;��˫����n�;U:��������w1)����R����N��L�.ݗ�uܳ�Y�qN��p�����L#\��0>��}gr<����F�L���������1����l=�}�{{ު�?��SՄ�}0��܏�u��R.P4 x��������=}Hr�V(* �5T(|%���b�)��k\�3&��]/�Y��Z�.&rHݝ�ÏW k��.���q�$�鱷��)�V+9e�M�2W^ݔr �cpλ���&�\�[	tD_G���1��R`�ޭ��<��b��5�Eu����$'u�H�Hd�FқX�a�	}�UUx}^�����W�L��ⷃ8�_u��,S�j��ĝ�%C���az5m(dr�;~��DB)!$�}]{�����ȩ�c
�jH�ޖ,J5�K�� CY6�DnY�;"�p6�wު��{ޡ�����ȼ����h��PU����I.#f(�"b�]���S�9���r�΁��苷=T#�z޶�<.���Ѱ�S"��c� ����\�@;!��k/���9�O�UW�۟6�~�7�~ֲL���6V[B���Uike��J��B��d�P��X��Bґ�l%X1(%��1���̄�LѠ���m��|�]��MuG	�,��8YWi�jؤs\�+��Y�폻l�'��Y	����N�-�1Φ" Al�lcw�b�G��Qr�O:�� �����0�bҖ���b�X+X��D���8����{��1˕k�Xqv�n�[mg�{Gv�)v�f��Tt@��]���s���8��^��j��������.���J@��P8�d����*K��>��[�h���W�2痽�{��kb����8E��hwYuv��7���/+j�$n�����="���M{����S���c����F���l�7j!YnYb��)ɮ���2�n���ֹ҃j�/v�\�n�}� @�  <.Nh�"��Ʒöй��֊fs�-s;�S��r�v7k��i_T�^��L��7�]qg�`*$��8W����}ZHWЊ����i�?YXUJV���\��S&�֧��n.�\ɮ�u��7X�3ae[O]0So*��Z��9M�n0��6� *�n`���,���Uu+*���|*�[m����2E��w��m~VtT/2h]p�*(��G@XKJѩpE�����vj
lB��HǴ�5���շC��DUN� 
�]���խ����`]b��ѵxТA�����yxk'Z��{��$�I��D�딂Φ��>�}�vk��:Ƈ(Q`��W�sn��t�ʒ��w@�t0�R�-S��4���I ��֛U�s͞��Y@9yM�\�N|>���@���W41O����J����s���Z@@nS��4���h���s�=�ڈw:sFCl���5������[kfr���Zz[���i5�W` �AQ_�x�n�J=�D�B�or�ս�Ug2��ή�<WRۺ;��k
%�2�hs.�|J�A��UK���,�����N���r� h��P�5���U��*�V_��ѭ>�V�M�7wUxP��p�g�.54X�])��+���e���s��O�t,�w"�Z�^����1H;Z��C��,.��٫�wg�~�����n����F3����u��5ں��
6�Ob4D�z����,L"���j ��&�yq����VSӈ	m���&�nMR���0 ���>��d��C:;55KVc/71]���]�@֍ˀ.};P`�ycΨ
��PsV���{(�;Lm'���t"�cE��|�`��i��k�|�:�n�_�ɳo.���n��(4�q�\__gX(r;�wb�ӧ	CNT0����4q�*�7�oŸ���<9�m�Vof[�c�7� [�F�V����Aܫ�Ъ�G�� ������q��]ʯU��J�x�ʣ���R���i�(<��-7�Qr��H�.&�Qf��+R�z���un�ň�4�>�Au�,��'"��Ģb�RȎLCi�wc!�9��c�m���D&�tH'Gd�Zi�{p����T����@˽��b����e�N�#�W;�F $ƒ�����95Mpݠ��]s]�y�V�jNu�}�x��ko ���H'�����}����s���N�ֆ�Yc��j̈́�3�1�ϫo-�W�[wq�ޢ�XWm\�����q�����,������eq"��Ț;�/_Q�[Ū�}B>l� ��>W��<�w�5�ͺW��t6�+�2���õ+�'T�9M��T(Ӽ��n���/1�陣��Tm"�����k���<� R��G,���8c�ޝ�j@� k��{ѵ�Soa���+� dm�W(�(���ɝ�*\�Y�5�G�.t�濏_��Ͼ�s]�����T` �b��{��Zgh������p�+J-ʏ`�Wד)�:󣥱��6g�&�C+{�躗�bx�&�uVm�,V�������V�?/s��׌�3���k��q4!RTqK��v���m���}��LUʧS���b��oҚ��:02�}�K�u����ھ1V<�zb"7v�]�V���9b;at?{��-����q��������r��PJ�T�hzf�2�,[J�.ѽ�r��<vz��P�`q药D{���;��\*�w^}����}׻�u�`�A`e���Z�dbAVE/̥2��l�-�0�;A����2J����H��}u��>��z���4�o]<�J˱mõ�2���6)ʜZ�r��6㵸����S�+nt�̪Svb����������Q��|�qqB7(�n[`̸��7ti�S��[����S�9��.m�z�
����Ul�B�<��ϱ�6�)4@��f@S䝝t�S{OWnWb�����l:�dS(�9�=���S��_���F�v�2�bIG)�	�Y��'h�F�Tq9�+R=
vE�c���#8չ����^}^��Қ&Jv/0�+�gNs\9Xю$��b����7;/6�uܥxHN%�q�=y��r��ݳfr󫖒����4mv1�\�n�+"J���j�N�k������k�9��w��0�X�$S��|6{S�[I ��,$m?w����~��o�w���>��M�J����7.�֫Y�**����a����8Wj���@|-�ʹuƟ�R�8b�7����:+�DV�G&9.�OGJ���OdyjU�H:Y�;o��^���gދ�mF��;bsf&L(�y5h��Z�r���c9α�.w*(r��:�X6�=α%�a��0p(�<I����J0���7�3�S��%���P����J�!��<�wh����ո���t�O���z>(���[LR|�r<�d)[��^�����{\G���	�G��.�l�Y�Ⱥm1M75N6R�͹�e���/��=5�K��"t�;/VF0 "��1�~�>{�9�F�Ғg#��S�� 5ٱ�.nh�Ζ��;��*��~WWB�I"�"�GT�K!Ykd*��`i5¹������_\���\�fTX{)-�p㬮���,ހ��W3����u2����F�%�ru���8)oE�i<�����}�::Ky�.<�^.��tS��q���C�Hx��8#}y��.b��wM��olJ��A�ꖔ2a|���y^��U�W��&�m���̬�ݗ�)�_{��Ri	X=�;��{�޼Իo��A�S~��W�T/y�{��x���SiR0Un[(J�k�%�� v��3�/-t�Y��9Q�aQ:��A�C��b�����Jy.����q��f��e��9q�7�ky6"u�ڤ9HL��|A`1��` �@X�=w��>�����tﱾ滛���(sUr��\�1ϩN�UP�l�ejJr}*z��D<��<�[�����������6T��,��1C�(hMh�DL*LeV1��2�A�(��	��.Z��"ѐ��2d�K�49_?�**�mZ��Y�,>�[�E���;�.�8oim;�XrwK�Pv�d�5�}�m��(/�jD ���*}`_��3;:�!�q�;�.�
��ʽ�͕��ڄ�&��Q���{�~����obZ����$ ���]5]�.��s��$�JuN�z:�9ZC.& � ;.N���8�RY���7�Z�ݸ�Đ�K�4�$��_+����wՠ��'��;9HgM��]�kI��2E�X���#ν��Ԑ{�P�rV򀦦sBj���D&��\�r`����oY�ش��Wb��.�������w,O텊`�Α`J2���nvh�lJH뒷S.l�}��@&�`[������=�UO���5��ǭ|��s�/y��L�r�¹�8(0�c�ol�y��5�R:������IJ���c����B1�
" �ŀ��z4.�u���9���y�n]
]����b��YЪ���W��m=C�m�D乄�V����e�yx*]�`�4�Yc�[ȓ�N��F��]l���-{��GL6NB���ьL��
��i��h�L�Y)�3/\���#��ެ��<��~�o���!�s�̼�cC7i]��SI�Gm2a���W�/�[�Ө{���ܮŪ%����ϵ�Y�钯�}�l�u���qNgy턫#�e���Q]9���u���hӽyKq����@��{�aX1���>��=�)���'y�L}҃wk	�d�rڹ�u4�:����@%�9Nm/{�����+�O��u�j���U�7m@T�� :&j�Hxf��pH.ړ���NڸoꪕRQo��Ws�����6�w6xB6@�e��zNI���Y@��@
H���gSњ��e�� ��!�׍��cK����i<�ZB"7�u����cތY�ɝK�*�wsn�\:�ѧ}�������%;��[���on� ���u>|�ݨ�]7���Ui����oADTī�I�`ꆻY��Nsmm{ު�jl�����R�����UVSi��.+��.��˴x��\Lr��6rcJM=�۷�dL���S��*"��@x���q��)ٕ��4�i���DT}���r�=Y30HJm-�u���/y�DM�6��z�Vj��l_ ��A�^��QB�*%}���t�j��@�"�舎T�O�f��J�{�EM�G^�����w9R�xD������E�a���]+�	N/]{`��I:�>����&���ԃlR,E��cnAa��a�yÀ�<���R�ۂR�( ��ց׼Nnykv��\�l�]�z����
�cjŻ�qt3��F8f�5/�IX*�����\bf�4u+l�M\�P@��7�3�>����9̨'�̹����2M���N�g�,��B��U͔4'&�ᔜ聇��O�E	�`,!������ox�8.���<v'�.��Og>�3W.'a�ݡ��bR��*�,��/��_z���^���j�/��$����367��p;Z�@;�u��:ᩖˌ\� ��ݴ��8��:Q�dxt��{���xL�M����+d@Y7r5sJpnꔭ������A����p'zA�P�޵�wEs�Cb����I[�����'1�����n!̮��e1|�EBW�7ώ�X���)r��ZUTE�f\��\�I1,RE�ILQV�Z0�-PUKL���~����Yf��IJI��:�8��c9b��{X�j�;��g�P/�ri��^�Pevn�4V<��Z����ejK����z"���Ԣ�غ�,��+�L�����6@b�q���h}覅��B�Poe&���.��4�el��DDM}�����7��Z������;��>�����6,�%j��t�x���X{va�D�p�d���H�
S�����G��)��}�r<�u��o�9�>��H�S(�<��6�wH�w@�y8A�!��ޛ�ہ�����\����qd�}U_}��戴B�$9t�#�����P}�����^��a�]I����p�#)��4i���I�Y�<�_1����}����qOa:^�x"k�Ͼ�z�\�-��� ��H	�;*	��9=�A�u��u��I,`�E��@�J(f��#�)�N@ߣ���w*3�?�(���Ӣ�u�v�ݚ͞��I96.��C/d��5� B�X�,�`DB1%Beգ��������/EuB*�[�����w[�<���ާ�عZ(� �Źj��ɀ�g����;S��wS�	Vw2b7{{$\�6��^�;���u�]���k���ہ?�@R`{�xxD'��)ճL�d{����V3'��F%�(f�W!��g�%�����86�mWI���E:�:�1��R�[gY�84a"""��z��Чt�o��%�Iވ���:jv�@Z��5� �AA`owfum��h����B�1�Թ�(ǂ��&2Gt�T��0{��{ɯ��>�u������;g(�2�r1�އ\���9��j�$��=	�P�_@��z,X�-U45A=��n{SY�X��DYd��h�&~�z~��ҙ�g���E/juB�e�H���^��>�	����`<FU]~�P�dYj6�X�s_G��DD5O�~��x��Y���L����Lh�Bt�Є��¨��Zָ*-��L:-����.���ޑgk'J�
_{ޮ�zf��A��}`dK�,Y�l���_i=nS+��_���z���`��
5WW�\��s81ӡH�)o�E�6+z�;����΅�ff��l�B���$���F�k��>2MfMu��E wt%�&�B��_[����0"��W��ݟ+ŗת�K��uN�U�¡r�e��,Q�bDC�Zs��h�R�yܚn���V�᫗�κ��4�J������d^�/�R��zv�uc.�bŉ��jv�|�{�k�gʬAW�P�Ld�y;�AUT�ϽpvZ"��6�1PX�~�����`"�Z���W��w{�G|BL4��������
ȱjѭ��Y�]��DKB�b�Ѥ�`Ȣ��u�ovA�w����o��CbT�m�c��q;����6��� �R�lڀ�}�Lu�w������ZEP�+r���W��Rn�A&^��Q�j$w��5��w�8�zͦ��q;�󯷯s}rv�b�r���f�(P�X1�ٗ��ftg O�p?cU��T�1J��2:L�;u��)sO�r
�z�ì��sNڂ�R�w9�!��)������k �È�J�O��`YD�2%�Ϲ�;����8՜���Gwna\���F�]h�>%R_E/���Z2���j���VL�0�Xj���\�R�évF�t�m��u��֛���@�����
4'msi2{�.����.�X��Cl�3 �NƳUs�0�-�������%�E��Խ�]��4"���0���]�.�ƭS�L:7��d��;x��":��V���@ܺ��K;��X��8.9F���P����G��Wh�ohK�`W6��u�1`����n櫭�q�!��E�V���iS�V�t���v"�so�Vۿ����=l��$f����	����:0���0i��Pd.��K�$Y}��N��ݒ�;�b�L���̲if�	&��zx��[����%�Cm��M<��i�ڮ���h�Ip�T	�vӥd㢟:���[��Q��*N�l삥</^:�=�u)�����V3[-��9��:D���r�Q��-0��bȠݩ����&�i�9*naUIR�۬\�j�c�t�kP���O�I.�ᮗ���e>�z ���*�UjU�K;��)��L^]�o��&��ѷ�Q��m��G��X��9�"�.���L��-3J����7%1,b���t�bɟF��c�u[mԴ�yILj��t��H���u�@ '�����6���ho٩�tk�K�l�ܓ�MR���*�������vt�f��o	���c&�M����v�9�����sHTH���g�\U�X󺠘��Z�nr�:�a�3u��P�t�huL��PUmh
��l��p����gG�HQ.7<�аȳ8QPb:b��?{�q}�}��~s ���e���n#:�����L4�֙O�?�h��\��X��`��R֪���i��z>�=�@�>Q�F8*������A-v{i��������O��d�����R%ܗ�0�"\�;����,�G������˛����>V��Daqa�:n�i�N�dOp�z���n�U����[��*A]̇��nw��+MyuB���G�����+�~�G�;g�ϛ���N�lK�:m9˩�G89�~eu�N�j�"r�my�ɠ)������9�7����ǿ� �,`���� G�'θ)�~ju��R�Lu�Ҷ.�Z��.��,Vo�z)>��\�`5��V;�Zs<n���'�����,;�~�����<c�k5ow����[Բ�Ua�\e�%�]��N�:�*�b���`ǳ��5i��X�t����u�.4�q�<�;]��a��(}�}��#�U�i1�W$G��\�d9�����n��
�\:#8R�C �t_��p E�͙�}���t��A��跒>����ψ�:�!�ɍ�S���:m�I�a,y�!H��6 ^#{6�χ6�i���zM�����Q�y��2�|1P���(@���\�a��uҝ�nwH�kgQÓ́P��۸�$&Yx �G]H�Ҥ�<��z"�������k��{�b�Ҕ�ݵ�0�IYI+���H�rg�vm*��hfUe�~w��(	s�fK%B�CU]^����B��N��Wz6N��F�g��~[�/C�
�]؈(N�W)yU�. �J:�uEt����z=���C��y/�-���?G��'>�T�fE�<>�`bWT��ں	�@R����V�(���*��}������w���Cm)�vw��QT�B�"�)j6�(�v�h�BT
46���=o�r.	<��!.}7,�-�
X�Wm>��t�jP#�Q��K}\1����SXy5Z�q�`	nW}�ʨ�G�S�����|�T�ml�Wj��b�L��*ya+��;m̪d��$˵K��΍�g���6���5����x����5iIه>����Ѳ�G}@���#:�Ԯ~����[��om�c�i��;��&�,�-&���.�,r�=��;+�/c7R�R%��Ì��{+tޝ�e���������(3:3�mk.�����������0��ʊ�RVM�Z�{�{�M6�'^�)�w2�5�G�#��� @�(A`1��������z9�����}�� 5��G@���+N�RB͔I����0�Y��2����ѵ�{G�՝��5�����"Y�{%����0�� r��@w0���W���
I��uy�N��q��}W��3�=�D�:�S�bcB��ލu�EE{� �Q?e�0d��")H2 �H �$A��0�}���۠+�5ʠu���K�4�m>��n+8bN�8r���_J���r��X[���U���mQ�������y��F�<2��&����V�'���p(:�
!��j��h��.��a��n��I<�Q�S�*�v�f����l�&[���!9ə�eLo�����1�)���`�U���{���AVt�t���s�S�Su5��B��U�<��۸q%�Ts��vKÕ�D8��9����>'w���ts�� �{ѹ�?�$K3*V��n�ۇ5p������Bp�I�r�����p@L�	��Dj~c8[7s7���a��E}|ٌ*2�9[H<������Y��+��H{;y7E=ʻ.�\aEfSڇ�T�z/#<R���k�=��hp�[��aM�C��C7&��W3��s �X�s|^��������PP�S��^���#�:�g����{�7�)�l�G���>�:v�S��Fz��9�mq��zV�~C���̰��,Ƽ��Q'�	�fa�$bH(�.�%Ld�b ��+�d�O��Tt/�m�l���Ɏ�o\��D���v��K{oz�vܵ�0��V�j�3�Y:�]�ǯk��Ur��o+���+kT�i�#�_��߳��g��9�k�d��$QI����� �n~ܐ��[��s�gB�|}�G���� �+�=ÉL��\�;�dF'M��r�X��(��������L=��(�7��<5P?Q���e��]�֞����B�x��F[w�
�!Ē�Ѐ��P �o�;c����l�����,�� 
k9��W������ĵ�d�ѫR�i��ՠ|�H��!A��z�F���E��0��p��DG�����?a�"}�/^�����}�X�3J.�υ��VD|1p>֥�	��#o9AL���]FmO��~���A����0<�+��Yߵ_CEݎT" ���2�\D�e5u��yQC$0ú//��r�+B���ڮ93��{�ڑ���s�پ����5��ϽM�ö��%HB�
�(AB�JZ���Nq��k4��.�J;`$�vj��闫�����f��u|����<O�/�=���e��(��3!�	tړ)1c�Lp������X[[+�n��(e�������/"�=�VW 7\�HnD�{��=����3����v󝀦e��=ݕB���oi��\;�rMƐ��j��;T��H�|�A�tw����~��{����W��u�ù����]E�Gv}Q���Q�<�Y1ǝ���pV$x�g8f���ކY68�w��;G�0��EJW�����"�7�tv��@�*�P�
�C ��J�$������z�`&r�*�@�K�<�1j�����G���e�o
�l������8>�[��)�@@4ء�.��m� �Se�=�@ǳB4\Dz�rrzovCg��������������F�r^16>��0����P�Y���m'���dJ�$��$�A�U�Sbs����5���W���%G>n6����PYI*H)�M4Lh���h?�dp�YvO�?;jR�tuu���\�[�PK�%q�0��WM]�sof(�<�9��+�x
�u��TmF�xglT�_B����&X�%9�:T�����(=R-Σm�#��U�1�Nh������t��	���W�@}|���)�߉�ȡ��������Ș���V���IA{�7f3�j{��
	I`�Oyܪ��M�뽇)�q1zc(�|n���nq��+�&a�ܗ�_�U=^�^��������]�2�7�fڥ�kʹ�/hPTd����w�����f)����^���o?}���pK����n(�'�yt�A}B�~Gjf��,�<ܗF��MN_'�uun�ۭ��8F.4��u7zi�G�� G���o�`'�F�4�I����'��O�����C�2����Ϊ!ONW�1"�{���c���VGV���4%Gdྫྷ��`�R]z"/�D
{~��󏲊��#I�53�9�JȤ�"�MӞ�X�41�=8���z x{�,������eg�t
��*�^E:NOm��k�C�>1k$Y�m�%ou^���<�uČ�R�S��13�A�R�c3z ��0�u���y�'k�g��$����:V�\cj��zc�m8�ɟ�ȁ=��_]-zպ۞$�S���J]���%��3Nmk�b�z���ͫ�.�2��.m�d,1�$e>�}<vP����"�N+�)�?v��:��-�X�������_"�A@� ;����w���-�v$�CV;�x<�����5]����w��-���s!���&��^���Rhw�UC�z���-S��}���-��U�"@���=���r��:2(��#��S������oc���'4'贙�ҹ{�QR�s�v���5�3�U:l�ӣ2�K׾u���M��P��IX��W���5�E<���w�j��\��.�mV���L<�np�{~�ٖ,_t�;����͔�Ŭ���ll��u@}U��W@�?�8n��wN�N@��z ��dRH��1�E�"B
�bZY"
�#B��#D@BFH�@F`��
����?���kE�%Y5ok��\n�1��W���g'���c��w9Xt�w�h�+�ԫ|k��u���-�Ot�Ǩ�UVc�w�V�70J����C�b����cc�&B���ވ�B�-�v�@L��'�ɴP�����!�����De9���d_����ڜN�|�T8U��i+��H�� j'Vi:w��M���rN��K.�����=[6�G� ����P�T�Q�����
X�RӣP��\��!��_-�g-g#-�D#�Wa|e*f�m�}������o����!y5��T�V�,�����.��m����ܲ�x����9/�g,����P$C�DA����pĖ�9O��U	���\OK#7�h�n�In��*�����=[�
�P;n��O;�z��(��D�Dރo�[��b�W�Z��3vO�O�Fݠ�o�
(���T��)�,1�ڨ�">�ϳ�y��s��}d�yI�U��IiO�?}�4��Li��#��/���ɟ$�3�j��̘&��H>�	V�7�,Zq�s3
*m�䪃|dy%m'�_PܑJ6�.�[q�*�-�%2������4�[���9�v�p��*ճ�v)o-�!���
��<*�y���B9b����^����DgU�%[�zпz$��&W�k��Z|�����������u�9���k��md�]���t��k=ɇ��ZʪԼ�것UK.��o�ӛ$�+��{3x�h �;�Y5
�X�Uu�	��W7R� a�A�DfL{@��V͢�����ڋR^�*��o�o��z=/��عO��{rc&��h��*��LL��}"'��E�q�+2����e�{0u�]��߄x����Ҽ���=̼�]kO��Ɍ膽W���]�s<���:����x|�R�P�qAkX|�/U_}�xKW˞��;����u��_��g.��Fa�k��(׉:1xx�|�j�%+�:���8���Uf�/��1Q��@*���[Xbn�+�r�.�2:pN_s�N�^'y�Y�7���u�r��y���C�
  ,T$K;	!�AbV��0�t�(A��J<����v��6��uٺ�{η�뮫2*㙧�.o6�������}�+ʵ�S���UKo5WU4��#(V��D�d4SU)mm����8���j�՗�PR�I�΋U�V]��h=n���7{7~�ۢ(RnS��pFq����_\8�R�)����\�eQ��U�C,1a���g.}�k�$炙�q"p"%�������7����ｿg�=�e�!�"G5Mr�<�.g5s5��ц�5�Ȋ��a�j�1^o��T�W]�Q�P^�^腙h�\��ˣC�s(�;�֦(����iʛ����m��&6RE�Y������iʜ����u�+�iϳ9t�3������{32�����ʀ0k2ϺX�1�\>2ee��@Tm������^4T�7\xkϟwq��}�}�t�{���wǖj����4�����C���Y�Wuww���Sh��e�̛��.Am޴�U�9�d��߄�giP���p4�Gi"'�ǲ�S�o.޺����­`+���T��*}>��ŸU����ܛ�d���A�2[�6�q:�'{�k��3-'��Vp�2��˙��U`S�Z��;p�m�W�Q�1`���G�G�0�;(o\y��:9���B�ic8�S[	�ϵ��"}�o#IUׄ���Š�,��ܝ��n��ic���[r�b-�{(����i���3@����-��m����:a&�q!�s(N�ޝՀVæ��s�ݐ����͹a�;�<Ilj�E��m�=Yr��N�1'X��}��Ɲ+"{��]u�䎷���t2���u7���r�6��7�I��!�P��N^8�	i��v(��{�%�Y�k
���\��k�]lVm �6���(!ʹ����S��@��m�G�U5�qԳ��Ǘ�gAu�1p�zfX�=�F��'8���5����5A�uAY�b��!��Q�ln;{+�"�������;��G�]\oy�w(L��@�i�Un�f��܊�4%moL	����JC�0n��(��:����WU�`��(��%��Tj�5z�&��͹�Qۊ�5ۊ�F�V&� Y�3Q��	Mzx�<����^!�v���kd'[6i�
� ��Ԟՙ��t�յ7$Ȏh�6Y6��ҮF�.a��)�k�.��b��'hr
�bd�q�-��L���٩��B=,mg����kh}�g��� �&�����E�"%�@�y6J�Ct�=�{ׂ���.�fͺ�U���y-W*4ʳA�%�+�4�m�)#�t�m�`6Pt��P�b��Pۙ��7��uݷWw�����(��q�9} ��� g�:���LN����:�PJ�~��(F�Q��ݷ�����W$3�9`@�D(���2gW��1�-�Vs=C=��e���	�D�f���P�˖*:e��w_{~�O�q%�i�~��ҫ��K{'�m%S�b� ;��QRȅ�CPv]�w��W�.8v?��n`�]��?��<�z#�3�z�,���IE�u ���i�����(���t+޻�\��.T���� x�C�(k,�\��qpr��H�Z�6'�1�q��s��i׽�~=9{�43�_�SH&w���=E�
��	��xb���(�3�o����m���KG���=e�յO;%8�Y��"���2��k����N��W칖�)wi�������~����}Sh�i�2�hFW�4l�%cY�2���5�D{۳����������%٬�P���@"� L��#���e�e���H�����}�QY�Q����Vu�wYY�.}�\Jq���2���Fe5�rj�-� ͞y(��d�����؝�P���Crf3���D�r�L'6��ݪ�Mq�d��/.Xw��n�`� -�@0�@���h.�z���>�G���M���*�V�7G2�(�S�<�����t�7 �.����l�$9�=ϳTc��p�FH�
�QDD*�"�|�}Ut�����K-��������j��7&uY`�>l n�-��5�+����v)�-;�y\V�l�ssT������".�8XQ����B �e����]�&{&�j^�o9ܵ:�r9��{O`5C	�P��\H�[I�E������Gf����_ow����+@;�WNq�� �n�ڙ.H/f�7F�H|�܌Y�0�&�+@W7Ǹ{i0�6�q��E�?{�o��_��C*f,�G�:g�(}�>�h����C[T�w��K�:�_���=�iwG�� �X2c
"�,YL�
��oo���{��q�%��Y1�͙�iބ!,�S�/�;o�\ �Y�	��k���N�Dk�i]�Ǘ�[ė,x}Mc�)�u{j�!�Y��T����qʢ���[z�����AibUp�yPԧ�=e���˖-��X��oU�s��.�<��YP�r6"⣻m�X䋰̖����@��ch���a�F.��ʕ�������r��N�M��rU\V���01�Ȱ���*\���=<
8��E�{�u���6;�Ӊ��:/��q"^��d��bAЅ��﫧uE�ENG�%�w)D���-�JL���;Oށ�~���:�6�gP��{[b_�mB��� F��\v�S�-;���b]�8���U���wي�V<\"�� 0�D����u�]O�FL�L�?|	��#�|�+�rw�ݖ��-`��+���6M;B�H6C�>�+*�׮����0�Έ�}��\.x!��`9<�_�׫����3{��$Da�k@�Y�6�Z�٘�nR�G (&$��-�R�$a"�82�`�a�liaE��-�쬑E���+aK7i�k�iՕ�yoz�4�{+n��r����o<�а�+i�Nf�)n�'o���brǡ�Վ�7�nvPr��V�A�Y��	�֛�n���-Q�݈:"�b#��0�R�tN�pY'��=����PV�����:�Ϯ���Ku�X�(kU
���%�Q�Y:`���u�ieP^n�ćj{<OoEOmD�ӫ>��@��XY�ܾ���#|0Ё�it@��]��':>�5�[���=	�-k�����k>�fH ʒ���&�舜n���}/���g��%�J����n�+�$T�]&p�P >�\�����gF��I��E�E6��(s-���}07�ӳ�*L���Ʌ�����jx�bS<�d�8�$��l#��)�ء��Ĺf�}�z ��pK�uEA+T��SKn���锔�e�X�9v�k��|zi��uok��h"1l�D����"C����)�:e�����{�h��փZ���") � �,YH��30fZ�4�"R�~YA��J���9���6"��%ֱS�#�:Hr,wrf�H$���u�m��YKC�q���@9��R9Gy��Q�9�w����h-��w?�b�����'��
O]�9��l�-�>���G��kV��ـ�e�Tu��#֧�t�й�������Y�z���Ɲ̂T6d����s�S�v�Y�omT��!Bz�|��U�8]�%hScmB�����C_{/��M��̋��=ab�����k�F*i�/fT�4ĺ
�N9h�<lXvNd�Dz=O3��kkDB˔ɑ�������E*�x���5�z0E��N�b�r����]�4�����(�'3��T����}R�t[\�Η��x[�?G��D��S�d�?�9�uT�eK4w*� ޖ��M��֠`z35Rf�e��w��<� ��e󽪥����g��2�qk>ģ���N@�V>�E-����l	RA�{�����@$� �@��VwU��pr���7����^���3�I����keWq.��9��͝�0��9�+a�q���Ք�:,�He��i�6��;�V.���]OZ���Y�ۿG���D{f��>����6��ϣ��FvR6̇�G)�.����9�����̕r,�9�!#	˭�:;/��*�a^L��F�����{�x�'릕;�N�>��"�N�W��2�s��i [�Tq�N��މ&F�Ε�t����J�
g���8��Ub� ��2�������Ҽ��P��ע%��*���5��x�s�m��V嵞@<;�Ú1��xj��Y�UD"���5��U?oF"S;9R�2����s4%��靲���|xj'��G��+����.��Z��%EL��E���2%L��z�~�/�|+�W��D������ι�P{r�A�c�V�E�܏.���I2�\���l	��҆U�D���:k~��|���@�g����J쯅O��  �+0�� 	"Ȥ�"z¤�"��4f�nf��*u+»V�x�d��ݽV�9Zt;n�G�ƨB�ŉ]e^�@ud��Eמ�S�W3��8���P��F��f�O���o2n��S�?��G��!ا�!4%����D�� ��\`�t���\�
��wʩ���qUþ4������x���vs�9n7��:fλUr�Br*�����(Ou�!��Lǽ��R쪴�k��1���z=��h���3��b�׭\�
Z�i+"����#CLN��9�����=cz��J�8w��)���y���=��W�׷��z� �̩��¹�����T�u��OH��q3�ˀ\���c,�U�H�����#�u�.����7��Ղ�eKm�hn�2Y~�s��Y	�`D+���Uw���ؕI����v챗=H��G��z��)�����_NWJ�<Gœ��7R;���I���z7 ��d�*t!�+�2�Zhe�2�8� @.Z!&	+��J̌de`�9��+I-�b#��xk"qc���N��y�>{XxT��_-�̶ڽ�td��b��(�;��&��y��Ύ��%�$��x9��������^Ǟ�X����s�2�$���<��@)��WkyoEZ|]�/K���ގ�XGx��s5�\��"c�"=�DRa}���\��
�RÒ�>���i��lܜ����P0�0�`�����&7��΂{=���1��eN8/_Ek~���d��B��ap�84��g�r�C7f��P �Q,��E>�ƻ4XN���M�T�w�[�����p�~�7�u�o�x�T��| ��x��*�`ӹ�[6��{4�F��I`��qc��v�R%��tY'�.#����}KM#+�p.0^�U�Fv����Ǆ��y�09O(ɰ�`�����{G�ײ���W�k�rX�
W�?!t F��=�&�i�{�������&AQ�Y�JR��Q����X�b�`���f���U�)�k��wg8k�],�:��[O�������@�5���h`R�b�YX;\�mV��8}ў�R߻w���-4٬���81z��P��fp�8�h�À�xo+��c=�C��-`ޘm�|�ɽJB`��3�Aw�޸q#������5�F��oY��l]ȯ[�=���P��0K}|%��(g�#ۗp�|qW}6���am�G4&��i�۱�p�r���ݿ��k*�s*�&s7����L��}[��w�hf���������:6�G�����D��D[�Av�Eg֑��Y�V�%�5�n��A6�g�`:#���W<��舮O2��{��q��G���=~�s����.���pe�s8���[�y���$��&K�����r�F�1��(��z�G{�Sl����Qe�5O�r��Fuz`�h�a;&e�1������]��nu��;��{M�8��JvOxz��{��|'���4E��B��H�k	{�e-����y����ekP�'���^�[�-���ʺ��nr�4�ؙ���.{���Y�EI��(d:�6���K�Dkwl�b�x���I1�ajdJ��S�C�`1��q(�˩	�UAb���]���Z���ɭ`6m�
�HS<>��z=��)� [gl������R�R��4UEc��)C-�S���;D ���&kl����=&����U�6���!��������!�j�S��l
�ė$f��&.���'�]�<�zs�g�;��G����+$�(n��DE�S�)�ND�j��ة�������v��u�5i��cZ�΄{@ֳqG��^Gj�C�V��A̕���GϘ�Wm��O�#>?��������;�M�չT05s����\�6Wk��j&h6���gU����am]8yj�F�u`���g"h?�B�m�|�w�
A=�x�� �.��R���Ìy�]�,��_z�'Pf�Ӎ��O��Dv��ڱ.�}4|D.\�n��]�s������"��(�p�ҴZ�m�+P�xo�J���t웽N��MQ=Fѭ���輤�-��˪
��]����3&��{4r�(�og&��"h���t�5����|�di[#��^7x��J!o9�"�ҙ�5�k1f��t���'#��[-�PU����w��SF�~�3�e�2��j�wZ9vw����D�l���.9l��Z�["��߯{/-��k�Kҙt��	7�kB��m4�0b�Į���h��f���3FV�T��]6�c�	W�LU����È�/�e���d&	߬���cSB��4�k�ys-g�x]C���Y����&��.�;�����}ۚܝA�(C����n
)2��ɜ�V�z�T����f{�a��[�a�Yni��*�ow��-w�g^;+]-d�QXo�]^�/��/*���g��_c��J��n�V�UW�1Hh��ҥ��t��t�8��[�`ĉ��h^�f��S"�p��4�4��q5�h��P�.��]���Ub���7���v����{��7z��Ē�0��n(4V��J�����m>#v2ɨWE��j�W9��
�rĄ� �l"�e`���F��8�j�,[5�+ח��X�y�����[� if<�����3Uh7֤;bN�C����`)�� E7]Օ���-���Λ@� E�K�)쵕v�-��\�:�M�����D7.��f1s����׺�H\|N+֪%�k��ԜsEA
�rKٛY�Ղ�� ��&�J4ʳ��X!�Ј�{(\д�8TLӵ���n�	nVU�r���ĺv8.�0��@���u+�����*�ˈ�T�L�XCn�k�����Ήrr��"9�rB;Xs��\�4�=ס3L���)���eɄ�ܥ�� fѵY-�N"� ����X0/��Q�$��9pֻ|,��gF�\���Ce]4��G��WIcZ���+��P�rЫn�.W@���K�h[D[���n��։�����0+/�U`�AWD��Z�W*��4g7�-�����E(��Rt3���҆���M5��}��^��j됴�n�0����5m�62�u�f �gV��d�(�v�<���h^��_i��u��Ba.Wt!7X
CU��hޙ΃���(��O��{8^���h�Z�7sOtV���Y�����)���&����e-�*�lV�.�L4�����	i�V��KL{]R�N�\�"�����YW�]�o���L�V�W��*��5'tg7��(��B��v��m��q�ϥ��B�8+�۸������V��c��(��.�[��������>b��H�s��T�~�]�L}��Z�U|���XΙ�Χz&���U����~L�8��2�'�ϛk�Z�9[��"X�Ζd�����]l���i�K?z�vT�ݒ�|�T9�.\�&��߱���yE���{w�:6.��
f�R 2��X.�R��{ހ��{ދ֟e'��\���<8�g�L�l��xt	'q�̝T ��l���M��y�����ջw���( (�r~�G����A'�jbB�A��a���ah\;B�C�K��R��OOR�@p�ZU�.׽�;\�6'R��}S�:�_)��zm�13��d��:9ΒG}�.)�{\� ]������Kf���Y<X��Q�ڹg[WqQ�<�8��E����Dr��/�M��6;$}�\������(U
 }	 	�Q8�dP?~���f�9�����+n�w���]���Zy�~�W��z�����r+��t��0B���K�s-��	�y]���X�˕�qɜ��ɣ���N����:;�5	Z|H�=D��RK�3])���O���=�.]�+����{�Znjc3�h��;&�jW0m]`�X5ݫ%�����#�:��\��A��|D���������[�Ŀ�3�a9(6�`�����}�Zk;��8�enIuV�����-YKyǱr�}s:q�ӱ{��
y���.�$��`
w�)[�d�=�GB�.N��9�1���V,��ǔ���5<d&�VK`��{5��]c���"�;F��e�G�>�F�׷�F+� i���Pkҿ#ˌ��ry�T;d����j#�#�����ˬ6�� �Or�-q��E
����%tkx�DD"�mi� �/X浹�wy�H��A.Jk�pp����:�������3%ZQ)e@,0�"1T!����:�)��ZQeVT.d�*1W2���R1"�$����B�111��0k��vf�=eR�B���;|pZ�b�ݲ����Kw�1N8@Nmj%76�Q�N�e�r�\t��f��9�9�ф�	ά���ufX�W�e�*�<Fz��I��Y��Qݵ{y1^Ɏh�-�0H��G1��N����G���e6���Y��>��.����ٙ���ކN:I�]S��B���t���i;,�9o���������E��[ꎆi0�UT�H��
SR��H�/oG�R���c9@�����N�6NΣ!�05�ɋ�$���o\�	� �ۥ[@
M�~������fb��h���Vq9r{	��͊4w�ljn�x�Idvw_��*�M���.��f������!s?@��.�c�_B��ӛ���X�3 ��D����^ّL1���I�8�Ov+�\<�� �L],��Ev��/���W���ND���1�G������W��P� ul���NT��iN񊚝e�K��'Hة��l���>��*���+jADs
c8tt�/�����s�X.�Ouչ��]k� �)B�ĭ�f�ע�ͥٮR��]��X�M鼆���R%�70��1+��)�*P>��mNZb=�U�d�r�����td�o�;�w���z��r㩄D�RV{<%�0+��C�L&����udۨ�錞V��R���]��<I����
��~5F~?0hڔ���`U���t���Z(8��`�.X�W �C���J�D����AmZf��=Z�q�4]D{��G��b�������ƵB ����/�7���I��@e����h�s�X,�����$ɥ�����?{	�G�뜄>[����@44nob�is�-��v��H2Q5�f�T���ju��F�Щ��TA���N�n+����z=��|wྯ�G�����pͮS\��,�F�G=U��H�6�]�(n�wA�M.��z�}��Vd�L����Rx�^M����=��{2��F�����{���ه�E�4��l���!�C����U�"�ޮ�v��gf�V��t�p�l��n�9۷��طN�R#J+��VJB�L�s8�Ѧ�2�	��u~\@�zy��шw�e6+��A�hͅ��������Z��;����C���#��,|�h::/�,��NNb�>T��p�T�� c�lvۘȜ̘o��9˷{��E���,:�ئ>ޏG�;�ﾏ���u�_B9�AĵHq�p*ܰ'���R��G)nm�x��:��ٓ�됈��ۮ���\�@��$l�_C��H��>߮���㗦���X�K4851Q�8Ip�&�?ty��i�pqa��[x�1��d�ýs5���/����������~O֝��í���͝~�����1���F��~�+r�b�ΪC�2�]��;�K��ִ���.^(��E��酇���������&\~��lN	d�XyR�	-�V�]0���r
"x�V� P�)�.��L#-�j�F+�,+(�m��[-*�����
�Y�H��TTb�f-���$�P+d�zG(��bu���l�c]k��v�k@�i�R>�~���a��[�|1�WmkѲ��s��6n͵|��:ylw(�{θ��}w���g�}V̀��7���Z���M�%7Ps_:��)��o��9303�mH8W+�E3�1jw<SJ��k������5�|~�Ǜ�V��Ʋ�2!���Kg�]kfp=L�����M�s�SL�d�0)s�#��D�|P�����?wmh:�p�/�~�Qu�����fL7�2v�D�Nf7�U�t"W�t�*=�77�ت����cR3�e��}�M��b���bj�~��Љ�����;�ȫ~�u��u��N+����q��%4���A�����UX��B/�	vD�^�q�F��*C�$�G�n�X�`��YpZ5K<�)'T�^��h��]��A˂�3�U�J�GF+ M�ޓ1ͭeCح����2�Ǥ��Txs�9W��=?iw���}���}������q��!#$ �& K��1�w7��ٮ^�]Ѷ�^ˀ;�7Qm��ď H�5m�����b\P��у'u�Yۓ��.�*������ˠ�Z�B�mI(=�Vé���zNz�g'Ltm��ܐg���k��A�o���{IPDjIӻ��BwJ�:Q2��ո��1�$��T\��Ľ���@d>�}�����|w��|p,U8��=����ѽ#�����t�+�r��%�ڏe�WlX�<����!u<@E}q�#�4@[��0�����1��ͫ�﫽&=�O:%���n��: "�0O8�9-�,YU0sK�tx��3���3�o@����<03��+L 5*�Ă�	;w��ڍ�ԺmT6q#1�u:n����N��i����v���lD<;W��ӌt��F�f�m굥�F�6�U9A@�WTv�)�ժ4��ʡ�Y�0�J�)�jcY�9�?w��.m�~�j���^�^9��X9J����J� Y�m�J���*E�X�	��a�0$�.Z,�Ȃ #X�¨[F����*j��i}��eÜ�_Z$d�A����_z�:f�R�n�����֛�"6�(_kX�f!�x�o������uvjnѫV�k:5�o�^4�hN�!���C��0�%u	[�w����e,�-n��^왃8�� :a5c�lӓ����"wj	����_;��V9������ꁞ�^�s�Ѻ���i`�r���?��,o���,͈g�ڵR��������RT����]����0��]��:F��(��	�˩K��ǭ�JeaUsɞ��5��f��G�у��v�v}}_}�닟���.@�H���������}�T��=�����U�����jL&O������Ӑ%L�QSLS��p���ݿ��y���G�"��:��,i�Bv�dY:q	U�}U�����y^yw��j��^ȧB�d��`n2\�HG�sG��'�<��Q����q=��WgM8^ӠԹe�APlG�ݠ���F �����=�X�&|H�YU!�	+P���2#$�.�Z��]��p�b�q��Z�!cu�o�,��'%G�tz������w.Ez�l���(+2�9��jJ�
�l0�B��10+_K���}2	�ʱt0g�wޟ�����ﵓ�p!�W\��2����g9�梭~�sVhd<�0�R���#^�jC}DD�;�Hȏ@o�;���ԙ/�9��̋���ʱ������p����Ɣ`�Yڭ�j��U���&�,Ma{
Y�u�[OfϽξ��I����y׈����p��2D�x��o�Xۊ�!]��B�{D�����Ԗ�9�)�xOn���|Ď����ןF�{����G,���ޭ#:�t�����kL�4��W[L'sU��1����3Xh-3�lV�o	uoTt51N�t���%:+~�1�p��o|'��g�QUZ5l�7�c*ᾂ�8tզ�Z�у��垵 mY�*���#�e UJ[�=c$e��]��	�����u}n��:c�2>
UIv��c��3���G�0�'�6��@�u��e�_�Xx �E�a�}��[ZVL���+ID��&V�4V��a���Q��:I�Z��y|�D�0��S�:���>��"m}�6Oq�f�\;"KAS;4��]�G��n_+}��3��t�n:lpK&F�7=¤��X���+uV�F )��^@��UM�D���l�V�&��W��z=xDE�x^A��j����X)f-�A8JمГ���!Н��*������fW���`u� ͈�f̃;ռf;h�G��P�?����x]}6K"�fwt6L8�;-G��6}"����h7���'vw��B�H^�3x��pR��;�$tY��fT��u���1�S˶μI��f�f�=ܧ!a��`ۍ���b�[�z�9S����_}�A�م���#��U�},�dub��
9��������;����r��_�OP�R�����ۂİ��R^V��J+���k���z��ݿ6z]i�~ʘ���8���kR*�SU��Q��Vm^.�w�z���P�ԮP4
̻�r�h۲u&��nwT��i\�cT�
�b�ث'����9>z}�|x�x����!SOn����ky֢�V!R����Ùͭ�C����TB�ds�����Å�E��-�r�V�@�i�#�����v�X���X�B�e�7�\6��@��ox��{��g4e�y�s6���j�����߹�ÏE��5�٬M}�*�����b*:�p�EF��L3v�C*;殴��K!B2ҋ�0�4��1��:h�R�F�m��+��V�syrŖɼ˂*,�{s֙����X�3���ִ;4�֓E`(�����[�[t�n�o��[��=���*��.��ω{to�.��j�宍6.�o�7�u���)�:�sE�n��=�n�E4���Q��Y=f�Q]��Y��X$v�h 0^��7X��݌�PR}�y������Bi�=�ӎ���є7D�j�U��,�T�AE�ֲ�&[�f���q��vt�{V��n&[��'�S8�Wn8�j��XR,gs4��\B4D�	o����e��̬�.�o����:��n�R��e��L����SܝƸ��{�1;�x��av��{H�\,���"`ݙ���s9�"ڮ��U���T�-m��{����c�%>	�RbM^����]p�d� >]]�=�,�sjc���ϺⰯx�����$�6fN�s��w�Z$|�|Q�.Eed�p���1<=z/]İ��M����U��٧BMW[[�	�6�v���"�pҫIٖ/�e��
8��f;�p
c���˲�V*�����n �m+��)�@�J�ޫ�<�_��}&����ҝ���խ"�2�k��[�eyK��ⲵ��s�Az'�|p7����^b%�.���t�nӛ|�n�O)��{}�v�J����4�J&R8k���X3XA���كT@V)��Ǖo����9���^�+�k]�|@;e�`����Z�vU�рe���X�E�\#v0Œ���i��;�����ֺUy�}b��n�E��ܲk`͑"����^����-F}S�^�4Ӛe�!Hq;�]e�4�E��$�3	�`FwE�o��������zV����A\���̨��缙ン+F�Sְlȫu��m����EI�8ܪ���(^��L�3l�.�듒�LD'C�c#��]�G	\�g�����RZ�^'��U�f���N���NȽ�4�'� B��n�!��!�z�мo&��������>�r�O���S*�QpE�1V�A8��[7���6���պ�l�Y.2
q�Z �����zi�?�e�]�Kt�z<��nx���R�'7v�e��3p3���
㥑���`a��l���s��x�%��um}�G����}S�+����='C'�7s�q��Ś/�]��bR�j&t���u_!���b�82��{�Q�Z��@R�&�k�����z#>����ƅ����[��\8��=�J��qɓ�bd��n
,���Ǧ.����|Gǎ�=~�U�@��ܚ�';�.Va��t�$�s�[͐8��R=@�c�yW�<�ۜ��N�-L�'��BF9�`��}�t�� c�:�h��z4){��r+:�SH�X��T��MI�Ci	�R�Hx�z,Dx�>��B�����T���Şc��2#3V���|����\9H�yUs]S�{t2%ݻ��á��R!���oi۬�Q1���K(���B�sQ��m�ޙlŘ����z @�����h"I_d��'x��j���ǈ��l^Gw]&w��ܔ�E��d��@5�z��~�2��)�tygJ��W�߽��lA�
~9}���m�� N���~��ƈ���D#�M.�5x|�����\n����\��;�Z�d5�[~ה����ꇯ���� ���W�Φ���~���Sj�qu`]:��jC���u�����Eb{U"pe������.�.�T�
�����u-�V����vJ��Y-�t�y����Vt�@�#|k�������:4���J#��i�&Z!L�o�~�F��V���(��n��=<�~�»k�F\}��$}.U*�4t�&��΅fY\vv^��^�{ވ5r��I�o.f�k����1�U�Q�tbC����w��}_w���g������B�Y%F)E��U5hH�
EP$A��*��@,�!+%�
A ��`�(��H�$�a+B���6*�[abg�ֿ~�]�u��m/��0�Ac�ɱ� ����iV��C��8�J����懓�W[ѷ�{\]lYG7w�9$+����M���	�tN닞 �<�nsi�ݱ�z<Cx��V9�ѐ_��^�pXT�G�[G�T� �L�= �e�K��e�Sk��÷�m9��<��82nzMN��%�y����y]����DGay���T��r}Yl0Y��e�7�:#�� �:��Dr�2�3��\\�AFat}�A7ên��̴4�W_މ��S��ӂa�!�\6~\)�Fu�T�5���Î�
���a�P�<[EB�2���*7K5�R��!�e�!F�YɄ�*��4,}7C��W�~,e�5ž�3!dw,�Ke�؜`s*-:�(s�Au���v������H�cu��fOZA5�k�Ƃ�3"�Q�G��@�O��}��L����6�D�։�=�N�o�{ZS�"ig��nT�w|���606g]S��\�rW'{�DG����&����~���t��R;�!��)��s{�Y�+`�_!U��W2�%���9���
wnLx��
`��Ou$/[ˎ���|:ַ-3*Cˇ~������~ψU�?^���FA�0�ʱ�r��>+�mdbcv�[�ǅau��#�\z��E}?D���ݕ�9�}�~�ޮ{�a�@�n��a�4S��N�}.��
b�C`�u����p�u��-%�����߫9��O7Nt}�P�{��oFm'Ӹ�Gn��x�Z=,��D,��� �T��e�Q��ވ���Qt�oe+�ԯj��w��!��ߠ��n�c:����:jvx}�yEt6LN�2$6R�j����m:�؝�d�P8����ɾZ� N�k��pcﾬ��YB����`oNcF�+��D�o��u.n�(���+�SL�f�T�^�Z��J�|�|u_����>���t큣�|L&���u^�Ȑ�L��<��-�둠M�Ͻ �" �1��!]"ᔨ
L��f�r�~���]����}w���K*�%����sȒu�mmC�9�mоA�x_p��9�Kx�[DvQ�O"�ͷ*G-f��o�k�y���K�0���O�#��=j�	��r�&1�;�b�Vj��fve�L�%=ᪧr�p�+ِ��6DG���Sםԛ��h�t�É�CM����$���1!s]eɟ�HHXr���n�9`���7o!/��������c*�I6�.w�{� .S�=�E���m�gQ�Tv����TVbh���ɝz�ԱC)�[҉�8��e�\@��@V�X}=��z=�#�kKw�>����W\����ܝ�Y0����xyߗ�н�F\ 5I��MM6�R-L�r�Ig�����;NM�����;΋|B�1���{�w���5�V��O���=V�gӞj���`Ad+[1�E�;�1\�M)��0�wcｓ^����{%����S�<�|�̤؂�����R"B(,��u��Z�������ߴ����x�Y�v	vTh�lK��`�2u���[.<zM�'F�j-u��{�S�;����"�z�3mצ��ٲ�'7U(w���1����c�ei�B��V���l���8�Q��l�Π"�$��靈��r�Io�6�R��kKqIZ�`�8���(�XL61\�.W!�q����-�4�8�S�f}��V�����~=5�Q?qz��q9�;��[�E=Dv����n&�\�-���l�rG ����o8P�y��x�?�S�ll�9m�e�U܈�RP�r��4S.���IS���bLg��+�\C����L��s�j�DM�p
�D���Q�Y%��g��+��f�N*�B�2��fvUE	�c�ںz�B�^��&d�BF�*�'��{'�'轘]��T��/�ݕ�+pg6���xv0nʮ\���y6(s'.H���ǿ����{�~y樓��VʲJ�����V�mh#s?o{��o����ﴇyY�������5<�,��b�7Έ`Zφ��P��۴qC�$�XX.+�W�N*smN��E)��Ep���WV�/�):��1y?y��~��te������ю�Fas�@+/6���}�����B���|�dq��U&eq�tFm����ҏDz���[X�qT�*
~Yt��I��e(k�v(�d��(���>��X��c�6���5[,dt��3,�UNJ��ޏ�""=����|X��O���u}���d�X*lV�1ݟ �-�%�<L^R�׃Q032/��w^;�"���r�.^V�:b��꟣Ҧ��h�.���A(�x���W!���W�����S�l fE��:u��������M�~��ƕfy��|wԵ��JD;޶��;2�S% R��ε��m���!M]���y���5NU��� �d������
�}�V����D{L�:�xVl�6�jʮ;��3����R�(�{u7��2�L�`THDc0�,�UD��%�J��@He
�`�X��ĕ(����bf����3�<}6K0vɯ4їyu��֏��A2mFd��ۥ�.�O��G�u��M��EY� �ĝ���|��m�;�	e�o9���G��L
��I�͙�ǫym��f�t_2\��^{�z�g.u�$�����*�]ήʐ�cy��m9�=rYسK��郉Wq�)茷�݉���U�r86�Zj��<�P4��&�H�6�v��W��e�P
[G��"��e8I�WI;5�b7Ja�7�6��{װs�)^t�� v��xұ<{�����&Rs�07M������0]s`0���P㦴*�g��t���&z�"���h�h���'���	^�G�z2^�?NH���!U��Ȏ�!��`LW3C}��cfzѳ�Y/M�C4���4���ʦ-A�.���N����J�i� ����mVH�78f���!���jT�SJė���e�D�	M7 .�������m�,������FG,$�*D+�.6�3~�bb�w����g����+VV�=��QV
�I�ͭ�\�j�i�ZJDl��0��<�^e)ղ]^��<�l��^�&�V� ������ye0m�{:�2�L���
�*z�Z�"K�HHoX9�ba��W�G�ட��7=�>9��`Y^�G�&�+Wآ�$e���<�t�c�4�ːd�<�[;3գB�A���u��+�0������ ;'�:���
=�u�{�X1���/�p7��6)�E�[Ĩ��@p&�kՇp�o��*�y�~��Bɟ�*!td*�T�3��%:JF_dPwtĄ�Qsb�i0���*U��t�p��i����uTSbL�2���e��ѹE������2������XL�d�.��i:�/\���n7�3��g7�X����7<E:@�{����P�2��W�r�oخo�,O����
���ca����c�7�aXF�ut��[=|K�w)<��yʹ�8$uQ��rcoZ��r�L�ߩ���r��h]]���9m�b�'w����U���]�|I�Q��i�r� ���tn\
��IvaVuV����a��̙Z�K���uQ��_�!��q�)���5���a~�&�͕1�!�^Lsq�O��zrM�}*����cw���$>��TW�eT�w�D��}R1�'-�ΚGvM�`��\��Ft�"K�#�Ỻ<٧Jf��9���(�y�P���{�DQR�n�-x�cuظ0^�2nG杕L�x��
RC)�3���sh)�ݜ��X*c��4��O#O'22=�D����ٿ����dwt}�?m������r����.(�^9��>w #h�t�`K(��������s�ud��)_��qnX�����2}�֮4��]07uZ�.b�B�k{m���+!��;ʢ
@\^����4XR��d�~��UUU5�߯GC�*ղ�*�s(��d��F��DܺŸw<���Ӗ�tq�O:���ĺg�/v���e	� A����p�5���\�#S�s�U��j�˕�*b���Ê=���_R�T�� (��Tz��p�� �u��_"
�V�@$�7�X����5u���f��Ri������mj���+[&wWS.��c�2�K�9j"6�J�Vo6*"���V�v�B�9YI�2�[���վ�k}�*�����N��*���>F����N�[t�[]�۔q�5�)�hX"��%�_3*�i{��(�n4�/�ШiuBc|is (�o��R��7���9�ZS�&3��9�ΗZӓ�w���3��Cv�9�`����t�������FJ�@�^w�6v�.(��s��׻���(;��<N�|������$u�l��
$��p��)1��_4�4ʕ6�s*����\���ӦYm���:a�3J�k�:U���p.�⒕���sB�Ǖa�D���>wΏI�����iΘaM\��pq�umǩ	A3wW(0�H�y2�F�a��uL5���n�����/�������f�girE]캺��W�W�GP@^::�=X	I�0j��)Vr�heE�{y�,Xi���W�R��C��qI��4�c7-���
nIjc�>r]��ѬY�ͪRN�����6��w<��Ǵ�.�W`A�\��k�r�mD��H�p�wsϞ+AÀ^e��yk�x��i��m;l�����\Ŋ��P��&��ܴԹ�e��-��X
cU�w�f��l^�g�u������G*;Ul�Z��Fs�����(L��@�I���_C��ٱ���(��
���w���'�,��rE�S8�:<���J���د�D���qD���S�Dc<y������>�X�Lh�Ѧ�s�p,J�{M�<i͸�o�6���n�ٗK��^U�yؕ��Z:�$���j�ٹ�Ry�[N�R��{)�N�,`(l�l�z�ݗ�<��n_R*ĭ��'ٙ�n�h2����E�c}n�1WS!�M�.�칉D�ͩÐ)�5�ɶ���P�w/��q�6�5b�8��թ�]���o�9������a���`0�r��9�T%�6����G=γ�s�K����Msܬ	r��%�m[9���qmI�+��c��]�{e�o�(�Ƹe����;8��e�]n�'Vf.X�gmܔ*�t�3�=H�%���C���}�#Z����̨��v�:D�S�|v�_�E7AC����������'�^��<�uZX.Z�碷t�`��f����y���45&_S[,!Q�y�-�%�3b����&�Cv���`}���u�=F�5z7�[��֫�,��H0b�b�޹պ��U��Jڰ��!K�/j��okc��	������ԗ=Ǎ�r�������S�o|�a4�wv5�>����Tz2r~��?}��̡� ��d�u�ߔ��#.��n����|퉛2Yٻ;�Kp[�j�Mu�؎U��'�b�5�{���\�x����re9�S�7}S��8�s�#�{R�*�7֪�L쬧W�33='3.1����ᩬ:7U�`)��i+���3���c$V��F�������1��;R?}��U;T�T�|�&��*��䲸�1y����E�P�q۴�V+�\t`�"z>���}t�?@�p������S�{
�51s�C�{��(�d�{��w��"P�\�F���_rW����<��ᝲ�I���
�Rd���4c�䙢�8�-߃��Ḟ����Vl�mÝ��:����'M���sb�O����
���A"�J�c(��E�,Q��m�-b�UL���j�j�aKUdX�,�ID[p�ʂ��R6R�j���d�Q*-�E#$EfR�P6��
�F"�~��Ve���2�Y13t�
+]�c�%�d���XZL��{�3�A��3�kl��1_u���q#(nX;�f��:� �z'�.e�т��q���`f)�l�p`�;�"�o�/z�uab)�QK&��i�]ԩ�<[�����S�L鯾1����t�����E�ː��U��Q/��҆���;H07�����Q��//^���~m�!�܆3��_��s�/����`�n��kIا;z�b��Og�fJBU���6Iv
��g��Zx[�+`\;���u����.�{�	�e�@���ޏD���ɀ��3G࢏�`]�s�-Z���ڲ�F�D�v]�L�u�Ny�Ne��F��C�LdO68�ϣ����P��d�x~ݘ�:�rBn�=	��Ṇ,��V�u�}���׶�sq�m�
Û4��X
K�~���x�I��{�R��{�F*h\��p��ΦLY���"xOW���~_7��� ��TAYT|�T(�W9^m�kF���/�N�"����IR	�AV��Um�65�/7lΘ���ol�1B���1RK�.�m�Si��*.Z���;�<�ct�}2f��k/~��f3� ~��F���w���x+%�l�4��,��p^r�:2b)D|Ū�V�L��}���;�8P�ЦP6�\��nu���}�Ry������J4v�|Lb��:m,�o83!Ӌwb1�u��6�HH��p�S�C�z"#Ղ�ֹD3+�1G��c	���3+&Ú�P��ۉ�����uF�a�kp�W���J59��M�a�}d7r�М���m���s�]g?	Gk�D�y�{��k�f��tk�Zo�m94�[��W���%1'�109F'���<���O/������9�Q��C���[��5J�	�����IX�i�[����5�ԁ����6�ji\1ɪ#����?�����.��ԥUu!�eib<Dz�D�����X��J�ANj�˯=������� ��ږ7]����nJ{�Z[X��&�����]k��)e���5ۈ�os�M�{z�/پ��T�]R��ɒ3��б+��s��$swL0���oY5�j�ٳ�U�[S�_�����z��ܵ�����w9���$:yi��\�T�m�
u���ݺ�w����'��0�6����s]Kp4�*�︴|e*��E�E$X���ᕐu����|�j��?)n�K�TP�3�3$ƅ��>�ڻ�}ۘ���! >��k���@�~�~����%q+ب@��\�L�2�[t�Nõ�O�̰pv�V֯Ob�
�R&FR���:�3�s��F�R��=��Ntھӹ��_Z�����ᠻ�����n�9Z��f*����DDuI}՜���.�ᶗ�\G��>��߅aON7�-9����T��O�^[W����h�#���:a`4��w�8,���:W�qW�s~Rg4�(�j��EG�'� !���_��orEQ3y\Ռ�Zn�mӽUܡGI��
��!yʆ:�� 9��ڷ�4󦲭u("��U��D-�ޘU���wC`��7k�A���<.����Br�D} j��_;��Q�{�Ԣ�OL�Q��&*!��R�!�h���ό�83���7I�:�I���x]��>AGβ�`.�S��|ɐuU&-�DWN��jS�4,��e�LP�%ʳ
c�U�i���;ͻ����oN�v5�/쓳��wN��C�����c����+��j^�Y+�F}��E\ރR�r�P��l
��L�G��`�1��p�gkǫ����Udt�#K2�OC�=[�����aF�Ox��<������-�9���=���`�:�l�]7�1<�X��h(liл:oy�.7)����k�̘�xNS�N9uH�#.��e���v������Ku�T�d8s?����G��f��~�����nK��Oj3z;�X�"  ��|�	���7O�֚ي���J���˘�jV�m�s5~��9�o'�����+�u��if�bW����fP�ۗ�7�.�%ۚ�\榓��1�q�G�#�"k}w|ïq��{����cS_|Pz�E��[&�c�6�(�#��i�=WАj�O!U-�F�\%�C�[ѿ_)�F��T�=�0�q�������UUUz��u���� $���G�5��7�����Uwb�e���r8����
�k �K,���Z��M��j����8�a��Ϣ~�DV}z-ܱ�Ǎ��IrX��EN%�̯Q@Dk�R+�\՚�ej��"�<5����Ջ}�߭��_�.���)��Q�� �Ϩ+��*�	�L�G�+nc2���X��a
�<�yr�=�z����'��Ma_e���M*��b�ܶO9�F���舍眯՞jfQ}-�x�����jHZq]��nZ6g�m_(v���?A��D=����T� 瞆G��D�Z�	m�[��H,+*@��HɅ�H��V#eV� ���+.\D������#A�	r�ff-�U���1I�y����m�N��G7��Tm ��Py:�pǹ\���,�y�>��u]�-B�K3�uڙ6����
A�ɖ{ ��W�ӵ���j�ݎ�����etDg��h���-�)|��X!m��T�s��2�ˏ�g}��k�l}���XhOj0939�6C7E�ޓpt�����4��K�O�/��*�3Qo�%o��qV�a~��l^l��xZV����[:���{Dn)~�ȶUr��N���n�	e!k��Ӛl p��'4�NQ��WHv���@t�������6�����]KF2��aV5�xu*����%H޸d��!�|��J�]9-��|��0���M��."3_e�����G�����}N)F����+�'-0�����L&dr�����[�T��=h#"8h�o��aʉ���+����n�������U�]��r#xL���X�F:� �u�6��n�"��%��/ÌG����z#�{܈$� �L*b`������9������w��S:=����f�]0������7�ijTR�Q�=�!�m�D���|pA��j�CP�טU ܝ�l�/��®=���2AND��.�R-�����Ø����nҨ�y�*wIN`�Hqs0��)ܞ�NlW��l7�]E*ܚ�{�}M5��,��v��}I�S�0;S-B��5N8*��0�,ѭ-#����ֲQ{3#����A�1�B!����Ǣ<����ڂs#��r��t�v�C±�7|M�� ,H*�qқ�8K��V�����y9/kK3[�H��'�<곴Ⱥ형����;,���@�d�<n���:��b���2s�Ŧ���-}�d��a}kN���_�v����1���Z%�ٴ.��0�x 2<%1uG]�i+�R�[�u���0B����Uy��Fz_�Z��#eS�L���i�SȦe֫���5�}��i���+R�Z�'���$�����c�m�>�\�V����G��,�ԫ����a2��v�Ȇ��4BS�8��kl]��L����(و0�MNT�e�`�o�E�t&�ˠ�-'Tl:���٨ofp��c��DY�i_�ǻ~�ϫ�s�"��f��`5
�`c�^��r�=�:[���şn���R @ �A�{���"}��a��>T^-}eҁN�����W66�tp(����p�@�L��W(��i�9L��̇�&($�W1U����w�
TK/8Ȇ�VIp5�u��J�M@��1}a�r�{�m,%� ��-���>��3�(�'o�QL��i��*	��1�����9��A��0��{��?K~�h�y+��|H/RH�&wX��؁���$	G�H�Z-�!��{��Z�� ��fu:�գlZJ�a�执�Ȼ�-1���9BlJ~��m�Vi&���f�k�0���߽�xI���{�ٳ���"�����X��T�R*�T�H%@�c �
���`�\�_��λ�iQx_s�i�����T���.�x����,ܧ���<��H��r�޿�e���^����]n��YW��^k��Ly�O�ٴkwз�})Dx�T=��u��L#=��+��A�Hs�˪��е����`C���-d���	�8��w3Ul���k~ߡu�:�L:�wi%�ו	�O �UNԵsH�9���"=5��)�ӭY�
���w7M0���X�gk��.�~$^~tFO���J�����,��L���p�:�}��(Z�Y"����S�N�kղ��im��5,f���d��=�ڹ{s�L�����T�w`�l����
~���V'���!��QՋe��ޘ�������(��8�F���^� �&�P>|�9<<�F���[�'�GU�d6$���mZ;]��� S�r��Ц�M^��Zd>�,s��3�G��b�@���[Ct�Ap7�R%����]�*L��������Z��G�7��A;;��|�������]�P#]�-'Ǳ�w�[J����aJf�ۭ�S9��
G�n��:�B��đBt�e�ՈRl��*"�W��u�m�c��Zu��h.noY��f�K5�ۭ:Tݥ�h�Y��
ٜ�r\�M��S&f�(bX"
SUd"#@�y�kS�)Z��q�0�>����5Z�F�����b� -��T�$K���(�]��w�p��V?]}�N���K�����zbf�*M��"oZ�{}�f�:�����L�N6k�]i �g]i��a��[�5w�]��)|��$��׶�X����z��NZ9\��w���˰Z����a�$H�-��XС�d�;���Yd\�AYGXLL"��P�2ULl�*�d�r�V��.e�1@����*(o���/޹җ�k����5�i�Ӛ�L]��f���l�:�X�8v���U��H�5���:��T�Ԫ�"����}��7��m�ܴ���ɳ�ֆ]+�e�`�[c�ڍ2��X�O���)��M�e�e��АhL��4�]����x��:b����鉞<���@�B� �{ݴ*�
�6�4��-1�h��L�����ss"\�B�{�IRM2ݾVn�����݁����/.Ê�WE�fa�8Hw�̛��t��D5[��@K3����Y��l���sa��0��"Ʋ��+Tkv��|'0"yb��G;y����`M�LP�\�d=��DD�f�Y��9�e�E���}��ΠmhѪ��G%]:��s��7D�[V�;7Q,[��Q�]/�p�o�'xCe�CD�b�܍���Х��Jԩ`]Mv`�h�WA��-�ViC*�ƥ�ob�@ِ���9�F^zp��B�[��ՠ3!eJ!g'˯O���#MZe����l��.E'.����ҚH�/�j+��.�\fҨ�tC0�Nk�eʹ������%�Ót�,����l�@�it����u��r�4q�a�|���RP���A6�ֺϺ�«�C��Kr�)��3�+��Vʌ#c� �8)��M��mI;a�v����*���%�ܦ�J	�	P�@y�hGCV�'qO�(���[���)�u�x��Ty�z+;A����ކ,�����mH��)U�)0��&t�������Y�ug�կ|'5��=i�ok��8էcs-"�V�����N�D��c�i��R���E��c�|]+����k/�%�X�:�;�f���X"��t	2����g�<�$�4���m��$N�w�F���
x�M�FQ+��!�|�O�w6g�v�`7z�3yݐdGu�oR�w�tNG\l��t̮î�t�$�����|P�ˆ�QCA�RC�Z96]�� R�>���G�'���V>���~���r��{ޏz6��P���qH��6�ch�H�	�pY�H�����\��K�:�޸[�㑷�-Ɏk��^�)� ���`5]�I��q���_r�+jo�dm�͢T�Q����3�si�@q��ħ�`6,�RgMu��mK��Z:a��do����eXya�aT�i`����us��ۦUU��:#ވ��)�P���)��
(<��0�Ê�8l'��@C6���əB�pF���%���ɐeKʬ�VH�<,�G���!4�Z���G�ޏb�Yj���y�Ѽ|3���K+��Z���H��(�E
Os����U�ո.��+/vY�+)����CP�3��iR�] �ܖ٦�d1PX�1B�%�41�̠T�H�`̶KbȀB+d�l��cT��eREu��"�im�GT�|�H+�~���F���t�6���6x7*K�Ǵ��q�eQ9صv�Ym�8�6ݍN��Y[�(��u�"�,n�Mu�y'/0�}܄�4{���v�mD�7�4�E�tr7*»gB�h������[���E#���?b�n�ڪ�U�p$�m�_Vr���q-���E�B&puJ]ʣB"��C��h�N��{6#��U,�����
��=�
���p3��V&8�*����Tsy��yNٰr&0�kgh�n@	͘ .��S9W# .u��z I�[܇F/��H2�*�*���Xɀ����r��t�խ�g��'�H3ZB犮���?���t���H�32zb�z;�%��V�+�Aۋ&�5��ji�R	� ���5n�Qw/�N�2�M��E��=��WB�C���|9ο.#�J�Yбw=�Ƨ�eX�����b�1-=u�O�����^�]�z<�G��H)Z�����ۿs��~7�k_u�ܤ��YZ� '�"ᝃH��X�js�4'5h�[~+c/�������L嘒�sM�6[9�"c��<;W%C�����rv^B�jϳuŪ�E"uN�r ��M�ҭ�m\�Yj=-aCH�a�j��~��w�x1���侉�h *]�ɢq���e�Dk����c����ɇke|7��zzN���7�؀{J'��NZ�-5�#�G����_E̤iT��"��_V����Ꙟ!"�� u��c�䟐��5ꉾm܍����DDCP��z/S�-��E����b~^�R�D95U֍}'�S0>��к�9=�֥�a��G{,c�3x�{�X�C`;���wge���E��cG�sdȌ�n��Z����G�މ�G[0�J���Q� '�(@rHV�p�|Ols}r;N���$��Q�-9."4G���눈���O~�����C �
�lq��f^_=�*SV�nR;W�3J�6R(g�'��{*�jT�����ܾ;K��[;W��݌Q��ʷܒ��rZ�f��ꬍ��ckjn-���B��S*r�eqY��k���ʶ�EV'�H�Z���0(H)�s
y�Lg|z��D:5�\��m������in�T!P���.�5�R��v;�FϹ�7|���l�j��\e%ͺ��튣�}�eȚ�AR\�I�0��������ӌml�3�c��LJ�aq ��SiW��x�祟r-.�_
����ޏ�7������s�p6Q�=�.�i��������h=Y-[�>=����g�2�	�:i��E�w:��2:}q����K$ۙ����G�F�@��H?d�!\����vO��{�r�`�U��MS݉�5����`�Gi�wh�[Xh�>W�`��������E���٦W���+5N�X���6�:�uTz�rGK����M��T�uҩh.I��5���F��{q��Ƿ�ٗ���3?^|�,є���@� ���)eL����w���s�}�ь-`)�)�j��Vsm����텘�����.���#�okK�j�����2c<s�}��i�U��K3�夑J�'�1�A��i�jP�[==)Xc��FJY��T��Q�Q2(�P��oUX�������W7q��6��N�K�8��nv��<�@
:���^� �VY�Zw�<��(��,5�DDD���j��_E��z����s�/�/�P���O*
���4�5O�F�vJ���C'�L��'yvj�����Ҵ��]�]�B:���j�֚�ÿ���1(��@Ǝ5&�@�.�{n����2��S8n�ӱ/���M�y�d��z!ܙ���H�ۮ�n�\Lr�cK[9�Wm�tj�G$�l���X��%�x��5&{}��r�NEk��SK�}�ɲ���p:+�Zj�Ժ�	3ޱ�حRM��嘝Nw�9��T{k�)�,+,T�b�BEP��1P-���N��߿_޺�w��j�[��E�Z2�r'Uz�(��9��yD����-kQ��Y �.�%�V��S������7���;Jyw�]�#Ow&��^~���`9V~?��G�"� ��2�5�-t��3�za�m�c�e�"�f�2��}�YT.GmǢ��pӫ��ޝ#-�]S���7mL>g�FѨ�1;Wl������	EԊς�Cg�5��{N������@E]7�O��xH���Ā��cb�%ʋ�^i{�F��s�k�mOY���+k;=�naV��>t��](n���o�%�>�'3�Ω�B��	��`���%�D��m̤��ON���{�	��YT�!�aѱ�{D���zġ��:�k������8�k;|��[�w0_\c�;X�φ/�ч�@�m١Ȩ��}�+����CZ���z#�s�i�X�yԃd��}3�@�%�2"Q�C����` �� �Da U�1�I%��EH(*�_ @�������rmo���J�qWc��6��9p �^�hnr�B�eΊ�!)��_4Gt�.[n����W��\��2��tܽ���]:>@�3��Y�/_��i�4�$S�鱈tfh��_o�@:K�}�Ջm͞�4�E���W8��кu\tv�Nܱ����#��
�*�����F��!���l�1��s�]˪���=�����Q�&2���t�
tDf���Y�+ѥA=Y8��ӲG])gL^�Q�����T"Հ�IWl`a�'���뼶�{6t��)���A�_��5���!J�=��a`ɠ��bs�DD{�Kn������3U0�������#^y�K��"���>x���K�p�i�nLeÜ%J��IL��NR{������=M�ۋ�����q��n�Ge�Q�
��ݧ��&�f^�0 Za�A򜝩�ɸ�<��dfu��!�v��j0
S��2��{yBԱ!JU�=������]^w�(��W�Ԅ%oD+N�t^- @��ǯGh�ލ����k���2�1�sF�)\�G&��9��f5N)�&�h� ���������積� +���	���5N�S�}�Ec��K+���Gϳޏx���Q,���I��P�DD(kiB�*���䓪s�;�{wR�F�����)�	D�(���J��m�L	б��0�Z��{��6*)[�^;�(�4U��vr���:i����4/�,�δ,�a��*p���:	�zgjr��jO�p�g0a�`5��l��R��>�D$c���dy�)��.rfa�o�<Oz���M#:߂;���/���G�=����ת�����}Y���F���x�7س� ��̔I
�=��	ʭ�����.�O:������DU�k����rt�l���$�\{��d�U�p�w����G�����Sb3�׋�Bɾٱ�:�j�<6@�1#ߐ�4�V*�#&��B+[~���6��C�!gl��yR
̕j��%l�5��
9��֚�l�u
�sd�^��e��f��y�%��Z�A1�����T~C4�VR�j�0g�d�j�[�<�'��R\��}���8�Ɗ�0ԙ�v��$!�~��_�֨��Ղq�Gn�to8�5Ӵc�^��r�C��d:�#��B�.����AFO)��Wv�E�ǩ�5�둻�B��!�����$<�G��M�O*��!��U�೽N��$`���iM[� ��N�ջ��:��QD�2i�(C��8A�Ѹj��)��N2�t1�4�N��u������4$V�;ڷ����J������Q�On�D�Af��r�@����u'o��;���H{*:��0 9;0��K��J�ܳ����Ɣ��{�=�
��*}�G�Y+��"l2A��gG�F��7l���$� (�"Ȥ�O�%�}V���߮�"0;b>Goq&2#X�M�b��}f�P�ϛ��o��oT�oTe�v1_k������ث]�-�a�`7X��c �}��&U�k���>����s0b+Jp�Ͻ�gP�0[��:ض�0]"=۴��
���$;)��ݾ
�M���0�H�)�N@�Z�ڛ��bw"""���N֣�٩i�3q{�Z��3�3��y�.N�D�ӂ�C@\��Ɖ�txV���<�������f��L��H�'����.[K�,h>q�k��ͦx�x*�+D��zUk�)���D7��Y]q��e����4V�嚁!Q���y�Gl2�C�'TYS��U*E� 򝧒��0]Kgg��f�r�u�}w�z�P_�]Á�5^��xG���A57�鲐����V�BYgCJɥX8=̕O_�>�h����9�}����]�@$I?� �	$�� �	$��@$��$I?� I��	 �O�@$I?� I��$�� �	$���I'� $I?@$I,@$��@$��@$I?� I��	 �O� H���I'��H�v I���e5�B�� V!�� �r 	 r}�![��B��`A%IKFR)@T#MY�h�IR  �$R� F�ERQHR*m��͠PE
 E�EDJUU   $J ��$�)TD�JEUJ�R�EPP��
TR�*J�% ����	�}1UQJ�PTD�\��J �6ҧ3F�DF��h�*S�e`f�,�m��=���S�j��9�]wuAT�����wb��]h.͠�m���JH��TQ�Cg���nwz�`繺�9�]y�� ����.�3��+�+��Q/{�����{ޜ�;�wYm]ܧu���-a5r��m��2b�ZҩW8�Q��]wcՇ�
�UB�R(�IU%Rw�n�;m'UD��M-���\�om���v��WZ��[�y^ѣZ=Q���A���v�r�����{���5Zk�W@^���-A���U��5n�R�@�J)TAZ��0��T�N���j�I�NXf:���UZj�;{=3��޵6�A&��:��\���oK�1�UZ��S�v���su�=�U�v�������䠈F�J�D�����\�����m�KMt�ۮ����/:i�뺽)�y�^�G�]�!�ow�\�E��v��t֕����3�g�(r��7�w[����{��ke�xJR)"�T����Hp���{��X�M=��7����[{�xuޞ��V��t�۰������t2Ѫ�ފ�Z��t{���S��w����n��;����k�=����Y������PT�HUAH�"G������n�Z���{�.��z��ӽ��z�U�ծ�������:2��5rݷj���W*�i����Vn�^�.�m����y���^��r�����\7e]�J��� $��@��\�Ζ�6���6����Kj��V�Q���{��*�����vӜ3Ol�W�Uy؋\zz��v����U�{N�wn���O+�oN®����˻�u��u���Ki���n����W8����@��P��r�{i�v��u���6�5��\�[گ{�{��⽷��ou�����u�v۫�[��/]ֳ����Ny/n=�\��ojq^�n��mzk�:�{z�����=m�M�ם�]�s:�D)I
��UJ��U����Ӭ��z����2�n=�/W�{۽�v��pz�������v����{ vԹU��ztt x� ��< @ �� ѣ@7�      "�ɢf�U@ � ?h�IJU10L*=O'�h   T�T�d0&� �{F��J�� 4  � 	I	Oj��4ѦO$�7[4r���hDj��bC}�5�@ 	dl ��2�DUk�p��;�	� �3ff5�����3ff�� ��}٘`��߆0ffd���f���S�333��0ffo��337����!��F�>�d�5`р?3.._i�d5%���٭$X"92S0CI��5�qD9�0��Y��8`$fh��0���QJ�4��Tw{�g_%�s�����I�1v͝م
)��K�eݳ����Mm&æU��g@\�����:u��ݷKh��27Wq7���s(]+�4���z�΄�E�%p{�1e�t���`D��N�6j�=�!��.��tv�*�J��M%,�h�IH�Z�R hk3\I#L�Հ�h�b�ڔ�*��@�3%�����k�%��u&Aek:ÖEm�ӏBմo[��:1����N��ߔ2�yo�T2���#S��O/��Ƿm9u2�gh�΍��}ڕ��vθҽ�qG�M;T�ڳ����"�$�Y�����0r�a�`$���Y� 60� ��(�C,�K�0%��2��L���:[��Tn�����Vz�;�S�p\.����ik�z{4�]�j��0�n�>����;�1L�'m廷���e���+wh���P�VK�Iv��؁ҺݙYp��L2��RLw#�um���]�+:���@۵��]i�ju�8�<����{jı[˼�閃+w:���*��P~}�f�R���pY=hdjvn�]&b�m�;9v
y�,��
�Weȥ�����nS�n`#MQ��L
7J��y�U�onS�	�U(*�����6fNU���iu��4�9vv��p���Q�qm$�0� X�r���h��&�bۭ�A���r����aL�qv�Ƭ���s��Y{���a� �ᗅh��G��jb��w7H��!2��gUnS�ڥ4�g�I�0c˭�����ud#g"m`ι	��#oX<��Dc4m����r0N�zf�U���R���uv�7��2�� B3����-�4�V�c���O1*��M�m�*�i�p��)C+4�P����@����J�EZ��/aҭ�Ÿ(�,��bǣbx.<��M��	�P%��Cј֛7�i���9*�GL���t˵H3����t��2nU�V�׎D(<'�׋�~k99v��ޠ E�p�ZD��aSsWt"`���o7B���I�����LdSt"�kqU���R�����席j��j��U�c�a�&B���	=,�d�[�c҃`Ё�2�!K�4��"��E-�h(�%Vʵn�Z'�z���p�:���Nn�5�{q-����8%���HEwWx57Sw#z‵&XP��i�P~�^T����Ԏ�Q%���*�\�R�N���QX�w���hT�
�v(�F��b�Yu��E�C)7b����&����<=��� ����;z�*a`$v��j��"��S(J��bm�y�����@m�F���]�Tf-��W��V�� �܁�m̴#t1��n������m�Z�`�ՈS�K������.j��Ǉr���j���kD5�XT���y�T݁(��*�F��t��F�Iou!J�dշ{.=�� ���or�2��%Bռ�)U�3q ��`����Jm��P�	���Wm,ۭ�M�qf��8\ڋ.<N3Vm���{-Rڅ�ff����S�ՕI��YʷgY�)+�B�670P.�P�x����A�b��,�1GX[�(г ���%����m��lv��%Ct�W)��ʚE�*Y��Lyv�4�X�=d�bmmMǨ��{�ֶ�Zơ���xh�6�Á-9��q�,�%��-*̷�3��j�j���ٴ�;v%�4��t�j��L��`��N��2��Sd�ZM
1��g
���l8�a�˸�g��5vֲ�PŤ<N�VPM�+m�@���<�9K(f�$T��c6���ю�cҨD��!�� WD`��35y4�F �;5����.�@��Vv�N<�� +�P̈́0�Y$�,*��V��D��p�e\��h��ƚ)GZ-R���邋ֵ�ٶ0���4��ۙY�4��Q�r��U��ZK QA�cj[2$���$��FbBe������Գ��K+K�d(���d�@�
��IV�j�Z�a���Fݱy��n;��iլ,��A��^m#%��5���ki]�#a���M�:�F&�� ���e��.򒭓Q�?,f��J�2���5�qñl;��ұ�խҲm*�lB�R���41����@*س[�� ��j���mA*G� �աշK�m#E���4-��Le� Ml���!��1����dL�C[�˺Mf�~!Uǌ�pYƛP�����NԨX�pT�-��wn$�dD�6Tw��oI	�ɕ��o�%���x^$`JՋ7�s`̫�b��uE +1#c���F�&=:(�)�ޓ��d��y�EP:�%�̾���i�����vl��Su�;�3j6j����ӽP�oP��+R���^�:�)f\ji5v��f́
�ܑS��@[.�DT�E��a�I��5k&��X�C�����m&�[��<�� x�Jx�����;��̦Џnܘ`p]���9�Ka��X��⛳D��s��l[k3Ǯ-�v9�� $�����3Z�&�f�lB��9Q�Ym���@�I=�ZD�f���`EH�(J�.ZJ�V/�2�b'W2��3*���J�9B�ࡈ��Ȥksr�����Z���=�^�AT��%��LH�ۚqҹ��?������d�f�Y��������ꅘF�Y��C,���a
2Z� 2����9�3Lӆ@4�Ds5��02-1���r�Ub}Ï{�T;�Ǳ���HR���ރ5z�e�
V��h���@:ݤV�MЙ�D�B����^lZh@�ghS%�/x�7��r�5�|���QV-��z`�S��f0E�}�["P��w�b©iP�Yk-*������le�B��.�O�s�Y�[��w%5աp��5�U�W�0�{�nG]�3Fer�RX�n�{�.��y2���zkks�I�.񗒢�1~H!P	�Bw)��m�u4]u�	9�D���C�,���.?ʮ�f�l�����[X�g]�j�q�ŝy�Wm`wP�%���X�V�Xʗ��; ��P7����mf��3��!��@��B����S6�fVʓ)n5W��_��gNب�"�U9Dvȋ����i
��!�d��!h�2�o]fVVb��� �c��1��ؙ�a�g��+M�<�AM�	�)�Ŗڲ�o/^��4;�%(^�#hѧ��熋o� f����ݨ"�7bܥ�� �� �V�ص��^= K���6�x�%�-��BZ�F�Ի2�o2s*�Ʃ�Ń[�i65Ge<�0�@�Z�Ň�yI)�Îf�7l3���e,���F322a��H2.�XZü Дc{E� 5c��ѝ�ί�6�	�̻�N�J;u��P��&�_��q�ُX�s�H�u	�l��T��,&Ү��.6ú��ۆ�Aan�e���L�E<�T�����8X����s���I=@i
Q7�~;�SV,�d�+���X���I�r��9�a�,SͻC^][���ཀྵ/��-"`fQ�i�!��n�\)�j��ī8�m�L��t^
]Wek9��U.�9)�1����ݻ�k1\I����9��y[�l̻X�S0�y��TT�SA�,��i��D4���ý,fX�2�K\U+��w]?(����n]�*�9n�'oZ]ۊ&m�0mB� �W�������Z�a��6���k6��Q�6��8*"sBwi]1�D�¯Kn�8�.�F����o�1�qH�lm��~�)Y�NSZ���{[r��#N�ͲG�LG�:= �pι�^�č����Ve�+3�X�w1X��!Z��d�%�e#{,?HZ�n�*����oȷ�&�1a!![�u����f�I1W[&�N5D2�+�K���t��1�Ѭ� ��RY���i,�}�Dwk�"��6�Q��Y��:��4�Z4�-����ڛ:CĲ��^�����d���p����Uk�
[�=�(���MLtw&��[��nV�32��N���Y�d��j�%H[*ZBzjKt���m`FbO+ug�wGt�4�x"���%�䲇�	K�hG����s��Gk7�dԴ���J�[!o2ƛ�L8��.�P���usL�c����1�זt�
r��ױJ��n�6��XrU��Lݕ���h^JX�ǏK;��{��"x>��zp�+%�0˼�T�Q�s�6���جH��MLq�H�x9RxC��!��b"�.V�I86��=˨5Y�n�h��F��/v<�6X��>4Aá����7FC�җl��A*���������f[긜Zt�{]��/:�s20	C��MJt�Bb7�5v�� �����(5d��(Q�Z+3K�.�@��l���m�f�	%��363[��B���I��ۂΥ���-�t��qG�ޭ�3î<�.�ZV҅+7��ʻ���GPެ�IEkktK����ą�^��7v�+b���b�[
Yt�3F淪�nf-&H�P�Df�9 a����1Y���|�����\���cF�*ɀ7�3��f�a v�6���T&�<�5����aoz�w�nROJ,F��?�^�f��Eڠ���H
=o��5-�*���e�pZ��J;a��䦘V0��唿Yl63t]Dr$���#�T�5z��Vٹ�ࡼIow�dv_�$Nܣ���k��6�v�e�n�h-SSZ��*@�]zm��id�d*)��a���nD"v�[ԁ?�����khJG��@+/ ��;��XR���/��ׂb�%���y`�QL�P" 4ܳZX��D��v�W#B͠0E�w�mݗ|�45��f*yB�*�op9F�1.�zEiJMA��X��N�U�u��Q��h̨�����h���۱��%A1��T[��Q���W,���RW��2���U�(jr���rӵz�j��q�g%��[*e4 Z`	��!�Y�κN ;X�P�1�����U�#T�bXT�O,�\i,����'��2 �x��e���ia�-H�w�F���Q��N�6�dn��3w�p��m=��
V��Ԕ�f�F�]"�u��M��xC���9;�K��fm��2#�6OFuɡ-��b����\��#]�-	*�l+�So7��a�\��<�c�ϔP�ݷ9R�iׯ52BӋ2wV�����Rf�-����%� ���I�z�8z�/�an��f����X������9Y4'���kY�J��|�
�+_�]���[.�i�s8l��S醭RT���3SV���$�Nk�������Ѫ��9oi�1�^�{d�^���ERf%մ�,���N�p�DO��֪vQ#y�Y�g���Tb̾��k0w���.q�]EA�Bu]������JM�BJ�-�i� �ct��(�i�?+{#�{u���l���a��T�8��"��V�IS�.���
�D��*��H=�/zMЭ�,������a�b*:D�B
�}�75e3�J'#��2�D�����	;P.��sf�WW��WJQ�"��\�J�C�� ��S�5�n�q�+l;���e�Bd�t��M��ę�-���4qi�z��Xуi �F������jC#a�[���{,�Vr�"F���*\���_����[J�2�"�*�M�:���	��vY
�=��r�F@K��X�n��V3�"��7n�cpE��f�䱺 ����S�L���d�nB4sPb�&���U�R�o��e��jUӬ���Vat-�y4T����_��L8�$)A���v��Rz�7�o�e՜cj��[��fT���p�Xa���{��m���ڰ�L����Xݍ�ά��j�&��ѭ���&M����%�޼�'�8TBiʻ�e
bR�{=j�̊�[W�kE���0�T�^R#	sp����k�Az��c�I^�o�%�]�vl�N�e�i��im:q6�`ׇ3���3j$2����m�����;ե�D8B�K:֜FL.�f\��M�q�,��5o�ғOn-��I�#on3p���no�q��L����բn�hX3�*,5��2����i���%h��X�2j���$(�z�$T[Cm�N�&�Lݗ�C-��K%���ZN��/���M���,Ihm�z&m�l~��tЙ�f�� *��kpи�hTeo<�QXа4���V��}��P�C\[��UDP������u*B#t�vbw�{x���kb�v��Ɉ���Y�3%�-\��
Y�F�L�y�P�2i!�Ҕ�J�.ۭo{H�l7Qj�W�\ʂ±��vBêi�ȵ�k4���R;�j����-���V����Mnc����5�ۣ�b��cX�J����[2�����El�*�ڷ3h�6X�Gj�j�#/��V��t���7����66�e�i�R-���j6Y�"[���z�w��N�;S�*QJe�
e���7�F��75b�q,�z�:Q��h����m�x0D��˽�����fn,�b�N��ƍ�I�V���x����~��E7$��ҁL�Z�aw[i����4���*�ŭ���Z�bXЇ#���0y�$Ď:utn�uk�j�~Y0�4P@ +0�5�V<m���?l�ڻ��F����R�U�ko!���NVvR��Ŗ�	X���Ż�� ���-�ӭUo2T���Ȏ�~�D% ,M��,U㻼�
z�wv��vV� )�yD˦t^#2�V躳��?F�#�6d"d	*ټ1Z�,���}��uA���4��]#B3.ȩ�/G�c�Y��� �^�	�<S{����M�K��_�dy͢2陜� |�x�hٺ�ƣ�u39ζ����7���v���W�v+�dR�c����*�zԱ�]uG%�In%8j�F��X�Z��:e�T����}�^)&t�y���7zO/-���e�qI8JqIH$�S�:�UZݗ��v^!|p����ݏX.z�m�^<�:7$o����7�F�H�I�$}$�N��$���7�H�I�#}$o����7�F�H�I�$}$������I'I#�$o������7�H�I�#}$o����7�F��7�y�I#��wr\z�.L�bK�K�N���%K�����h��8Q��Κ�4�r�9���r��kt�S]�j�4�_(�H�U�Ӯ�Ww9W\���XD�wuI'Jl��ݥ�'''�wt��9�Wws�qk��[���{����*7�Q�Iv[�sMr)ӝ�4�>��+�.�#Ir�m:����E�Ҙې�D����籽�!����2to������GѴ����j�s9(ҏ�m)�x�t�^vbK�&nG͖�[�Im�ϥ��ǹ�$o���$'��rIѽ�{V=�΍��j$���us��}N�s�}ʹo;wu\�u �l�����-oH4-f��̱�&ɯz�&�Z݌�&L���3�yZ:����Ҽ��`��+ZM�v�����cFNWN�S�ɽ���縐>���z���4G�7{���ѱq
�����bQ
��N�R��X|��ؑ��3�ѳ�\�v�b��Q�s��J�2Ѿ|��;;*&�U����ͬ��]^���h��j�-k�қ�ϭ�x�7�VK��v1.��ʙD�B^|�%^����f��
�|�.�̪�ქ�\�:D�^	�N���M�(�e��h��O�6�����y�t�C�8����2b���wG�t� UJ�]2����ukV�^����vBlk##�|��.�
�Rot��6�%+3��%m'ҶX���յ	��bX�T̻]�+/�]zks�B�(Tu-��z�v�����J�q��ݓ/�j�մ��J��b�H��m�T�<���Y�&��]n�B��4w��Ӆ{��H~}P��7[�t"fY��J��92�����7r�ɱ���s�;�u�֞�ʎ��ުYA�w�4�a#�t|z�@UZ�3($�^덢��8������P,���.w��y���7��hv���`���l����,�6�!FV­v�ß;�}6�<����S]�y��_�oŴK\W�3b���'��6�jnr��y�m�g�|5���9��RW2��T�WB�6����U�R��I��f��+ݒڬ05W���h�5��U6�Y��^�g�MɰՇ���@Iedhs�����c�K�;'�E̳oYم~�UQޮ�{��K�l��:h�wۜLcv��������xl�%�,�$sѦWnP�y|a��'��*��43����mb#oi+u��ԫ�'`��]����)��*��>��;�{�׈��j�\���z�Ҥ��k��iXUί�,�q�!�S���0�y
���w��	�V�=؉��k�Q�(ss�'��ee�����V����݉��`ja"��	�W5��d7@�.k�0_5�f�ܲC���5pX��:x�b��t��kf�ua��TtTL��E�v�[����{n�Qt����vF.^��N�ch$��,�8V���S�z&��f=��)K��`��#֐\̙�G��8i�ʒ��4V���4�pB�d;�[� �{{�.S�h��Z����\�����w�3m�7ې��8Z8�yq�-7�U�3�b�2r3:�,����e�q�ζ֚s���G1�����K� �Kp�n��Mw3![IT�1���;����L�Qc��ci�.�A��_�z}坚4�SYe1c|�k�BoR�@�����;��)�0we� ڮ���nQd����!��k3d�U����f�K0z�T�i�4����e/*�(o�lޫ/�S'��D��(@���W���:ZEeǬcgZ7�4�W1� %�FoH��u@�-��V�ܪ��`�>=���Z��o/8��^)�~uhdf���ֳ��Y�T,���{��c+cq�u�Q��{rIl��W�Rҫ{
��C�,xI�\d*�X��2��y�Rj)	S����{:Ғ�uu_+"��*Q�v�K��oo��ŇÓ��s��{�,����*�WRK�5Rk9�V�A�/��`+�����{�uJވ��wws��:ʧ��N���zg�N�|7x��ۤl��7��tW��	b�o��{YPlw��Av#�t".4��/5��ke��Rɼ!�ѭX�<��۲�c��3���wE@hڲ�j�-��C	�87ˮ���Ko�A��KY�}���X}]��u;��Z�tR:�Dp^��jM]e��k��}�.�3z����ņ�X&ڱ-tU�-Ώۇ�]�6����=$K\�o�Z)�)�ƍ�er�a:�����bB�81�7:�6	noe���`]���fw�Ү���6��v�w����R�Wh ��:�L"�7�>sH���\;�u5M��֕I�x6����K!(��ҦiU��g��؂�N�v��oiu��3HV��t-Ž�q%Ŭ�+r��O^K�r�WwW:�ہF�1�T�͉�7��GfC�]mMn��v��GFY,�IWmX�$<8K��R-���켘sr�_5��o�����7��C���a}�����t5dܴj��j���d��vau�#ǒ��pL�,̣5�����]#��'r t��f��kC���c��''V�l�����]�g�D��8�E1�>��y�#ٗ9�X�^%��k��Cv��g�sO��цT��$��gj���eln��1.O''u%������v�ӫ���[�A�qѳ�����WV�wImf�V��W��e��*�����Dڿ�YC'��)���w}g:^�7Y������w凯��[0vڮ#z�vIP6�uZ�E�<�-���6�W-.��x&�[m.J���Y�z���G>��\ǃ/!�Ç�x�h<��/ygf3�6X��Wj�d�tjT�����z�n�_�C؟V��+k�p�ӥB��x��fT|Mπֳ�Y2��6?=�I�δ��g�)y0�x�!�V�N�u�6+tr�ۇ�>�ݛ����h6�qpb=�c�k��K]�#�p)���oK����=�k!g8Ų�eb6��ݮ�Kr�%���"�9�,��2��Y���R��; ����2�[
n�wYk4-e�����/6G�w��e`�����̮ǡ����O�a2aC��lqu �N{��/6��2��$͝�X�el}���N����`M�#�]��$� &LWΣ��-_�-���#r����C7�_�#���:�y�:T���.�w�W����Z�($�ix����`�uݽd�p��� Bw<��n,���M7\�w�2�Z"#j�fg7�ʾć�f�V�+������ƭ�_���Y�\:���$|�N��n(I�P],�;�xL�sĽ�god�3����L�-�Vb�^�}�O<����ݸA���`
!��'���Zw�`�]�Q�����o�}Պ����B�d�q֗"��*�,,�VTYJQ�/�x�]�ene���8o���΀Υty.	�M5��^��*��囸lCPi"�tI�޵C�:�Mɶ���e<w�j:<��E͎�q��]�n���A���K9F+�Mak�3o��-oU���NS��ҡ�s9�[I��na]�6�XH�o��WS�F���-&!plC�bǷ}��f��&��t�հs�c܉mT��	�3'B�cb���,g���o����q�Ø^�5�u���<��%�B��XEJ���(Ջ�2�q������w8�Qv��<˹|h���&�U�͝�F�8?�%o4l��i���	����܁-JA̵��=ܣ܅�N�p�fP�2m(;G�q�%ŝs-�.�q�-0�[��9B���� R��\M"c<:�}՛1�il��A�[gr�I�m����B���9�?�t��`��s�=ͬ��Zx�.+d�t;�|�n�8fܱ��7R�A�U��`{����n�ԓv��ݯ�
�o�,�7�-ljSw���I�A7l��O�꧍RJ�I]���g[{Ղ]�k(�c�p�)u��^$jăZ򝔣�j�5xGT�G�sv���Q��	���ɲ���Q��q�sS��QBww#�n�+3�
��ol�49̗���9����ë1�7����T�%�c��ef"��#��j}�{{F���Ψ�m*[i`�wS���[�b$ɑ�o:��P�0�������A�������g�8����p7�aN�V��Q��ϸ���:N����u�hpVyuс�2wh��,�[���f�r�kN2d��y���8Q�M_^k�}�bo1���P�j�'m����nU(�]v�C�u�r-}�4 lYCK'{$�`k���x�Z.�Vd�x]lu�]�Ci.b�����V�}z�*�2�|Ry:+k�c�{]+'+��$Bk(f3Z3 �jfS��1��9���7Ô@��lU'U����k��?ڑs1�<�:4���I��K&��ݗ���v*�k`�$���)M�{Q+0I�y��������>ڙxAVn٨�',�f�)s�`��Mhe�D�3���v:c^ԣ0���>y�aI��&7�ԟ?�jl�ܢ��wQ��]�fu-��h�'�%\&�2Ď�Q���G'�:�eD�%p��`Zg����Gã�Η�7Y��,�M�`г'M���u�gfr�͡�UG"�����(pFl�8��^ Ym����]�Y�cH�,8ӽ����+;�;6v^엗ƇN=u|ri�l�Xr4��v��r `���ҿl{�T� �N��ަu��{�9r��JS"���t,-'R�+v��7�Kz�M]�NR�9R5��)�l�jջH91JT�`����d� v� J�bņRæ��{�m`�U�{2Q���1��E���H"8��4�����4�9Y�$�Zl�@v�=�77�=RB�u%���̸�/ٜ����Ֆ� j���^�G��1#F�[�'��K�ҳ����*�_0�<Ue�Fbl��er�܋娯��^g �����]�^�{& ��t��cN�87��X�z�`ikw{XS��:;DX�pd��ވ������� |�:�ل�a�G]��9���:�� ;O)�N5ƈq�|�;���υ�7"d��6�.�w��=w+Vr��us�|�+M�k�I�:U򠲬�mV���tp�jP@=�Φ�����{8���sI.�yu�v�����|8��ݹإ���!0��)3EɃ�J���[���z�J�ؘ�"ɭ�w���C[���y�
AZ�o����5�صG��$�������^����d����e�pW^5�u�SjK��]�PR�v�L���˰��>���}Ƶ(�n��r\�n��*�e�<,��rj��ǧ���(�O�k�[���7Wjӯ{qej��+0���]�Y\붗��յ}�G�E*Ŷ6M�X�up�P�J���cӇ�8$��3�`lݭj��
��rز�#������̱܉ �|Z��a�-#W[�/�gs�������6A�z+��f֐[-�"�#���η#�ɱL9�V�jݫ�&��ZY�ܠ���ea7/l�v�&��Wi�jP�]�������6i��h�H:��g<��6(k�0��5I:������o���������27�1.�Iv�XnaO�*Vγ(X��֫�FV[�誹0�q,:AԿ!��p���(̝�c���ӡ[����+:��K�����$.���ZQ`�Z̺����Z���:�`fyVw��v.qX὆@p��"�x�3�/��V{��'�S:�gS�-ӱR�NK�S�ʈ�Y��i�*��N�:F�.2r�pu�9��'�����p���<�-Z7�:������t�X�2�x��^�mT���¯��y|xt���8u�Wl��ǹl���u�u�e�.޺ȓ�&�������O+k�Dz�
��w��%b��N/=�[׃�:u�Z{�RƸ��߀������������{���A���m=�h"�P ��(s�w�!�B[��v�o�*�r�H��8	�h��{r�V�i,�Zl�<ą0ӽ�4�+<������:�Z���F<@,Y�9�\��Z���B��l�sxpt�N��V�
��¹jz�R��w_td��)��_�y�:2��F)gA�0䖺�/0g0�ʘm�'m���β�'�L�+ev�z.�e�}5f�[�]F�g	�z���1�fY�j(Q��ڸ���':}!-6+.P�Z�d�:��gQ3�DQ��u|e}�y�QN[R�9�)_q�X+�˧�9�=�s�Iq�(�`kc[���s�k��SU������h����:#]
T^��:ﲂK`�w)v�k�æ�Q�S-<�r�bX�Cx�vR��K?c��h���MYz�R�t����^���5j􋎳��C�4��yrG2�㡆e�t�#��O���׉��e�h�CM�`�̱1��B�"u%P=p)}�M��qV�2�<�9�cvש�՛Sp��Y��:�w署�i#��E�6vr/]��Kd�p��ej�\��5O6^����oX�Ṿ��P}ߛ`[��r��t��]��kxOA�[Y�^c�aCB�j.���;ݔ�뭹v�~�U�K�J����3��*ކ���i�LS��;��v��R�����B��2��-	wè]��H#���4i��=��L���%�v�H�(�Α��m��5x�K*_H��K9��{w9ܻ�E�{E��Ζe�I�XT����Ƨ.[�������݌���N�.�J*��^�;�Y��CJR���Y��u��4��>�L���HN�;7:k4-�7:+��A�ꛀF�9�
��Fu���H��XU2�ҵ�Q�Ǔ�45Ek��-<Lo��c����`��e�`�_��otwd�����b�U�w]h��oc�`b��u�v�J��٥��4Q)� �@r�YM*C׬C+��E�{l���k�Q��˛7�p'��89��M�{yӬ����'T�U�=*5=XZ�5gv�4��G��6��8�Fl*V����n�E���w��\�S��N
�| ��H�
�+���Xr.ਫ਼"ɂ�Cn�1����xb�Xr�]`COnl�wmcG��{6�2u�j������B�r�'�ƍ٣��0�0ffo�����`�`���f����&�� ���F�D����$䍷�\tw@���GO����M*�6GN<�̏u`��n^2&�]��$�];]��b�Z�;�:�R~y:�^�m�,��%H��c�kI��@X�mΥ|�C׺4	3]�r/փ��ZC��=������]R��f:�J�iw"�;�����.*Q��]j���;x����7+Tf�I��5G3q޷���G�t\���u�j����\�u�i�q��� �/UNfӬQ=X-�C|��l���qb�{�w�J'i��;���be1�=|/��'u'����6ʌ����u�,�*�ڟ�A�+���{�v��}E��u��_��F&�du�\�#K!Lr��jdU�8L�帯v�v�pW;�gy��C�2��|rٳ��*6�Svm�C��-����עP�{NNk�@@��!�h8/���H�ˬ{2�*�t�C���<�]�MsM�B�
)�1g�`{Zu��.�g��
��V�W	�kNpv�E^�<�+��6H���9V�f^�.ʄ1��$���wc�r��`Sܘ����̒��\l��lM�LΌ��gf�Υ:i���ʳs�"]s5�jt�	�'�I������N��	���ZSz�D����'�ۯ�NˑnG��G%��Q�;S��Ϝc�u�um�][/�!�VS�eP�:<�v��y�ލh�Y�=]U��&(��0`�70�}�e����^��jh��n�.�	��4��b�:Rs��N�Mq�o�c�$q�d|t��Vp|F�v��9��V���;�K ,��ӝ���[�Ԯ�l�=��C"�����q�����<�������Ye{�[�h+e����o����*��@=��v��9��%{��<�
�hH��:+Ee��|����S�>tn<�7^Jղ�+]���F���,�w���R�{b��-��V
�̱�xb�/��'�U�[����� �
�qfc�{��K���_:��=QD��j��:���Z�|F��_��AC{(^�R���g�ꕇ����^�xC�+��lZ���zr�����NN-�	��^�����sL���+�Hn1�߅���\ �����IT'qEOw_����1�	�N{�Ѕ��<[�o��Vf�5���֣��%�=L�ٹ&[��W��=�׾��Z���(���^��M�{8�8��>��r��E�V| E�J��H�&�XNY�}����%�+�[�l����LZ��������%��F�Z��:��?��c.�k0�t��$�W0�|r�X��Gk�&�`C��Ԣ;���s:��ҫ�6�Z��S5���,;%M�8�:��a���N��7y{A�O�ޮ����2�_���T�������ҳq��~�y�T=�Bꙧ8�C�<Z3i?iZ[�+�����E�3�4em7w�-gʺ�w��Z�"aػ-��N+���H]�4&�!�]�����H[�z��/;��J6����X�X�V�X%I]ك�v3$$��.�-'��J�*?	���F<ǽ�˗��f����DZ�Xj���z�0��[vrÙ��}��;iX5+�M�P� �ph؇���r��1^��X]�/��N*�{�97��R;�0yO�dqx�=37�eq5�#��t:��u�C}�O:�G_	vE�R���m������L�֛9���.�r�P������q��\�s�r�<M��������K�s=�Bm�V�<y��;�F�9k�T���]mK[aX�$��9*Fq�J��{�qy��܎p���m�քx.��Ǹ>�-�`���g�|ZS�xi
7�ʹV,��ch+����5B�X���X�� �;�dv�KY/�EZ�X������%��vo�+�u���8�W�2=��>���r\7��2xpZ��)�7�+�}0lh�GӚ���٦��+���_���؜��y��P�\7#4sM��ɛ֒�W��X���`|�����t��@���H�d�ݡj0g�=��bU.�3����´Э}ֲ�� Pg�=W�/�Vw�p�{��ȖJ/�r�.�-VI/-����;V�Yu���\c�L_wkYP3��z���!�5��v���'#>�Sn�-+�},�tc�m��{�ku���~�~O��{�����$��#�l]���>�aa�æ�F�f�Bɍዊ��� Y��/+l���B�}�����<�oo���znn�s�>]D�WLOj��s�)LT�6��Wd�^h��:���$���lZ3�.�qr����
W(!�����w�YZo�9�	�����TL��:�e�a��`�|k��	t��jM��by����N�h鋝B�H�]�c������T���n�X�*����'H�����swEJf��Sh.���ن��wp���+{	3(�8�1�;��6����V�~��(m՟7u��|�Z���턜{�s�꾧�5~;oy.Y��,p�U!��b��ubϜ{��9S]O,�!������1mgZ����\*j(Ջ��ʔ�[�������[�)�[�}!jȳ[ݶ/�h��E ���Չ���A��o�|.^���Ƕ��=� s-9(��Ky~;YN?
��6�>S�=���pZ���!
o2�Y��ӯ:pWw�,u���e�"�,cj�4ܹ�V�c9Ϝ�ؙ;}�{1��/yW�"*�(���3��CGԪ�^<�U=@�s[0ɺ��f��M!%��vܼ.�G��t����2�v,�� Uu�2�*k5W%_R{��!~�ƨ���T��
���E�`4u]��1d��s;�8'Dm��M6{������p���ʧ��v�dk��m�學q�f�����V�Aۏ�=���9MIc�u��fX@sz�IG�煊�gq�ѻ�%	ԩ^���3y��9ų�~i�l�6Po��m=�\iY�l�.̥YX?N)�Nw,n3ͧ ;�wn�Wb
�\���5`�ݖQ����xp��a佡Y؟A-�W�?SW�~�c������1�	�S]pB��wWn�(�$�Ɓ>�Y�zl�n8j,�9M��]��yn��}'�y�E��2�Q|�8f��\Co����h��ޚ�{;�FmK!��S��@�)��@�|/vE�Kq�.I�M�u)�mo)�Wm��CӐ{�>m���F�J�gS>�1����W�ٝ,m�{�z�[��;�|+Voy	�YD�Gq\�90��M��9����ʭb1-=�r{���w�Ƴt�]�+x���O'(��'�
���Sf牯a��7�����޹�� �>�u���RG.�����Y9��/x�HhB�-����������(Edp��oDf�N�GP�.L��C���S���R߽n��&�ELƃ�{#.ƫz�ӏ��n�r��Y�+ED���}	H��ѻ�">ٱ���Oi�b��u��&j����[Ob��=��s��:��K�[�sV�PM6�~���[��{b0άA^9�
̡�'�!rK(��Χ����}��e��t6`}�b´vV̜UҴU>�iǮ�Z̦Չ�-��D~��r7Nn��z�0���_��y�g�v6��� ��O�k~��bg���޺������O��-a��P��=Jyd��^��q҆ߒ�s���������
�B�W%��{'d�Ɯ�µi7�1��%�w�x����:f���䱽<������g�pި�S�ڙ �m8W�o��R̓hh�9Vx4EF❁�Q��V�Il��DNnѳ�,�办�����L�(���u�Q��so����^Wmʺ��S�5i�ѱ�ߡ�Զ�V����h�C{{��&2�%���G�B���n�M�=��]c���i�63�Ml��C�b���l�����ݿd��F��w�˓kS�S���ܼ��uwb>����B�x^U����g��#�6�(z/��/�KyGW��ޟ�����b3V�V��(�>N݇�ޚHU��Mʳ�!m^W7�;�"F\xD=�ItC���Ŋ��<k�S�#������U�Z�o�6�we�]K�;���y�������:r��*Ĕ��/6�o1�_V2�q�}�vgT�.Wl#����k����oX�c_<�z/�+�apB�(s(^�Bm�Lᰍ��Y��3y���!���ۻ~Ⱥ���Lԭ�`���]2��N��&�Ў�ՒO#���ڨ��������K}G���&I���,����K�j��^���e��c$o����D{}CL���+�*����x�;��w+\n&_<�ŧ7Lm��4m�VNfjd�q�������E\-�ٽ���&��N뼴n��T{f:`{���J���t��R�(۰.��A�=��d\��̼d)%(�?h�K�w��` �{�������u?b��gy�׆g@6��s��f���6��+��b�K����-:\�.��=���=��ͺ�7m��js�xj���;w�>������]�I�3���cǽ��O������8u4�
��c�N��FJ�F�)��oʙH��W���g��hq:��Z�:������Ԏ��f#u�;���f,RQ�f�ԩn�ߛ��a�*)�{�t�O�����U�HC�
���O4,�Q��F���鄮��yC����� �1�(NĤ�1n���ſY�T�����m����X^u������������Ag,:w�iSSW�>O���>��@�������E����7X����d��o�z\\�R�Wg��%�ɪU��vȅ�m�fb�Q�g�t�Ί)��9FL�F�۫ڑ�4��Z;vZB��U15Z�*��_�|v���tY��b�|}:�f=g���td��xd�W��� 9�&��~����J�S= Frѱ�
�tGM���&*�lO���#4���K�a5�!�l����w_�m̵y���{���;v�,�_���]y5������.�z��
�]n`��6Ί��o��Κ��V��^e��j�g��t������8|�=^�*Sw���q���^�
y��+]%֧6����(V��<�Ç�($��
l=����5��j��R�V!�@��F�z�ɲu]M�4��HF�PƊm�����.�(`�<*-Id�hK��M�5�Y�n��_*8���$N�����8��i<[[�q�k����o�6̼��Y ]��OS�+:Y�7�m�Վ��EY���&s�q�]����W5^֯՞�v�̊���HļZ�]�	�(\؟;��g|��Ψ�4%�E�ԧB39�EC��]�3��{=[����օ�d�̘�F{f�un��-	��C��Vޚ�	]-i���:s0�[6�����O�4��1�ι�
��7i�w�ٷY'6Ŏ�bm��;<N�	�[�i=S)�m�x��9�oǵ�P��P�=O��2��[ �:T@b��~���� ˮ�Ȗ���!�F�SIT��{N�WZ��i�/6{9��
X/�
��;a��W��O�u����D{o���HV��M}t�~#y����v���5�d�1�+��v��U��b'���(謽F�n�K6�!�=��&���y	Pi�;+����05�/W
C�/�WTN����ƇEQl�@21�o��"3�'˩�*DZ�9�O-���;���R�ZWH{�u��3b˛f�@��[1�l���0.b�:s�����u�����:�k��Ed��!���k r��䝛���h$�StxH+c��c�3�YU���G%.l�鵝�ٖ��W�nV��r��M������6)lH�<9�{� �Hc�\}5�e0��%�P��0G��X�«�F��WN�v��zs)�A=�0�^����ǻ�Հ��Ǌ4:�1w���Ɵ�J����R��(���g_���ꖵ�s����zn�3x��O��=��;HY�w�L΂�^��$��� �N��*ХQl���W��G������ۘ�?��N�ǽLV�����%WM�~��椖�#}�
����"�%Ӏ����&�����P*k���/y�ճ�O�Cy���/>��XewVޭ�&g��!]��i�P�Q� ^���P<�'^U��w����8�U#�¥쒍����ESw�ܘ��:��g7���y>��=.�;R�� e�cS�e�u}��ރ~�s�;�{�<uW����ˡ./w�E4��d��E~����Dë!a_Ut?1��-�4�HP�IhQWru���yC� ����!ze=ݪp��q-Vh��l�Zp~6GZܤx��F�i���p��鼯	sA�wm:�t(6��y�q���8yf޺��+����[��ӅX/��)Y޾Y�RK�[Yu�����(���3IjPB�+���_IYagY.�i]eXZ�.,��!�IԾ銯-�Q��p~|��;J���J�wXk��a�:��J��Be�L<��̣y�Cr�'��	���鹐<{�K����Fc�;q����K{�i�zs�͡�a��&`��غ��3�]����N�r�tS�p�K.�n�����F�¬�Fl��:��I�2�9���#�k@+�N��[��s[@=ͬF�o�k��p7ViJ���	)dF��*�%��i�3�V[³'Zv�uյ;.ח�1|�$�׵l$�����+f!D�������0b�v��u��L��V.^�MGeiB�ڃ,[�q�E�����': ���%l�pq�]j�F-)��Lf뤻YC�3mw�K�hkzrѺ5y'N�)Wm$N�s�
�[��5Ǣ����p��Z�4}��K��X�o�gA��Q���j-c)d�Cd9*=��d��ʽ����N���9CtpM���vQ�Q<��1b[�gn�ԭ�k;.'Z�w_Rz���vs9̼���W�k��R]�qL|��ݷ�d�B+A�O3���;�J@�f�k�7�u^w���Vo�;O�ӻ�I1���|#�9ջ�ge%��F�t�J�����L8r>ݬ�����o[6���0�O���%{+�:��%��zt��V��W��4�i�.�"mdY�'a��-�:��
����5s�mc� ��tc�`U��y}?ag����Jyo�q���=���"I�w��#�����Ӡ5f��Vө��f���s���e�z%Z�g����e?|��M�e���v�������-``�	�i��%��b�Q�7l 6-�zi2-�h싑���]�.t���O\�iT��aH�t6 vif���^��J�et�u�&;J0Ed�c+�c+�v�_N����Q �~�х����/B��wk޾��>�nek�B��3:�8S;�_4�­�M^9�gW�b���ʖ�[���M]ٳ���:�"y��Ŷz�*��w�2����L�F:m'9����h���a��w�3uS,K'k�Km�<�ӱyh0�W	��m�ګHrAk�儑����u���I�N���dر-ؕ�ok�坨�%�)m��ʞU�]o����
����ڳW�J��&;�F����+i����1�=�pob|N�V�B��ч�f_T�*��b��S�;m���w�w���)���l4�̦��v����J�eիKmmV�m:}�X���Vq�q�ȎF���MNΛw��d�x[�w�v�V��� �~�I��+r>����苈��+�Ә��`���җPO���h��v�vu�
���h]Ev����&�w��󅻸�|��S1L{�Nv���9$x:���*�4�z�]��z����{�*��d�T���_�C���\���{~���,��c@���:�ُ�e}����V}-�Z���ִ�c�'�K�;A��W��u��VTI��#+#��p_���N�r�i�ZW��ߣ���B��R��e��,��]*�2�2z�(0]<v$=�~b����
�[�!�\�k�98�WtQ��Μ)m��Eoܗxe+���o�/�n�5�:�T���5Bs�D��<N��"�������7+�+GN��8f�Vʹ=�Eoy0L荻v��!Νg������Х��ڝ+���/0Pv�;���Q!��Bӂ�|}�O�^ʏy2�����7µ��v	�Ҧ����j�S�X|MBѳ�X!u\`�Ǹfc+�߆��c܁]s��!��O^vC�_�N���)��#����gw�;����\��u�~���"�G�؏.�/��C���W�t�&�gn06�_]98�^�y�J9������j���X��-9b	3.�aą����ᵼ'C�F��%p%a��L���مu�z{T�lM�u<�ݵ�Oup��j5+�����ސeɬ�ݺӣ,�k���[i�S7�jc]�ݪ��z&Vմ�x4��i��|���E]�ǜ\�;	�S[�6���%u'��W��dE���eʤ�4Tb���S�˄F7c���F�mI�J`I7`��{���݁0����:����ԗ���:b�7%u~u��l�ؓ�YV��Lo�sT�b[#ѿySDu�/�\,�*��>v�zrr����S�;@%Ie}��!�r�{F}.��x^�/|�p�0Z5:Z�ۓj���P��}�?���V
?{ZVq���-�W�<�w�ff��[�
5���2ch/E�f��PN��C�aY�}64���8��R�J���I]⍽�F�w��	�No�}/�2b���d=�+��O��:@�����E"��� ��}��U�}D4ò�G�8�,��Mק:�³�vn�x:N�����4��w�y�i���lTYO�*ΞU�'�9ɿ(��/��][:�_�ʩo�aHK�fȥ�=)X����OxY㘬N�h��?S��2Ϛ\,g�9���|Ν]~�����ޞs ��#)e�8�E��.7�h�?k���d�i4A�.��oXz��ř������ܳ|��CbL/Br�J25�>���&�ɯ4u��P� ���<R�.��i��ʬ��2u��^Z�k;MoLeud�鑋
/�k-3��=����d'R�3����ow�6�
<e��̡CH:s*n�y,4��fRKiU�V�.������[Ĺ��n^T�j#H<M��0�,A�3�D	-)���G6�L�$5����=��rs )0��Y�#$Y����:�T(ң&�.�U�n� �̋	H4e���v-�����l�׆oQ!�������iC2,�!�dCq���dF����"���$�!�W{��B��5qG$�<�k�i<�Y�i iaz��QC#���%��ɀ%�����Y��4�И�4�N�#`�Qa�4�2 �秲�2��>��X9Cq�9w��**�����ۀ��T�6GT�(^x
��n�$j�>4-Te�Sڪɴr���v�C6_�x�ژ��<��[渝�Գ��QEL��Q�%���x���`���R�7#�#�/{�(��}�>�L�-�	�����:/]L�?m��y 2���~rc�8�y�3O0aJ���t�~�N�.�ޖ��y_�J��'��_�;6����+�����+=P;6j8?�{����TҞn���5�&
����9�N���=�[4v��)����0%U��<�-��*[�����Isrn-�Qa^ߓ]����k�m��
��>��u�l�g�$k�O��2��4<^}�������8�{�!���Db���L�⣻��e+5�Ϙ1�@�L߁as��k�o3�lc�WL��ߞT��(��6���u� 9�.�j����e�4��Ƭ��H�,]��h�un+ý��_>��d��e��^Nv��s��K�F�X�C�L��ӊZ;- s&Sz��]�(:��G^����8�Y���D��_VТ�rx�Ü;�tn��x��%�����G���9�+��H??�A�S˲:1����_z�W��=��o�~V>���t*lZ��YΨ�;=�.˃�l�|y��%1��^j:�&��u�y��X�����w?:��F]�o��L\�R{��a������׼fSR+���f�'�n.�*�n��%�[!�/�~q#?Vފ8h��z��N駃���V	���h�'�>���P{}y?>#g�Fy�yU�E��f�v��,��8��uroO����{E�o�� ��؂g�ş6Pk�u^�^4��pN�U�uK"�H�k��w|����B�ES��/:/����oB�<4ȟqu� �#�����3����fR�������s��av
au�~5(N���>��w�;�j����ٔ���6	~��3qE��29�K��B�W�tE۪ѫ���gBow�I��.f1pZ9ѳ��y\t���]����l���U��r��HF,�`/R8R�dVNR"</��wh�6��j����Tf�ҏF����rE5Gl}[�n�p�<�N��,�osrf}�X�-9�*-=vu��*F�ԨlTCj��!*���;f�֜躻.�+Dݕ
�L6Vr��s���Z�$��u� �Wwz��j�ya
�ef��C`�oT��G�bsu�Tܘ�N����}bwif^}��A�>�h_���_�8g�pr��c>5�v�|usT5yP���*�����fj�3�(�����o�duŽ���9�i�LF���3�z�������\Uc�k��3ݠY�6bу���"�9>����}>�O���6.�圏�+a}�:|�K����LQr�uzE�p���.�ޯC�W!凜�"����T�������1޶|�e���o�ۇ �~X�2�*X�Ӟ���}W��!�͓�~�菪A��Z˘�÷( �d��^���'<�N��f!�>�'5w�z,�g�o�W�4����or����dlWx[�w���<O��A��a���h�:�O��������g��ȫ��!�{����U�uN�@>�h�Ȭ��p3�q�O:���k���S�P���G�ڃK�h�p�v/���|�Gc-�h踚.��7ɂ�-݆���h���!��-�u|ڕ�Ph�w�zU��E�rIqb��T���ͺcݣk�NJ_�nP��zw�gUvXݹ\���
�Jrz����ǅco�g��󬱚FU���mZ���z��-�?oi�أ�Iڗ�K����5s��d�_�ŕDg�9L��W����-rV�{je�\�G4���Xgca�Kz��Y[v歁�?�/z�~lӉG�nXc���'"��NXL`�v<Ҹ�#.D��}�s�{�\]NJW��>ߐ�qV���gt�q��^��]ќ��X�cC΂� ,C�5Jහό�tM;�9�a>Y�ܓ���=�)\����'Ն�:e|q� ��Ka��,A.$���q��Iw�Aѩ����|,��*Ӻ]xA=9�s��>�IZS�i�]�C��3�w�tWY�6���h� �Y�:���V��I��=B���9'o��|���Z&����Z�za�On�t�&���j]�B���?[��S۵k#39��g������a�ggn.��\#�l�(�B��~��)���ݬ�~�o��+%8��j���Q�=UQ��M��;1϶G|�v�ϯ��9����`/eBv�ǥ�s�~�+'��<����k���/����V�A�/�yĻrb�O	qy+��'�̙y@�-��D��wth[��x���Ϯ+%���L��wCu��`q�Vs��!��O�-ɼT�k,�v�fbk̢����ֽɻ�~�CI#�~�/8�A��{9�)=�E֎r<H�n&&��MRB��}�b宝�{�6�<:�f+}S��3�2�a�[�Q��7Ҧ�E�5�J�� ,b�5#R��|ˬM��=�yW3��W.v����iZ�5����^ʸ�&{<ڗ^�)U��Q��5>���-�M���,(�u3F\%�{C��Kn�e_�3�K���Z�!���|~Ϟ�`W�-NiX�-�}��
�����o쯻Ȼh���`Lof�T���+��9s�^'v��>Y�l�Dz��U-K�kP����d� �FwB��.�����%Zv��H���� q���^��´A��heq��L�C>{������RŪ˙�iI(��[�tW()���8�yw>ꐌY�H����@��t�%�dہ`\�,q��}�b�;ELf����~��K�w�Vn�k
����`ZW�.�v�=��GR�"�����fv,p��cʘ8S�n���d�|i�P��7���8K�[�}�9zn"�����z�������p�e���^]yD&�І:w�q������F�/p}��(E&���nh����))���WօyJ�^�y'��t"��-��d�K��)[�o�R�lU�\��
��$���~ۨ뢷;s9ը޸�V̀�z����d�o������PB�ŵxjc�OP�e�Xg�ݵ�F�Z�7��.��յ�-Y�D8\R]��	��zN�%8�w%'���t}MAw�U�%V��N�ى�n����5�z�����>��r۔xR��d��w^�9�����
ٙ��K�����f^�B�,"{��'���-��Y.�{��$�9���j��X6��xfv ��rM3��.�Ŏ���f5������;}�C��,hXz�%ꦖw�t��' #~�"�iVa�&dxϫ�sKpU��m5 ��C%!��;�STJk����=��&I��I���Ք7 M� i~���j��r;/8VY�����-�ެ��n���ٽ��أ���.�����W�[^{���Dm�I�s&b|�G�
�H�=U.j��>����3�
�S_�7=`n��.I�-ҳ𾿘�5��]a&�vN���GG9�p�L�|E?�#�d\v4įȘ�T��\����q9��LQn���;�a�y��Q�^�ֹ#�g����g�:ҟ���^�WC1�>SL�h���w����u�^S�I�ۇ�CGw�U�b��`ڵ��	��9�ׇ�O��@��9_�[�g�>�h�zw[�:��OO��X���p������]���J�]ag��[c�`B�?Bz����jGݤ&qF^(݊�cf��G�8X�Z�2��q��F���f�6��9�����{�S˕�k���N����0�ʎ9o:���3W� f�[��b���nÁ�jWp:�M�a� ���z�-Ȫlc��sa�.\���d�c
�8-څu6�DKr���w��:E>&wΒY*=~�����Q���X��k;wbTs��|7S�Gf��(��0�u&�e��O8���\�3}nbX221Z]�LGw�-�o��R�>�,P�3�~�����w����۳V2�u]@��L�`�
��1��B��2_I����	��۷�j�k�;�K�0n���$F�33�{T�y�遝!9��y׊�n���)��������;緎��-|� {]�~F�i含v�>�nG�ۘ�� �;�Ozfn�&���+�f;~���l:^�Z��0��Od�|�軳%�HE�M���>��m-rͫ��LQ�0{cq��I��#�<�9ϕ�f���zx�n斺��$��ͯ{�̧ink0�/
�b��m�-n��QJ6/en�*m{-PPlۅ������yb����
{�PiO�.��s{���3��?b�fgƗ����.f��R3�l�o�OA�װdܔ�[�iuiKh��:���zͦ�)=�J�o�`M�D����4�(*_>9f��J�56�U:
�Ω���N����n�Mє��]�D��'iT���nI�]�b�n�G&ŋ�q�����sv�&��4_������w�
�e����ab�9b��u����w%��dom����s�#��߱�_�o���_��f�'$�ζ��n��v}�%:R�̳�Px}��Ȩ?�!��0��S/�͂;�k.f�I|��q1t����ɛ��s�G�-�:���g�E�m&g�x#���hV7�CY���C|��+V�M� *+��δ$�I��]����ȋ���i�+xƁ�N�+�EIt�,{�Ů90,߮A�<o{]�{�>�
9��1]�s�q�r�rD(�ڿX�>�B��߳/�lF*�7<9R�n_���y�iA�|�ż "��Q���f�V��1��&�K:��1Ly%��4�+����MÝ��߹א���&�mTNV^�J̞�J�`@�]<�����'r�<.F�ϩ���Bd�j���@���]R]�)UB~`��%���v�wJ��Ƶ�\h���'5�3�:n�KV{�s�Dh�ϕ6Gn|n2s����羊ex\]�,�>P���V+��"<Q.��������w���o.�Yk�/GxO� �J⥎�s^(��>c�%莄G�>?�͝����en;����H�6�\�Gi^ˊ�{S�e�3U�z��eds�*�U��km��ax$ePf�[�T�`'��J�]n��6HC�Yd�F��(P"�r��w�̢CL}e0G0���F;9� �y�81K�ش��1�k�Y�:�����dh�6nBo���k���F���cFs�V�ԗ����5���}��Z�]N�j�V��A�)]��%=���5|���P>�Q�[�B#�0{&�m��+�X!�l��R5�kMKι+GSZ��ۘB��Zy�W4��8���:�!:^_f�R��]����w|h�&�y��wʄ�3���u��h�Ǘ��g��d��R��윈�h�E�e��v���6�#kHa���J ��Cz�]`����Гxl��-	Kk��Մ�E��J�.�NB����%���Q�T���Ii�N���To�y�p)H5T����e\����Y��UkN��;�!>u���ᜟ@�?��׆��`��"��H�u	���z��1
�#�|��V��
Y��O������-A�����ci�n�uG5r�arv7x�-��o]���K��, G'=�����hVu�U�EcB�'��5X�,�E5�{��^��F�J�S�ڳ;6,tCh�3gX��Fz랅���,6cb�<V�K���S��b��W���W3����Hqs�Hv{X���.�ޚ@d�5����s��G<��0��A�]�⧵=�aS��|���r�rr��z%�X�"g�/s���.g>SX���o���W�MZ�����`��A:�ᳶ�����*��P�0N��L_�z�U�瞝ϣm��wt�Gd;(Q=��2e%%4�:�wofl��hh���H5z5�����-�w���]�پ]�Ȏk�1p�H�/N��ԛ-b�!M+�4�A���xE@ej��*C�>�f/���X@[�N(I�s��)�_\�	7v��|�A�g^E �
�Sy�t���b��wA1�Ԛ&���������U���g����� -K�`��]��E}OTk7x_,��	\c<���]��ە$���l�5)EY3z�bͺ���jl�����u�O!�6*�Ed[�v�p��ީ�:�E���Պ"a��ې�](4g���7rԔ�)�4�FY�$Ǽ�P�GhG1]>�6�eB���������nNY-�md�<!��6��v:(	+wQ�WP�]���:�u�r���3�zw� �L��G��^�=?K[�����ăC�Z���Ժӷ���B��nZFU��Gd,O��.`+�nQ�ծk�(�j�h�ݓ-�6���?����Wt�`tOD���r5�ZG_Q6�a]ғ�:�5�,毆r�9ί\��qV:}�N�I�f�8�m�؊6�� ���XmDL�Gr���}Smm� ��>��G)�vy[�
�����d�E�;�w��$�Z� ����ܬw�{+e6�xk$�uk9�����].�:� {j��`NM�^5	�lBڵv��t��uEƍqݲe�Rb��eݪ,-=%F�/7���~+B����7ML�k]
s�u3��:�o����!�#���L�����e�<-6[x��"�SoZ
�e�XFi�*�N���`z:X'�TL��f�W]kc!�jTn�n���*��_��̧^"�"�*�H�Dx�4����Z`0;�����Sw��@f
3�d�H}A��� <.�Q*�4<��?W��^Q�c��W@E]�/mL���9u�nC���D	%=���z�V�.N���L�Ǯ˪��̜V7��.(_>��!��꯬g�C���X�����s`B瑇<����W�}E�~4�캉Iܺ
�1vLI�*�Ѥ�9�ex�nz�<�2�h�I\��2��}3������o#��ޝ+�\�]$ϒ�]���Q~ԕ��>������v���i��,�jC�jNd��*�Ɇ�eG�����lț�{�$k�^9N���4}�ӕ�+F��j�z�ޫ�9TҾ���AӦ�jv�fn���7�U΍'s�}qy)<$yyY����{���ѳ_Y�"@�3��ԙw�Dc5*��LSbyО�]n��9 S��{UP���T�䏩:����2o�n�YCʚ҂E�[��3%����疅O{n�Ċ��NP�ۑ1�A���f,�A5W��+�o⽆;���s��u��ym�'`{$&yx�,�:ܫ�9�*'�t~<j}�����Ⱦa��K�� U��C��W#���0��а�:�:�*[�9�����:�*�d��8���&�,M�T�6t�\��������~�5�+(s�#9�m��#ve�C�6mK��#��u,���o���S��v���n����)=�Gfc��S�#�.cT/YCA>�ڤRH�s�q6���J/��{�#㻒�ǋU}���ȥCsI�R;��E'f��6ص@/@��ӴN�B��PfT�:E�Zoõ���K������:�}{	3���^K���DG۾r�yba[K|���ߵ�χ����S�aP�qRmwsv�}XW�9N�5�\+�nW�*���s}�z��WH{��>c�f=���Jz���z�ζ�Xdw� 発Zy�[�c{�?b�U�5��{�Q�;8vo�`�j#�n�o��e�U�f��d�Q�.��՜Қ�{4��u���`�l�P���A�����2�V�_���t�QӼ]������*�q%���̹�=�������*��y�r����3:�w������Y�r���v.��eYB��{��`���?D
�n�UL�$(K�m���U��j��l����
��+��U?WZ;E�u��bwb�gD`���U*$��?`Hha]�������(%��i�䝃2%ȕfn��hH�UT#�:�|�3�ru}cEb�x3O[^�9��i&��=|c��6Mh����;	�"�5��8�ַ�)�du����ӂ��L�;�R�'6jř�E{�ّn)����`Zq�E���6����W/c�:��t�=��k8U$��q���+^M^�G.[�e��Hn�nN�9E�;�!:o�骷6��ɢ���C�V������8�Ζ���U�gX�6;u�]R^�,���C���8�hg+^_}�W�����>5L�]��7yz��9����qwF����#bME2H��NT��������٘��<��*�j��Bu'm�yj�.�AR���v� ��t���O[�-M`Bڙ�a�+�럽�T���q����q�*K��v�O�*+8� �Z���I/��p���3B<`Ti �,���#�ՙ+�,9>�ޞt�K	�f�Wn&�T*�\7l ���D��n��sv�|HQ&� �#�Ċ<T"�#.w_FW�㡛a��Tx����B�h��7�,�>�X�M������Hء�Th�v�'mUx�-����|υ�ڔ{2�1�������Dq���{2���T-ԏW���\�r�Ԭ��/ez�T�&����|]�j���9�TN��J��[��$�X�z���of
]�|n.�)YT~�����v��J���[u�aP�a=R�XR!�51�*������]�F���66-g���gO>嶌�סI
��̝�!ją�������}�cG���@�]QK@!��c-R�5.꺽JC�}Q��b�<��R�΁���÷��oE���-�]�I�w����Q_%���"�%�ϝ��~���:��
TmG]Qڽ1������*��Ծ��h��nr����.�뽠^����0a��-Xk��헗�C&��T�')Ltr���N���vp��B�}�d�lKu�S�ޝPX���K����p�[> eG:Y��w�$��ֶ~�:xȝ�f�h=7{y�vLì�oJi�޹��}e��Q� [���.�gtjj2M��6fث��G.��c�X��>��w]݌�+�8*�R2s�A���<�P��eL�ST�^�3�LT"��;� �b>��C�_��:�����7y�ㆦ��p������fkW�ff�S��fV���.{�kA}q�0ƹ}�ߍͧA/�6��z]|r�i]�n\;}�[�œ�v3E^��	m{�{�����>����+Ҁ�u�����7�qr��s��;F����7�DĴ�u�������{�|�#V&z`����̔=.v��!mei'���Qy��0^e��.m�6������eP3k��"G��r�j�J���c�B����o7�κƊ�5�~*[��j)�WbzQ#�G�6kC��^&�\9.O%��j/�a���Q>�חptT��Lf��Zk�Ӽ��)!e��T��їk����M���4z�#�t�t��np�;E�;���bR��3O�����A�y�ozL�s
3K�cN\�����r:ȉ~flZ�WO���+Mc硭�6��L|����#�m&�o�(gg2СuR��6r&D���g������Y�$i�V��釸{�\kK�5�¶N����$m�S+k*umm'�E�r�#�%��x��啘�`yM���"=�R����c��נ�����c��:J�Z� 2��U]Ļ�q�Br}�������L]4���\�l��3t�Jm��]6�:�ͳ&�מ�8t(����P���خSʹ�~��5�?Kƃh��������s�hK.9�T�p98nWz�.���u�"+m
-hz*%��N�A}F䟋ˬ��h�o��y���yjog~����^���15�ueAcs�Z^�O�G�*�c��=�Iɴź�Fx2�T�,P�W�6�Qz��p�ND��)k�Aha��N��b��C!h
�ވ�?m���,Q�c��������Tg����t�K9Bs�=q�P��M���4��������j2m\�ک�k:=)K�C2l^1�8�y�zU+'�2G�N;10K9b�W��oz����&r]�l!��=����leIȼ�q�����r3�Su��|"��NN��u"Z�V=:*2�#p������I��8�T/{ٜAZ�YܖU�����c<���T��&�ͻ�i��+��YX�.�%�ܧT�îף�\�J8U���Aݬ�r-ɂ��;�O�ܶ����,��������}�d��Lto�D��=G?z��S۴~�n���v|����d�*$�'8������
��P~eܱ;�`W�甌1�>���\����s�Ȉ�ʯ#���0jcV���;ܥ�qo.}�p^bY6�H�������u+�Z���k7$UVI줸T�*M5��dY��4@�/R�Z��܍��X��n�W����&����^.�=�̂.�p{���k�};>�/3�JeU�������W�\��m�zį�K�a!/08�L�:X��'ٛ��K�T�|͈�7�C'ى���8����99�n}�VeG(�䷋ا4�:y��<��&�.�̍A{P�GSC��o�M�����Ihb�*�vo=��:����]Qr���7z5LE��"}���N����pd�^jb]�T� �I���pDQ��ct�^�픠�Rr6�wSsN�BLE��H�?*2�c��B��=Þ���9꩹���T�}��e���@1�z�����1�x��+ނ�S���.\Ϥ��5J'5�Ep$޾�;f�l�<���޺EB���*7j+^*γ�1R��ڻ�i^���槌����4�L-1�;�vO/](>�����y7p(.3ww?��5*����#lc�T����!���y�󋥛�ˉV����\g���������=:~A_!R�}IC~u��͢6���WuHج�N�V��b�v�*d/���[5�y�zf:g�8+�b�ssO(�����T�u��O�;���/�M��-��g\c�oEw(<UM��n�'&���,�ٲ�x:A�&�O.���S����;�/"�HS�0�m��1��T��e駂�V\�����"�J���a�3�V[Xn�W��z2�剪�w����3�C��Yw��E�uv�[	p�J僚�O��U����^QL����[�!��G`�*���ȟ��dn���j4E]q����}�{x-��[��"��R��<�1��
_a�I}�t�T��/c۝)�ɺHVX������o�{�����S9�����{>p#�d5t�=j���%��"����&:��bJm15B%C�=G{U�t����[�ձL. #��X�b�Iq�����ly!�86��C��4K�9���G�&�U�+�^S����V]��z�e��ᗒ�8��ӂ`����.���)V��ځ����c}zuSCw����w���}}�Ձ���O8[�V�)��GЏK1!<�T��~�u�tP�C�5Р�;��;B�Ҹ��L�a��4�rw˪}^����m�Mx�\U�3>Ԕ����UTu�&��p��AN�e�8XnxH]�c�����]��yg��49)�}�E�-^h]�R�Q�0�^}ɡ��y�Q��q����s�`+�I�\�&2M���:-�㐑�&�9���8C�����1�k���h�y��[�y�Q���d�x�S����'t�E��U(��άB>�1��]=[��"n<}���0V��|�mj)ԛ�D+�3�K��o�)�V���r�J���f�GV��ڷp|^����O��"�Ix��3�н�Y���t����b��$X�P�&$tK䮜�64a�޶�z�]�YY������L [۾ټC{������w	���m���Ewrۃb?ĭ5�.�ɻP�����Ⱥ4�0�deaP��_]s�9�45�2o������0���̥@�� ��Ρu�]#�5�F�N�FɅT�Q�����Ψ�:�ĺ�u�)��;D���l�8Q���a�8f�����D�'ӄs���ܜ`������n�^4E��qp�uY�lo�Q>G���T����a��x|K��=�򽊌*�ދb��5-xI�qM^ 3} U��+�E��W��ފ ,Ћ�?��ZDP��M��R��j�Pf�AT9*���n��ԟe�� ���l��p���9�R�2�l�<�n�R�ln�Z+쨆��|dF�MqLo���a��F'2Q�����7�(���ע�"�q�J�Z���R������#��j����=~�Bۉ��z��K��kC��Wc\�|Q�޶��c�E���~�?O9'u 	1��6r���̇���!T)����w&��������e�cx�s�aP�DNf`�Z��\��<䢇��Û��&��T��],��S[��U1◌f����>���Y�}'�i���iUS�������9>�^|f�%����{��<��f��p���W��1:�~�����e`���/��k�T�=��/�A�v���2�%-�Rv'Yb�,8�G�XOu������2��/z�ǚq�en,~[*l��tO�u���cu�Q���y��;�Q�v����qWKb���5�\�L�g/��of��,n�kX�{�����,��C
�8O�<k(�h	�����/}�jf`�b�*���Tb�F�q�!#vJ4:���|��u��]}���u��e`�_L�*��x��Ϟ� ��Bz�:�R<�
�6l;����<�}�	���n|ӰY�m-�w/�R��3�'�B��bSP�}��>�P��z�~���rd������{>��k��*A�]!]o�EJ�³��f��tx<^S��$�=�������瀈ǂp�2��以R�3ʳ�>};��T��pj�t�X�#'�����"o�ҕ���1ٽ������n}���ɺ&�a��{��N�CD�]�`�+���5]U�=q^|k<+M)ɬw�%�����1��lh�[H�=�1y�m,�ö㗕ɻ̻*MUO-~�!ۗ�y�wW���?	}:��������W�Z���{��zb*��/j�D�F�u.gu{ �r�m�]c�qX���ks�1"n�5��7��/���l	��ɱ((�,�cU\"�%vq��=֧D�}�n��[Md�g�⫫.�WY������vi�ewmdw,B(��H�/s�E��2�1;<e�?'��S���7i�WS��
t��EG�
�%L��Բ��g����*4�*S���8�:�6��7�bM���k6����X��+��U,�ծ0��o��E���]h�J�Q���MN&'\��X]�n�z��gV�5�N>��3���tC:�����L7����!�乵��������c��P7����.}*d���ĩ��j8A���O�b��(��^k�nB�/D�{57���\2�om���\����O#��j.I;�O�r)�.2�Nfu՗�g����dyŉy�ᳮ�Ō���O�_H��|�_[7��R����v�n�㯠3��7�}:r�n��ֽ�hON-�½���rH��.���1ϸqi��y
�d^�8���k�Y�Xn�"��i�t���QN9��]5n��ݻR����b/��٣��*xx<�v��`���dB�By{��|��ܒgِ�o� 'n.:�݉jS/{�0OfUF��|��'y�>��8��Y��2wr+[������h��2�G�3���=JU��y!�+j������e�5Iry�?SWi��n���e�٩�9d�<�����Yw9����tOT(K*����9�8_p���;mNL�戛�v�˻�!�wO��CԘ�e�4;�з���u��NP���73Ⱥ�*�h9��&Y���7���3��,��x5ȑJ�J��3���-U�+,�:ܞ)��C�J�xf`M�W�폕z�!Ge���п`���t��+��@��dTOr5]4��L}
��þ����h��)���"��4r����V객�n�Y�ZU#����-5B�#�J��ik�������XN_���p榈p��Iu{��0���y�/�r�H��.��!�ƻ���vv�<��xC$�F���QML�0���+z�2����hEs?[�oj�#���l`�sD�`�lqN^��x�H���G��ޅ�1W�R6���nf�V�P3����D� ���T�Xҹ��vN��\7����T�҈v{Ugj���\�8��
���ml8^i�K���k|r��,������S�GU�҆VbPV�]E��ȬZ�*��e�è�۽�:��7]�'���U��v�0-�����]�
T�i�k噿�]���Ԓ�xxm]�K��k��8�m��d�{M�ꇚg����5����m�[[��DQ��g]���eLw��1k���wV��0���V7jCulS�{'e��%��ԵI�n��is�ӡƗf۶i���66���:K�Wmjnh�<�9a�����5W�mn�3�L\�"��S���
�Α��~�Vf��3��n���J��Ⱦ\���/�/�����zt#��5���8�l ��[7X[�`��U��0�x��x��H��Ve�Aiv�@�^�7ܑ�)oD[�kKۊ�
�.��J�h/,w1Y.ͦ�?�Z�\�*�Y�x;���L����]�9@���=���4s&�^�|�b=�sOI4�*Ŧ.nH�F��&�#�+�f$�#�ܻ�sn��;����#�^���l�:�d���n��5�WJ�,C�v�e���q%�t62�B�']��4e�Y@Ԋq��d�Zi�ȥ����2&GV�y���N�u�j�܉Q�{��W��T���ށ����]�����*�ej�X�{O����I�t�4ҹ�n���Y'��S��R����lh��L���C-��׆�/�CH���ǌ�9�b�N��r�&b����`=��_i��N�ի���Ul^���Y�Xf�"3�FzV���k�\ő���,�~�\O
���!Ԣ����G6��f��Wsjat%��}3��'7Z�]��=K��ܬ"v�w}m�;d�x��<�r�7FGYc������(�_h�#oR��-�Ԗ�ZA@��wM���}��3yK�ޯOx��h�0�nѵ����O�
���lO��\6��[b�u<� ى;��]�I ����H�T��
v9ft� ���1���^[�f��)Q\q�^���A%��6œ9���拖��+��|D(�!����pۘ;���#����E�����:�Shp��m7[�B�<�bN�VK"�c�Q����C�Eᛴv�T����	]ݬ6��}�ηgc(w^�`�Qw�30V���EHu���PS�`�6�����v��0f�|xJ�\v��+U�{X��L��E�^�slls�[��˝�������Վ���9��Yt�v�ڽ��n��˻�\eq��M�J�g������^V�+3G6n3Q�
�2f���:]F�~���qRd���~T���G+�l>��J�S�U�{�P����>��>���/�Y.���m�{Zi�¾X�-^��~��ɰy�����S���2�Ɠd֜�ҭ<�#��%�q3�n��('��GoΘ{tQ�\�ɝ��ҳ{�Vx�V���6�7a0|d��2'�	��B��ӎ�>� �0^zC��o-Xc^��"�;�ri�ٓ�r��0��"f&k����Ҽ��,�}q��|�W���n�˖W]���*�k9WQ>QuS�Ջ;Kё����è�&�{�LmӃ������7}~
]>e�� F�עJ���d[F���{���:���^�Bo)%/ca��.��QQ��U㇮t�7*v`O���i*�O���o��!��5��V.d��|���Ӯkt��Ǳ�μ���Y��|ˋ#e�|����y����/.H�犱�`H��z�1r�,�SUF�u��MFmx��'#�!��J�v�	y���`r8'�WzU�5���ފkz����ɭ��5d�Ud�Vp���u���B���_��twg�S�u]�T���gz��r9�Jb���!e��j:�� �,TK+��'��9��^F�E��=���x�.|�v��ݴv�74]j��Vu�: %���d�P�����v^.L�nl��v)5`�3kZ�-�yl5����r�Y�ި	�ض},��F���o��X�Wfj�##�!7c�.�;rԶ5;�Doi�y8��������>=k4��f�k,fYU�q�^R�����'*�+fCC�����W��^�>v�8�a�(��3/]�������{�Y�G�~��g�F:�qx�V��sE���I����-mϼ�F�r���[��/vk� ��k��>�	�n��V-G�d) ��
�v��-�B�>�u�tS����dx�z��zmNp��~Ƙ��H���y5����,1uZ#!�c�&n��j
��A��T���f�3*É&Ax�$��W��=��B_^5��{h�}N$��^PG�.��y�S�+˜jϑ�(Vg����ߖ�᝟���x���w@U�I��`%ڗ�oiT͇}��ˏ�|��ϡp��$�ӏ��=�c(U�y�w�s(���u���IaJ ���?!ȧu���|�ʨ��S�n��g�F@���敺��bt���&��czR��p��.���J��C�~���7�5e�g+����<vP���O��y/apVU�*�Mn�z�ϲ�P	�n�|��{��R��K:�9k����k�c]|h]t��U)c�>+��;5��H�SD��H��;�A����[��N��(߭)��={�!��0�霏%���+-B Z�Cl�_��1�W�������3��HE�r�����EVű�'��ew�sL�i����!���x)�!��v�M<�f��\�kf�P9~U�	�";��K�r��R��*��6mKz1����֫6Q��C�y6�@}|���S3v�qݿ6��J0��TF�=&|��&+��}���WD�= S�7���=����y�w5� �� ��ɽ:*yxm�U�KhOo��2�͉{N4g�q��{Gr7�5���b/�X���l�}�<�<����#��/����nȦ�U�y�[��P�"�jnA�%�ܗ�CV���c�z�3�'���a8 N���r�|'Φ^(h��Ռ���|�Z��
�Dϋ;�!c���sв���@��p$?.�Y���"�zn�e�R�g�&@�Y1b���රim���y��[IK��=�g&��^tۤ���w�b�(��/an��l����{ߵ��ox�F���	K+`�kB\�2�g���I���߸:=��pr�F���Dt:���h�;{���3p���uִn,���z؃3���п,��zz_�F�g :�Q��T%5�����U�V��x�|���C��.����-���޷��_NcFqɉ��!*�g�v�f��΅?Oc��J�*a��036�;�jx6�씦�x�kr|��뀇٭{w�o��Cܼ��} ���'i��d!���G��/1�¨���JW��$cۼ1��|R��8f�N��f�e�X�5�*��S�����`:�ڦ9#�c
+]��ZŚ��<s��ݤ�F��4�y�Fĺ�ض�m���-Yjr{.�0K�o�:vHw��fH�Uq��s���o'앓�Wrg'�W3|;�j}ޅ�_*ٹ뚃t)�J��%}n���r�d܂A�Dśޗ=�+�2�3U�;��1٪�}Jt�"�[��W���$N@}&�L�R=���,��<�,��J��k�E�x�z;.�n&�r��y��G�g��W4�	��<��]R��#q2`�l��&)e�3Mq��T����<�a��N窸��'	H��m�[Ļ���P^�d���Zwj�)p쐉��^�|6x]�o���f
H���c�8�����2Z�N�9zcӱ�gwS���w��1�(SQ�sڐ�r�D�!�2-������\Q�v��-n;{�} u��}�
������H�T�C��<��B$��7*Cgp>�/M��&}8�'2��e��[7�^�^T:f���s=UQ��U��;��O�����Nn�~�< S�j�5F�f}�B��᪌�n��+�u,�/;�u�������<�F����r31)�RiWfWhUĸL��;P+�:�����*�@G�����b$�H�#Хp�<=�R���0zh�	���1>xcԱ>�Q�qފ��$S����#S���4Fyh�_�geb˯�����we���
�u����"e�lh�+Wj��h�f�q��\��&��yϳi�t�q%9�9�aJ�7�˦����ܘVU��֮��E(��{��#o:�Y{S�Z��bW?L����{������?4��Y������g����yO����rǂ�[0��bM��0zY����B��x��rS���9�"����-jZԅ���L���E��"�
��r�/ ��� �_����PA��u�|�G��,�qxV�zn2�7#-��ڒ�M��.��y���2kN{F����NM�g�t]�;�nb7OV]�w��gPxy<��o���	�O=������S�{�F������#}g�_�Y����뫷4�={r��#=�Xy�D,��G��C�^����2�E*�E�j���F��ؑ=T|�x᳠�:Y\��5�Z��ꥄB�n�N�K���l��P���X�-g)��;�<��ޚ���u{��0���^P�11@��po�+h�X ��5t ���m��4�V.c�fx��q�@��F�CZ��(��r��2��Y��r2\��ʞ�R׫48���{ك�#��;J�[���Ur�ٔ�Q���g�_���F'I�a r���o��{�o�ϝ/��W9�]'��-���.��r�yAxH��̩Hz�X'�d�.�ޮ�I�l�<xۊ�Jv�<�6�"TcM��\/p��s���j��;��moQ�u�k0�冄zȥ'*�w�b��S��-�˕-�R��|���&�oo���=����Q�腗��<��I:*�v�%hN��������!����^d㎒����C����.^�X��A���GF���Z����3�#FiA��xC�m���isDw@�*�D�ev3ո����W��3���KQx�t|�� �n�/sי�Z���q�7���,�O]*���*���]4~�F�6����wR�W��S��z"�RǣFD�K�S�
����bs��Tl��r�'"�<�����^��Z'Kl���F!��Q����glίm���N@7BsD�T��sḡ�G��K/s�@B퀶@��R��g< ڍ�C�U�86����ᥑ,�w�:i\�eb>p*n���/��O�xܞ� p�M_����g_�w�s3�kԲ��W���3�UGL�3Nc�'��H���oE��Z���W͑�e*���Myaw�.�b��X[s�&;�A�s�"�:���T����st|��5��^t��2��T��U0�h9�bw��{Ă�����uU�RU��C>R�	��2���������F_���Y.s�2DO'ׂ8���ٳ!t���KD��+��`9�V�f{"���|� `�%�vI�s�+FgY�(	ц;�6�{���G������>S�Fc&��
��φ�ܰ�-u\n_v�j�7umH���W��mJ
�\����T�;ٔȏ=�)�MX��%�n^���F<�{!�����<_wqum�ȹO�0N����d�X���0��򻣹SInL�b�+�Z�/8wj�����}����Q�������%��}D�p>��������Rγ�N�Ƨ�>���#�Ⱥ��Q7w�̹|�=�"�D���kF�׊zwN��ƛF�&{��s�p���5�Ϝ�Y<F\ķ�v��g�>y�����![2-��O��8ʳ*wʤ:�] �K��	�c�TW���;s'7�x����d9�,��2��xBN��^���Z�������p3%��
���Qh�߻Kljb�_G﫦3n��=������`�����^;��N14!��턠M���JQ1Qwpp�Pm�'Zf�W���ܳ�0D�3.:�["�ϗ�g�*U�d�YisΣ�D聓���^j�33��/`�F:��l���?k��F�z�.3�q�enft̮�k!��b�]�wj�Ֆ$�5���G〈��lF�e�;�2���.֤�{3��?S�9���_��O��U�_Z7ӎ�Qc [�1�3;�3���M�Q�u�3�]�^ź���g�R�]��+����Έ(�FwR��)iǋ~>|�Z�>���>8p�|��C��ʜ��n�b� �b�8.g�y���xΏ��:�Es%̹K��e��ܺ�6�_�L����P:1J�듬�C��Gu2T媢��"������xh���1\�sVAR��ߋ���uZm�J���a�]Z!Cx�.�R� �U�O+_t�Ccu�_wRq1�z�hǮ�����@�f�����ݕ�,�������s�7��bb�G&9��n]��q��|�{W�<o�3#
������YHRT����t�3�7bצM�Y��Ư^5k�c���3~[ٗ���g_��&uŅ�X�\0]�r��P��7�������A#�-�Ⱚ���=�^���d6�����"�{+�q6R�sԜ!�"˃d�������,��R�5,���A�c�k�tD9�i���:ٗ�%�&:T0r��N�$���;Z���������ߐXP�d6�v�񭽿c��fO���T�uᘙu�/�.���:H{��~`lm�cͭţ͞�Tv�{��ԩA\�{�pfW�fQ��G�z9�g7gM�T i��7f
1�Y�1����˟S�4�� 1��'Tìˉ=-�W��ɮ�Bκ:��$��{*Dc`��Y/��*�̴��v*�'���=~�o@ fl��m
H<�ԧ��E�s%�S��r�Y�14�cj�#�9ܖ{�;Z}�t�F���1�w�.2<`�فsN�T�4�]4y�nT���'k�@M{�A��<���v���ZR�+37��9�V\���B=r�)<@޻륍���s�uqa:�gQ�����M��'�L[�1V�[5��N�W�Ѻ�"k{3Z��{rd+}}|&u]ǜ��(RT��:����2����Si�:�`����p�b�jΎa�ێ��Yj|�vK
�"r8�j3*u���ǡ,��S�v����*߮��#��Ma���e�ٟ�{�
����Or.�dĉڽ���wY��l�}ˢ�{g8rB�jR�x�U�[�*^��N|�i��Q�6V./b���0�eNȟ�Ҋ�W �r��.���$�ܷ"���h��t6Þ�cv�U��L�<A���
H�Oָe�Z����1r] �fG� I�ܺ���Z'ی� Ic	��&�L����0���f�r��K�%FJ���^��-�����w*��=�-,�Q�0M����Vwx G;���]%*#>	*��<U��*���G	��{�q�U��ƦR�% ��r�"U��.X�U"7�a�#�_���5����Z��ZZ�0Q��}��v@4�d��;�����&������`3Fɚ�@'�1��ϕmN#��c9�3Sܚ�d}�WpR�̺�7�%F0U�(׏]q�JP���
:�p�>��9�z�}&2v�<f����9�D�Y�:T�sW���X�R�qw�꯶�3;\ǲ���	a%�}��u����z(��9�<RAV"��x�ٓ%�R[ss	fBI�j�^PO�bR���뼰�qu��蓔�6\؇%��37��vu�]�sC�'A����;(����T]bO�Nƹ�_!����+�z��˨e��'����
&-��V����MfRӶ�0זL[�k�K0Opw�U5�Q��3�aGb����ڨ�}vf72���w���=>;84������nϘ|��{����MH�N��="���Mf{���Q|����/���Cu9S��xOm�f��q@��A�j�zl�o+��0o]V�1��(�������Bj��D�Ҏ�4_	u�Y.�ǐ�E�����<��j/�@F%����eUa��[��Ey��t�M�ل��ݘ�*fӄ�W+��m݀vׅ̚�k�͈�Y~?��L�\j;�V����Pu�9�����<{��*����c�z{h��O$)�{+Ux�;��yP�l�Ba3>�����N�~�^*�`�&:<�ug�0�yV���;��rG������n���\'.U�8���N�@@������`�.⑝�eeY�1���2�^|w���\J�s�r/ѷ2���D7������}�{U/�:�������T��S��f��U\U֌�I��s0M�G�8N=��z�)����x���.�����͜��t%=�fgitUF�0�K���n���1��<�Ss?L�|\�A6Xb^���|ېj�]��޽���jT�:<:�R�j�q�]�!��l���[�*6��Y�����n�*��ͤ��[.�EI3�^���(`�gjj�6/��
j�;r���������:Y��Ĺ�a�֠r�n�+)�5]��1m��ǩU���%������{�/��(�H���Ĝ����na�T%�F��t�S�;�r���$DT�ZW�aP��R�(1X�,�C3��/xw�6LZ�9�9�;��';�����p��N�.�劗������q�v�8��[9��Ġ��o���4���Ikø�ŉ�5T�[V�p�kA�q�ݭ�Q��l�R�`#^EAucũA
;xw�
N���Xt��u����p9O������k�,#hr�Y:́�������xg1-1=Z�[Z�+��^u�ںu���|ݒ��:��e�0u�+c	#1�'���L�7n�b�7�W�1���՝�
�_H�t%��*)���6-X��1����]ʑXK�wO�ugX�~�t���ؔ�����<��V�kkvZ�V��R�(�f��-U������t�.:��O�s?5��u������P�x)u<T�"f���ܺ%�F��JAn��e^c�bS�`�Y�]�I;���(s�ۺ�8qh��B�c�-'�K��u{@7����/����]�̉�Vc�	�k�RwB�oe^b������<�#m�Mz�*�;"�V�mrTN�1��ɑl�=\[�$;�ړM]dN��{����چ�����Q}���uټ��!Q[7�)h8*��SWPf�C5Y���q ��8cx2�x�뼧D���N��Q�v�9|��o"�у6] z�qblڍ`�j��+P.[iQ��4+f>��Ԛ�ь�z�ν
��V�u�|f�U�ה�r�"�Mˀ�jԣ���\l�We�i��0�,iʄ��=�]�����i�U�FX�<���Ҝ
�(�V'��F�,U��ੑQ~&�{v�K:��c��b\R�k&��v�-���8[ދ��f�%[��Z�N��HԠ�������}v���	�b��n�׻B�ㇹA�Gf+w��ԉJ�;��h�pAXάx��V��H�ux���h<��+-��A�ޘ��:����`#���I�C�Q��}6AMԭ�ub��wj�4I\�׳��󮔤�)�5ڴvM��c�*EŇ΅_eC�^a	n�w������z!99��M}	���y���5��D��d�d=;�{B��\�B3n��ԠZū��]Z��(��SW �ꄮf����}<ٔ�X��Ì��$1��(�_$�uݵ\sĔF��\@nS�ռ�U�g3f�+�Ij"A��_V!N�Qk����U�6��~|��8M�@� -\��i����/���;[����]L:Rs��Eok���sܧ=E��]X�S1�hj�[�w�'��՞�5w-uwT�*
�ӎ�\�������[��u�ݷV��|M}�����\�����׮揯/��Ҹ��go���v�F�޷.7Խ�����.����my,>�	x��}c�#�����H�D+}8��GD��0xť,:�q�"b���:�˚N����[A;q+({�꾼������I�po�o����*�٨�������(�軸:Nc��:��gz�Բn}C.(� �f���0��M<��u�
�M�Rw�	nEõ���=�.P��s5��7
I�����)�U��k����^�t�M�`Ch��s��
V7�j�qU;�����<���ޚ��`�T#��xVL���|��ڟG��[��P�u�SN��у�y�H�j�fm
<�"
ێ����WV��_�<�M=�`��k�E�>)E{�Ӝ8��:T�q����:��U��tj}���zT�	�L��$�U��[��S�y|�5�������ԁ�A�W��؟��|j[cֲ�?x��V��@t�gA�m,����z�b�2r=U 	5��l�LQ��W%�,�ڻ��5��	���=�����E��`���p�Z#īƺ&����j9j�NS2��/6��0mM� ��H�$����tt�YO��5�v{ ����ʱ:��+�I�d<��j�*���b�<����:)�����H�}���&m��|�ƕ�����u�ڲJ�#�/ﾆ+qM�Y.�M/p�c�*X�3�{��8Y�1�Ot�UKwg� m���_Q����3���t����gp��G��G�6���e���t�b��R��8�y��A��OϨu�̊)f[���"䴽1^����Ҵ��)�O(����]ub��u�4�+W��X���I�����A}�j-�b+�o�k�owZ̉`Ǩ�^�sj;ܶ��?�}��ʟw�&�Q+�6�ma���͋�5x��!M�+�n�k載2j�e�|�U�����7�=
�uDS��˽F�0��N�w�y|}��0�~�~0\����&������գS��S�
k|h�]�8��@d��W�i��}=��Xn5������?�M}�σ�Mمx�i hEo����/3�٤�խ�����6/�@}�<=��JXU��=�` F'	"eSI^�8>�X�b;>�m�n�m@�L
葛���M��^�)C��ɢ��<d]��s��;�]��7�bS�otf.%7�3��f��g���E͛� ��jU
�����)�f�*η�<7�o�c�u�����$��>P%�}�R�/`���wM�<Օ]Leu,���+��Z���z�Z�Q��5V�#��=�N��\��m��9;uU���}zVt㠬�"1�17�%��Hɗ�!Hs���@�Fed)��Fܩ6�_��È=}���7~�䳢�nz=�V`/j�Y�H]A���0~ւ�C�`%F��8�w>W��
��g��Ǯ���e�o�&�����Cu��Goc����;�e3
���0et<re�Y��_��n�8�a*D�?��9�vQ|o�N��c;`�r�V�Z'�r�)��[g��|��#�n[�z�{�Y�n9��o���î��ʚ���c�<O�}�&��<�(�ȝ徫����<)��I�i��e`A�U�.��������k�^�Pyq7�]�[��>�h�Ɏژ1�|�Fݬ����ց�WM;�8ץ��P��������t��ʺ?U�f�B���Qgn���j*��7�I\�W�c�jn,LU��V�ڤ;n�=�`��W0�Щ��������}+pۙ�Nq##�3��Ū�]VUWֽ�ӏ��^ʳt߲��e�=�`��|2^w�)�8"}��j�8N��w�z�~���0�^�tt��Sw�����zp�F}U�7{
)�
M��~
�0X�a�t\�umL����"�������,ϧ� �J�3F�i�x7��R��E?��Pc[��g.hyڔhb��DR�i�buvա\���W���O�t�������V�YKU�yr�����o-ص��;�]�K;acd�x9���0���Vb�!W���꧹�9+�b��TNt/��e�+v�����6����3oĩ`���^����ǽ��F8��&����z���@g�8J3�'!T\΅a��<8�������b��{��	�RZ�]?Ϩ�S�k��u	1qi��h��ؼM�p9ոL���n\P��+h��Ms��G�,_���_}IS�Vb���g6��a�CY]Xc�B�	_(����粜M�tR�9���%�\%��u�Xm��P
�h���s�G�\���5P�`�g�����`�9ܞ�{/�	�n.w���^ˣ���e���X Ji���=Sq�c�b\A��j=%3����Ƀj���Ϟ�X��o����뷈S���2Θ�k���M>�k�ּW�"ȿ-8+�x��X��B��sqW'5�����Ӯ�x�v�<EN(G��'�����jN��5d1f���y=!ㆽ��h��}J�v���rR�3�ȣ�'�t!�޻��g���X��W�t�:�;������~��w�s������"�S�ss��7����[�	���"����;L�At����dm��n����+���d��<�����G��O���§5S{���jo�,�v+���;$j�N�ɅB�6A�ڭQf�RAʊ��"_.�=�3�tn���bmuv뇇 j�9�^Tpn���{�_uŔ.�w�:o\zE���&%�����"�N�7��������!-��J��U�����D�j�uK]\X̵Vx�s��u�lفr��~�����@�pԽ��w���;5�~/��nY���'Y캾����?	~�
��Tk�A��Xr7}�ȶ��{� ���sU����p��G��=�-�^J����k`[��֙�QS���6az��}X��Y�r�ܮ�?��S�RN]zn(�?���w�_4�=��a9�v�#J�>�U]�csBE�4##�V]�M��:��{��Rz1F�e$�E��8(�ѧr$_�N򜡕s���f&;T�3-KiLɍ��'gm��$�D��N�/�����ٙs�_F	��azN����)'�7=a��2�^�h�uc��XS��[�3�W_'�r51���GҍdU�l]�Æ�پʞ�:�x���f�P�s���d�~���&߶�1����$|�N�R�E�I�0H�ӵ'/���r�g�6��������P�[��*��0"���e�K$,��y��4�lD��o�r<wJ7�w,���L� i�2a�Mk�6�,�l_?\Mq3+z����6K�f~#b{ա�Eb��`��G�b�6։#Gr��
������Fw~jV=�ݼtg���*���� ���E�$�d���3a��:�;�z��i�8庛5�uӤ��~��J4�`�u�()t�U�;]��D�o5Y1����ͥ���8ly�yn�]�e�:�g��0�N��,�\2����׾`����Gp��D�בr4aDQw���2ڔ>���D+J_�x�#+���tBޗ^����v령|���}���u��iA����| ���l�HI�.��s��4��a����{�اz�
�Y���d#r3.�vjrR</�]z|>]:�W�]�Y��MGX������\e�#�G�V�]�w��P�:u:�^w��-�J 	�&�?k�6�>M��.��;{]���ʚ��ɨ̯!��PzE�ӌ�z0���*� ����!��>��:}!�'��_O �	�5sV�U��C��U�J�bm(��hJN܂]�ճL���Np�o�w"�D���}=+gOL���v���C��˨4-R���l�yB$ۻ�t�Z,�7j]ZY\�U���mW{���O�z��޳Ї�B��qy/�l�*ry��+)C3��W��,8}�S�C��|O���,�Ҽ�����5f��/J�'�'��㶽CT�HxBC�m�U<yn�W�ɇb}�<�D��˂���6�N�
�� �G<Y�8M�wA6�*j�u8���OrS5n��v^Kq\v���ݳ�Xԅ�����{��N�,���g{[���&��wm�8�zy�Imv6o^0l�]P���v�@:��Nٜ�0�a|��&0g[�9%�m��H�3�]mދW���#,��{½�۴��O=��g��(�+GE#�t�wM8�boٵ����x-߻��?|����v��r�Zٜ[��9y�N)���B�=Ց] d�P��\�N}:�@u�����R� ���K1��K*SU�s��.���BX�qq!mk�%��tP�Ոs���'����<g|���Gt��P��j�|�}|~��󧤞�{d"Egv�n|�� psXD�|kט+ύ�Jc��9=P���Wh}���w}�1��6��WN�}hz@b뮡����v9ё4��Ux���O���Ğ�����ar�5*�>u���| �Գ��Z}�Y������U�Պ�wT�&�ݪP�L+ @����y���!Y�	�o��E	��<��Z2���d�`�e�g��毽&�3j6��0���So�O&z�\�ܮ�5�(i����U�^�[ز_�|B�0���}���[2�Y��U�܇���]:}��B�Iw���<.�G�O�e�6_c�n��c�)��m���R�R���:n(�f�9�G8�ר�1<=�\�>QS�o��.�W��}�ǱX��"�M�B�}���FK�&[�;7���F�;k6�o ka���+�sY���M[k�X�)�0��*U�;���z���YЁ�JC���$߯1����:�5W��]ټ��Y{���j�����7��ڵx%�Qc�շO����k��КlO����S�:U�ͣ�~�:3�^�u>k�yns��vH>
,;R��
�]{��9wy��ITO�6���j��D��g���>ػ���%t��z/���^j���37�<��Q����#��/"j��]��Zu<�3��6�9�u\�s�(F#��B�hDtS[	m�Ǒ��%����ُ�p�H��5��g�
]�:^�.%��3	Ly�����q#�^h=����
���°]�X�!��7�VH�O�(Y��v�jET�uu�o�#�F".�v�:OEoQO������	�6"G�[��{���7�ƋSL���#���B�k�7����D���í�O�$J���V��{�e��=���!�Мm�|;pmq��>������|�tl��U��q��H��Y"��+-�><׵Պ�3+#�Ao�F:�-�OV��@�qi�z�����ˍ� Z11�޺�]SѷlI���#�M&����.p�����[*�ܾ� �-��G��<5aCOك�V��0�h�B���ޮB�$����N$�lI�w��"}xO��F3´����yj>���vk��Ӹ�D�:��y&\�g�P��I�������ݶ��i��0���ph���A�&�v�q�����e�6�����@�.�{83{ݷ��,�Q����P�h��k����p����k��+��V��-�������
��[�>n����P�{j!ۏ���g�=����Yt�8`Y�X���c�'������dOCp��O�j�|l�ܰx'OZ�`y������Jʌ�=h�bq
�}@�F�͟9�V`g�}F���֩�b^a�b7S�2D���+�q�.�WOk����on��z�z����:g@n��6:���=̟p^ɄDd�y�|r&��Fx����o�Xb˫!g/�(����F��)]��5���t<��ŏ.��;Ry�ڹC(�m�s{�jy����J��/^�s���b�_�����09�T.<�կz6~��4R~U+X�}�I�5�,�rg�bN�l����)⻡쭡F�'<.�;�k�b��'U�z6�3
�\ׅ��7Q�b����v����T(��1nF������;bNL8���)��Y��^IC鋗���/s�����\=��6�������˺��o>����}ʚ4�����۹�m�>bm7�s�wj�^�kا/�ԩ}O�lƽ���,S�R5H�<.r��]��,�y,V)T�h=T	QHZCj��>~`�Kh�F�x��ȭg���p�&gPʷ�4D�6Γ����v�seCj�T�jSW�8�3n��y��ѭʳ�J�}�B'�+�ٜk�C6N��3��n��7�Z
�Voa�F�n�NG��ə��Z�8�#�mɓ`jsU��Q��U��WhXF5��G���`�G1f��Ƅ�MC�g%�z6/$z�j�DS���m��R�O�F� ���W�m\J��M�q�P��.��A�-�_3t�NG�����&n-r�{�<��Y����;<���.\	P{ ��a��{����5����Hu�Ğ<̔:;�9kա�xf�9V�7�Q�T�Wċ��)�J���{��r]��i�$�2Dϝە�O)�}��3\f�HM�.S��7�5���0��1�(<�gԌ�Ѣӵ��L��X1�!���[�G3�˂��w@�^p��^�M1���ŝ��1R�Z�F��o��
H*+�Y�(������}�k�˻vM7BJN�/yTMG,��b�Fy}0V܄��^apn������@Հ��}��y,���r����sW�|������V�t}gF5q+�{ER�o�pO�G�'��y�.��N�Fn�Z�:ɣX`��n�@~)^�K���)f��9�g�������da��,�xu��b1���ҍܸ]OLR�,� 7"e�[�-��04>y�r�p\�dK�࿩z�l�$�^�P��"�-&�~ ��Vǋw��3hv�����������M����8�š�f6�G�X\N��v����{�Ck���U���iޭVq;��k,u�Q[�� �Q�Bf�_~6��/yp���[�<U�f*x��j���uԭ��o9�Pգ)t�2i�Z�$�|�w:���%���
ÿ��Q��y��"h�{C�1u�gf���St��<#Y(��V�1��.ݩ9��QK�8���@q�L79L��;j��:.�Δ����;zk�Z��*	|8�tP�;f�z8۽�vx�8���&����2!�@G�	��ͫ��9>��㴵����+�o{.��Zib�=7+�}(���wA� �e��,�GhYְй�����e�V�[3�Ҩ�r��I.˦��W�i`T��J�X���H��;�r]Fb���n�Gwf��
^���NT�-�ӕ^v�%lQ9/5t�!,b�����[|)]��gjE���4��G�q�M|΄�l�x?:�2�
��H�|hWb�T� �r�6яi<Ԩ�]CK��6�]0��x2��lP�R�v�?s�&��i�+���jHV�Wn�ĐZ�ک����Q�b[Y�ژ2���ʊb&^ڧ{j
�R�`�г:qh�h�J�`\��l�u�+�p���R�����Xݥ�GSmӤ:WvVn���� ��J�^i$���_a���o����}An~uzt�'���R��!WH��(Z�Ӥ���G�3��;�VôR����U�i�}��c=Rl�3�����)����v�ݷ�'-ZMˣJܲ�wE�"U���VL�]-1F��y�n�W|s����MZ{���-8�V�$��ͬ7/k� �dt���]��4�V�3�+L���PnI~ۻ����1j0%����ڛS+=K����WM�/c����E��Y�ǃձ̬Һ��9��kV���嫞 �� Q��tHK�X.�q����i��]gi���;���e�7;�:����[��������p�w�bLY�A�v{���N3�lqg��zi^U��]�7�>q�ېL}peț4�2UҠa�n�Cs�F�@�IM*�:;ok����PE{YB>������^�J��V��k5��[|�b�ͭ����Ӓ�iС�.��#�-�qN��yu�q;�h�	��:��`v��f����i78��+������9�a%�vl��]i���'uՉe-�π;�����O3��vm��F펒�YS�N��t��M� �ݦB2��vl�1��O�)�{���l0���:�鰉�����s��[,L����O�ޮ�n�7�å*�nǣb�J���Ff;�=5r�M��7��
�,�I��ղ��]ol�=�d�����.�*ˬ���X�F따&��y�H2���L�	#���\C[/�]2v�,�7}���RG7�e�H~��=�L�:�Zq6��ۮ�;w������[�QdW���Id�������f�.N�J���F����W��2=�\���/M�u����A�}*_�Ǔ��Z�3D4�PQVK��f���1~�����Ç�+�L�&+R3:�Y�ė �[8�M2FlO�R���i��am�g.���n5{w��\݁�y�A�q��8�9c~�Ü�s�� �y���!K6��j�{��~ʰ�>N��㟾�7���)+�5~���Q	�~k��WԺ;�k�cv����������vʝ1��_�hx��i�KQ�����`#�]�~��vy���̛�d;B{/�=VJ~��(����mV(|&L�)��\5�t���{���9�"�����Og��I5���K.�ug��L��|�ڻ��˧�5�}���0��=�/�%Y���^�-�(V���}�l1�����ýgWq*(C���=xo[���d��`i�>�NV�|�鉕���y:���{8��˟Q�c�ou�n�`�綫�Κ.5�Y�|�ʦD	���Y���x'�]��'���f�Teq����uw��5��E��:d-���D�_i}8�BJ*���V��5noef��K�W|,��ouI����*���2�f4��2�����BԮ�BƜ�!1������C���:9��(�^ż����i$%ٮ���y�'B����o?9i��S����'M8�$������[�������>	]���|����xuM*��}��Np
�-&�+����Π�W{�gJ��Ы
q�ؾ�7����ji�v[�7�c��7�ڇ�pc _�U�G�Ξ��W�����W���8A^٢1ڑ��9o|t�����h̺��y��X�ݠ~�7a��!�S�GAcj��vc'йS����jWud���p�BT��~p�7
�V�m�VGW��T�c4>��o�L�{Z�Tk=2��S�XnCh��9gz�6o��g�B�_�٠����m˸���/pG��j�F�>��E��bFm���ѵ$n��Mq)/�1�3�,����,K����ʫ��݊߇g�\g<Zܥ+G
b�I��.l�M���h����3B �9��g�2{����.�pvaD�[:D��s;5Ob<�.h�E��^�k��(	�/%T{� Y�輬Ԝ��+�y��(���0gT�-��$]i������M�(0�k�n�&���?��۪;.�	��wavԴN������>�>��%�>E`E�Ae���Ugv�%7V�V�����Z�����d�L����*��/����X�'^��p;�W,����ύ�a-���+�6��Z�)uFtb����ؗ��
sgs{���Â�p�T�0��o�.�ה��ں��ᴕ-�]J�d��<9v�ut����g!���1���$uqL[@����G��'�:{z����j�1>�!Ot���<]څ$z�����yOP��`�^��g�+��9�PB2��e^�z�·2���ا�~3�U0�5a�Y���R�>/��}�G]ܯ���Q�o�Z�[+2���[�p]�;Wګ�]I��>Dx��P�$6����ul��g�_b����L��7��ڹ^��5<�b�sj\���9<�r��ûn �n7�D\�J��)R+��OR̪�LD�L��_�Az���Ӻ�	��©p��sڜ=~����u�y_2i��b�{ysLxjU߆g�/��KB}�T��)x���j�8�$D��>�b�p�}sq��Yڞ����W��2�lg/;�k�9�X�o�2�i0h]{٥���;����d�2{;uLj�+�IK���iL�Wh֦l��e�P�]\݂Wr�:�_J�b}����h2��������s��Y/�ze�cW˫%B���LeM��*s��dH��W˞+��
A%:O�A״,�i�+��������:�	�˭��ml�9b<��V�fU��ǩ��j�� �]�39p;*�G���t��wh&N;l�?G|V"Wʂ9+��T�ٖjq�o��dm�(���3Y1iv�Իu��	V�VY}�H`��Q�K5�Yɷ��"nsY*�E'�.E�i���Q�W��[�E�WJ���~�RxA�ݍ3YҢ�90:���˖�9��'��ȊQ����lFΞu>"����$P�mv�鸺Mv�fp�K�Õ&V�^�)Zͧ.�׹YN���w"-ng7�Kqp}t[�8{+ey>��Ls(HO]��՛f��<ȉ�8b�|=���Fs�,cs����U��yp��.ś�t�@�`�?	u���M����{3;��r����p5J���M>s=NU��~G��ĩ�/Ӥ9߄���N�b�_2;d���e�WGن��q���̿���������~�Kp�Wn��2�`��_��I��p�3�������'�b;�$��:�9Fw����/[&cwHa�G+墔�Q��=z��o���{̜���Y]��Ď�����d�Hq�PR��0��/��ϙ�ö+��	���<��Jؙ<8/F�W��vb���~-�"���Zj(|SR�T��ĩ�/�m�?yu�Q9�㒂UZ�72܊��,>DI���V/:8=�l�V5�Xf/:��%�}��ؐ>����9��ͫ�HV�7�
T]xY�}r�+h��k��]��ͻh�� �c������'d���H�8�Q��4Z��fN�z��X���f�lv���m��:�m+���J�[��`��hU�v�Z�LS)��������ԻK��SZ+�{5|��Ϛ���_�q緱���`z:�����<s#���fV���Z��7Y�[��_t��}�z�ң+���1a��׀U֑
������V���w�^NqQs�J�!SĕV��a��۰�yP2z灉�Эtdd���n����[�QA��q8���غۄj�j�.�"qy�}�4�8����~��/A�������0�/|���@���0��1^Q��I;��:Df��JZ˪(��)��Ce\a�V���n�\���YO���$sܔgooB��`�_/W%1�b�7:�QT�q��usB�f������:�D����oy9����
9^�T�>�!&TSM�;�R.A�R�)��"�^���9�'�5s2O��*��9�u-1�UES�5������3C��h�馊�wǧ,鋍.8ѷq'}z)z�U�߉q���ày՗Lk5��H�(׶�x�V����K�u��[��젮^���u�;�����*KϰfQ��my�u��F���_�Ӌ����#5�c����zA�1��VFCǙ�Rvw��~��[��I)T�kk!}�Hsu���u��J�5P�BL�cWt#�WA�M%J~	#��DP�yS��v�PC����{$�h���L⸷����U�� ��;�-��Έ �x!U��"�轫��<*��M���Y�M#K����꜓^�ݻn�Nibl��]�5�ǔ/_�3}=X�����N�t���<����!Q�9Yy?>���҈��w�⵸�g�0:�g�<�>5.[��]Ojȸ�����]��N���
ggjy^�����X���e��G�E��QX��*���*�;ơ�vnN�3��Em�8]�2��Ǹq�mV�)�P!a�7Q>T2I>�Z�0t��g��;P@�s��y�S����5�<B�������;v%**<�sr�T�Q�%]�qB�[Uc���Ϧ��,aB(��(Թ�����c�W��)0��dT�_w�8���z��1-�!ܠ�x�ǽX����=$�,��#�:�@�ʖD �)n���M`����O.ә��>
���_��軇�j�����J˽ɽ�\�Q7p�G;���t^�*��{&�z��B�ʙ�]K͟�&O`��7�����^�Pe@����X��H7�6�v0oY�fl��L�f?v�a����F����ԳϤ�ٔo����1|=M�<W�m������l���x;`s��l�ٱ�Q���hn!T}n�ܨ�7|i�V�˨�#;��CfmcX�Wd���_q�L�MFӸ�XAcγc"���킷{1
ν�d�8Ps9ܶ�e#}�i�+ܾ��f�M�J���VQ��l�B�'�So�jեm��ѧy��E&��'+�qr�S/v�'�z���m>3�9��~?L��սDD�+G{Έ�R♉�6j
>��w����H���N�>љ>�������zE���3z�n�~��}?]]�)Y���և��j���٢���c�(��k@M-<������Tq����jG4Ӭ�p|�z����hx����yl6"x�A����PZ��Gg�Iyv�T[o���i���ɭq�σ~ء�L��E=��L�h��Y���m�S�f�~�����m�_LF,�z�,��G�r�2���񨳹q1�?2�^	����q�4:%í�5�o�LQ�&k��%����c�r��W`�5}�gɥ��i��6~�1ʗ{ L*g� ��(����'F�w3��ѱ�eX���4^���2_��J4�p�m$�mF�*�i���Yů����c8ڧkU>&�=�P�<�T�-���Ӗ�V���S�q���
�c���¾&{ʯZT$ı���˅��/�M���s��Pz}���o�T{��)���)œ��|�>��sD.����>�<]s�[�g0X��הvf*S홡�e��
V�S�9�ޗ�\7HP+��f�� ��j2Z��Sc�h���K���@n1y��՗7;5�J���2	�	bs�o3tg}:�f���Yt�l��WO�m���V��Ձ�>�h0�>���m�C�՞r�nsyA@M��O�p]�r���:��U��;j�i�Ur�*E�w��ۊr�����+�s9�K���\�ݨ��,.{$�<' ��jq]��oX{�C޳r�e��#�ѩf���ȹqU
�n��5���}�Յ���/��q�k���va��K�<�o�%��@���C��)�me*X�� .C���_�t�׶.���=�L��:G�����_�ܳ&F�p���}RьQ��`����o��uKӓY^6=$k��Jr��S��|��,[Z�t,=�x�_a����V�H�������G�"j����^�DV�I�|(7H�q�������TnmŞ���\�zez�Bۖ�����ʋ7�5��ΚB��Lj�d�`fQٞ���t�]��#Q�o��Q�-�^`�G+hwN� ��ʤkx���w#��x�+�>^��S���stN�{��!'J:��M\�ъy`�>�nL�M�'�\�K ���]�g���j����ݐ\9����3#�z��d�=���9�M�<�khlɃ {V+�>'=r�����2�]6^ҟ�lfۙ��qz�o����ja����u��p�y���Rg��/�\��������U����|�ъ��]fJ7յ�̰q�Qڥ%/֎���R)�(i����&���ju��X/��3a��� �ý}���.�
8��c7k�=V��'�Y�ю���%���<n��}{��ɹ��v���g����-��v���F���TWU�v��1z�� (���>���F��9-F�ջfg��rb[�h����;���q8K��p%h��lA���bd�@B�1�e
� �'ӯ�j�4/R��ˎZ���`�b�ʷ�+�8�T����ZR����֥�U�A{R_�����^��,�;a�L\̷�e���yX��D[���8b�N�� ����]8��}��r>�mx���=����ס^���t�jDr˚���} Я(��x�'A�>x�-��_"{���^y��47��/�Ĵkoj�B��:>�t���9������cοc�Ɣ�<���O^�s"-}���xfM��^���&�꜐��1s��#G�m�R��q��[^�!���K��n�Xg+��u9�tY���x��0;o޳�����[��'�����Q��TRM�.ծ�핪�}��4�q�\�b�1fEL^���&=��[���w���SȽ(��xF{-��on�X[�����7YJ��~}]N���U�����@���~���[ۥ1���W��32�ٓ���pgC�q�ݷ|w-t�F@-�Q��񻷈`����P�:�N����yb�C�ZR]�e�]p8S�9�Nؗ+�meōZ�u�Ԟn�t{&�@��!�\��ɿ��
mv>��-�w��"��.�zygT�Y{X�]j�	�z=Vqx!��X��t�k&7�����|�q��eW���W�=C�{���N��;��Y)�y�!x=��E����,�Z�-��}f'N0���͍�F��zp�pV�ev3��PV��@�͡��|�mִ>��ώ�VL������U��H�{&t�2���'R�4CQ���]Pz%��N��}�������-�닰�ub-M21����ޏ��~�V�#���6�{���TD��3���f�˿�D�;9޶����)��A�6���IQfc��dN�߄��ګ���ZĈ�20f3��"�TwX�����wJ���OهY5C�f�M_��'�SҹNc��+=�<;[�W|���1z��l�i1��4��A~���N�f��ަ$���+�݀���.2�.��N轖����o���^�L��q���DeZ��#)ƛ帣�F�U�>�ŭ��]��j�hrQ��S��l����F���N�N'�<�N0��2�N�>�0�	!J��y�Mxޛ����o^��}�E��/O��O�UWX� ���*��e�yȺl6�G�����uʂ<��{�� �Q:z{���ҫ��gru��RV�Ug�E%e]����J�Z���l=��-S왳��Q\kh*{�[(���[��:ͮ$���s�V�p��[�-��fr�ր�k��?رU�Z��M_vWI��u�y�;�oP��������������url~�Dmв��ؔ@n7M���o$�nm���]#Wqk:u2��י�;�5ܹEre3Vo
۽�B�kj��IKx��إl��9)�j\;���X�5Cv��Q[@��a����\��d�����=KA��/vƧm��-�P˾����ô�9�5db����v�]`����]�9:��-��U�`����Lͫ���[}�V�432:���yŅ�ܛ�$E��D�+��[mv�&����l��Ӫ��Z�L���أA�CxD��),/���K�љ�v[4ݻպM�a��V�`o���f*��`�Һ����ɓas6���oM��Y���݊��͵�K���K�ky��3�e����ih"�]Ե��gUܭgSb����\�2Q�v�*:;\k��
���[L]�����N�|�׻�bރ��9Vb���cvˮ��6��tY�x�#�A��h��D�E�wܕ�󹉥�̇l�t=�a�`�O[z0m�Ĺ��#c㿊2�W���(e��2��wme8��}$��$��0)�a���[�S���ě�u�H�J6���y�?�)�(9Nf��$p��X�,D�l{��h�����f�3�r��r�*�A1�Ew_@��b9�ЗO9�j�"0�U�(���g!6v3���#j�g_t����r���;[�&�P���u�bkg%{�L��eu�շz�}c+^��5�Z��tbWjAY��qh�3�^��2�WrͺaF�j㹻�wrp���"�ӻ��b�l�ڛѮs��I�f�P�/�,�A�����=wٝ�f�W΄����r�IopZ�u�3&�/Q�ڭZ�9!&�;��^.�:�O�W��{7F�7��n�FZE�;�N&Wa�E��`�a�H�n.�X*���],�L{��q���w���6;�W�R�M�� ���k�#uѡ��f�C]�\�~��:WJ�{�+v�n7�:��.v��3���)�*���b�����ָq9֘��U%eb�7H��;]�ǣy��V\鴓����e�9����XU&6N�W����`��y�1+��71�*v�1U�P��^�z���u�����v3���MjQ�H�[��Yc� ��GP��:($��M��h�	�?�n>��VuM�j�u�ЗE.˚0��}.v�m�;�n//%(	߽���;J�X�F�Z�4[�jp���W*��@�\� ���]���M�l9�͵�[�}6ն
�y�6��$+u� �]h��ͫ�������f�)
��f�R�0"��6q?�:ys�J*6B��3}{Ӷ]pGJ��Yw(���J>����7�󸪬�ث��e�Ψ8�ܴGb����o�:�|��ɺ~�h�6��sQ�j.�Dz#�dA�Z���\(Ol;*7ޮN`6vk��,�zOь/\�^�����wv^u���A�]M��p�*9�Tt�Qp��\��zqm
>�K��%l�d<̼|�oy���f���o�2:_2�,Cπ�]1�a�R��eU���a�~jh	�}�u�/;s{�����NP3�4L��^�o^e�H��}�:��|+]��;V3��1W�D-![ewk>Kse��8���aK�]Ǭd�ӣ����.� �� ��`j�����6�Bb�/NNڟdy���H��t��̸���R�.���2uuǖ)�7�&{�$B.��Ïw��O�۷����u������ý;:����z:�:�X1`��ᗎ�����:�眾CenOI�W�9��
��~�EBK������'R�\�EF0U;]T(-���g���E_�}��0���T��"C�3r�����\��UHu��yFC�jz�|�5��4��Lv^��H���?[#A !��0u�Kr�^vE���O�h�{Vy)Z�45o7�)�o��_nn��:a�'�wO��vW~�\Y�^ne��u:�g3���A8�]�}�Nv�k9��fe3�:�n->���g1p
��hn﷖i�����~qg��꿏�`���1�Go��8a({)�O�&!�.A�\�P�*T۽�WY�/*;��
��补��ߠ�)=���8/�����Ǔ�[��@�N��е}�8�����dS�w*��;���\od�ȷ50{8����xX ;��/NTݫ���zh��}��v	s�s{��x�W�A�s�������Nfhgl��E�M\2x��z{}�ѓ�Ck�~�ɾ��n�
���T
F�,����=�nX1]ּy���x�a���{n���6 ;��<�ܱb�ib_��YɆ�U��G����w��PbT��*Wf(͹���2�Z�z=8�5f+rj, <�q0��#�h	��pzD�h!7t_��?o�b~�Q�#�[��=9/�n}���Y��Wn������x�O[�e���[캞�����w�rJ{"�aCx���qkc4t7k�8~o}����������V3�/֑{��߳���pqv0|�)}�X�$O{l(3+_z�D]߮�GE���Sx�WlH��N�pf7=�`s+�"5O�l�G�)kǪ�1���EZD��{ia��H���=�O� �ͳ�Z�;-��i��z�u��YR�yIC�89p�w[�eJ��0�a�)������m?�2;�����5�7�5�>b>:q��躽=Dv0��Lk�kw	�&M�7��C�������;r:&nh��CH;�4��~����5z3&����x�`U��c�+L�W��2�����4����������X��*��P�;���GM��3_+�[�v�:�G~�����X����&�>~��NO���i1ǝj���oQРBb�8A����ӧts��
>���Z�[/�N�w�l�����3��ݞKe�PkϱP���s�ls"+�����y���0c	
}�&�T��m��X�b��ŝbbg�U/+|�rNn��5�ڶDv�s�����T{����.�tb2ޏ��z
�q�wvx��>�h�**~�KĬ7h�;S��jN�˅-�F<o�5&%�^�^��X\�3&�%RZ�*��7=S�K�lȭD��f3*�NO��j�%fux;r��v���>�`��ӷ�f�sO�U��ǒ@��51f�P�0��֏{%�o�`�r��q݋�S- �{~�$*��]7	��^�3T+�Z����Yz�;1�
�C&'W���/C"Xϴo������4�
"9��OF�����\�S;�X��X݈(����bOgnEk7�}ӡ�� ̖��Z���=��6��yGu�S:��iJŬ��:m����$S�:���F*���.=W�:T�Cfӏ��F�,��I�{�$���^G��7s�{:�	�Ŗæ�`\12�'�P"+ Ѯ�c��:�]\��;s����so��S;��H�77M�>u�g�*P�����V��e�0�Mّ�v���˟>�H�̈�����Ï�Ә�k�kE]d�mF��o��".Z����>���&�^Aم��'�7�2R��0D�����;J}���l^�4�v�'�����$�ETa��� �\{I�����=�L��`:�Η�Ld�^F�HuQs];�oɯ'�U���;�����Յ�睶;oj�ÅOb��=���a��@z\]��F����پB�X*~���*�#}�����v5}�n����������|.�S$hUYf���u���;��t��+E8��1��Vng��}Egh�9�耳��i�V6Ώ,�qӆ�m�2'��ڑ��dCޔUV	&�̿I�T끃~���FX�П�p�{�o��E�U���G/6���*k-ŤV_@ܫQ�a��2�S����D^žyYF�~F��n�Z�uNc�<�"}V!��OxE�^��^h��ƾTP >��z�xUB�Eʟnq�7]p�SB�c"��}���FY>��G�\&��Ҭ5}n�F*�� ����~�y���m�q吒^6���jn>�9\���q�FƷ�,��K+���\v��%'J9��WC�p���� ���wy��p���-yo�_��^���SHVs���7D��gn�\ӻ]A��@�6����M^#!թv~���ո�����w��s#�d���s��bg�,N���V����ww|as����!(�����#3�M�ٞ�>��9����xnNc~��ٳ�!S��w��m��t�H�W�������jp;�S�R̘�y�鼆s�;��f�U�9���;���ه���v�/���p�a��ޭ�EU��x�Q9�f��:f_�]�S�i�e"�+M���1=Ө�q�WyV�T|$I�$�C���"TG1^G<��xo��w��To�Z]��Mc�̬־��^蟔�tD�����De.��ݾT��e��|��]9�o��&kr*�bgxU�㮴y����ݏ��j���I߶�e�?p����]OE w-���Ƽ��H;T��=G@��I�f�8��ϔlƍ������i��P�n^�<�����6]���Cvk�F`}K`9O���㪶c1�+�[����Y�_U2,,��p{ְ8=�=vaG�n��_`���O��dA�k��-�{�(@U��m��uB��ǩ�j1�/eM�n	j�{8�v�{�:h��3w ����j����q�����q�tlZ2녷��k�z7��-~�a�vm�����񧏸��Z/��Vz�����-�h��V��G���rl�Q[�;n��eb%9��ͱ�oL�X;-t��u��5]2D�{�_Ln���^�6�n/��[�W�b�[W�����`|G
̯y{��R�����s{cp���%'��ЎlO��]�Yn���Cŷ�܆������=f_���;�
OV���Sy��X�Э1w�#�bl�̉��^)_{���D�P:S�$O������34ǫ�.�����u�ۋ�	���e�,��8s�ܭ�Q�0��j.���H`��y�;/���b/�ϔL�9��O��TP���U��(�jaX�m@!\���U�`�WWb���tz=+�g�}��(�zC�FOK�7��@�G��~zV��~20�DF�߭ո�z���F�WX��3���G+��� �(w��_S2{�7'��S���up�HI���99�a/D��{��CT��Q�0U�{ݾ��sQ�뺼y5j���F�_�]qz��ϳbwT�I�����(B���x�(��~"�6#ًf�}��YC+r�´���ʫ��[�|��o��)�À�\��s�]|^��-s6�ýU
Ѥ��z0(�s������_���/.��RYo������	�^�[�v��I�����%�õ!I�u�~ۭ5���ky%��E�U��������{�]nu�B�nA����noT�䦫�)'r���a�h;���Z�B�9.xw�wK����ũ�R�� �u^�1H��wʵ���7�`:�巘��gf�ug�͌�OL�'���Qŕ��Z��5�6Q)��y�3��7���U���D��u@Ѩ{]jeŏ��5缳���y�{(z�����r!��Z�h�5�EQx3p�֊k]m�zb��g2�0��_�I���iB�����:���L�Yz������BW����s��\��4�~�B+#du>NgB����ݧj'��ԫ-�q�Y��34�����@���_b�sի4��(z�1�4v[KhE��3a��ʋ��������x��A�3O��T2G?|��y��TUqYy/�񹪈��o���<��pr�"���Aždŗ�b�|���[wG���K��.5@c�z�ʛ�ӣ�h�Ӊ?�i�s����cj��E��Eև�=u�IK��W��j
�f��Y�Ex�wU�����֕}͸�h~{�H���o�M4Boɡ�)4d��tu����ʪ�g�e�h�<:�m+���}�a������\�7����±�~�R�^��;���c�J���n����+-�{R�=7b��dd�J����2Z�Z�����Њ�����9�n5��h��4�Gr>�P%�mL�yJ*�+�z�w]�tQv3X^'%�n��\�î��hs��4�d��U����ՂVQ�I�N�6��q�U�����׊��z����9�]r�.�`��	v탾���-g!>'gF�Ķz#��4["2	�����<�yǍG���۔�a*��No�w�����3s��Mf�m�PS4U\Ǎ����ð<Q`�ŗƐ���������&��K�wX�YAO���_�~ߟ%��D)����9�.��pT��W��^X=��w��N)�$w���΃-T�/�yc�Z�䮵{G:x��^zW��:5�KH�ǘ��dS�����Od������S���O.-ujE�M��1��h-�Wx����{�����v�#Uu<Q\8�����>��x9\���n�a����Sb3��qbi$/�,��Q0R��}U�N���>�L� is��9,A�#�s���~��o�Y��"�#}c_�t�Q X��\G����Pe���{`�֥D��7dg�Α���jD�C�K���[����F���⟇`e��\kgУ��\t� �l�wrX�+�Hҭ���݅�"=��9'v���]Q]}�eJ��ã�u*I��<��Խ"�З�n�v����~S���h��"�݊���P��=n0�H�r��Vf�w9�Run�N�¾�.n�T�\e�TW$�ak#�GKyÛ��\a
���\��<y�v#G��m�Mm7g.��t�57ku�dI��K����dW\μJ�=�c{���ە8dM��dzK��:@?3^v)��0/5�fG���W�ާ��Ӫ�o�<�X{�,��]l�f�{�v\�q�N}9dm9Hy;t-�����s3�ȃiG`J�h~�ǫ+��6e���'h�E���S*��^ž�GE�3O�C�ö�:m���2��s��U�᝽�[Yt�|凐�k���?*c������'Zc�u*>E�� oWݮz7�0�3��&�쵿b�U��ž�Ƕ��i1�!�;�Tڛ�����Q���;a��ީey�4��]9sK�mzs�&a\��2]D�И�3��p�����^�`g\?�:~S�0��=y�d��Od�W]+ ����q�4sq�y���߮:j2��A�z���wj����v��*���]QYk������YK�}��G �M�ɀ�dxW5��f{�DЉ�S����e��fLgg��ۂd��>.{��CX�D+��陭����-����G{]�i?v�vq��-����r��|��T5ԩz-��9��w@uB��t�ɉ�t�ّ�̳,�*�&���r{�NKb�:��c��:���9%\��T�:��:ֈY��y9��A��U�7�:�w����
9x6e^w��r�y!���{k���c�	��>��b�������Pr��z���H�:�%�0���1��|_��b��[<'�~��K��#-ݷ�K�k`��9W�[p
�����Q���f}=1u/���=Ϸ�V_Z~�c~<cZ�1����wl�M����6�z�Fx4��m�q���;Q��gu�����s��;�Z<����}#>���՘s�������
�(�C�-�*|Ջ����z�t*�ݐ׎W�:����7c`�"�����Ϯ$|�~�W��-����V��>�Bv	Q�4tR�g%�{�k����b2]��"��ݙ�э�ُM�]n�w�\t�=k4î0�^��/s�e�.o���3=}&��H��Q��5R+g���᮸32��(��57nrF��/�N_6�(Ҳ;pf���@���H�e�]ߪ���k����l0j��q��2&���y�ë�g�x�
�}��{�Y�
�<�/t��;ү��;�)���vV{�_U�!�ئ��E'�3^��$)��5+�N`2U(1�{ξz��|Ha�TkvǷ7���]j�4z���/�k>��5��A�$��ȮgqV5?�s��T��3�%�/{Ŗ�7�:U"��c�D:(��/�1/�Qzy���JY���%� XQ�#���;9饀���̛v���"�MT�Q�#����jf��t�������ݓFK�������w�F�C���|`a���`��S�r������3�tɜҽx�:Yͧ��n_nH���f$�ξ�P�}�k( ��Iq�����e+�Ty�o��:�uuD���wIo]�{O��k%֓[��$F������c�ZΦv�q�i���x�Ԛ��X���ð@u�"y�U��HWY���lm+���k��.�ZiK޾�/���o_u�����ց&s�6�{�#��պ��Cz�9FWV�┝;�D�Qt�n�1�w����4 ��t�U��[.�SZ{%fG�ۿ�p��F~�5QY��%j�JR��R�;x�#zV�X���iUq\��)�̼Ʈ�YFp3��V���j;�'8��#���mN՝��.�4�k��/C&	�C�&u�����d1�_�.�<�Wqv�F�p�:\�y��.�ު�n�r�*_V����)��K���*��ܙف�]{���uˉ"�WC��s*�fQ�eݗ57Uaڨ�]��ؙV.�j&����c�u]r vm�x��M��S�������:��#Z*��Now)�&��n<��>	Z��ӷ�y�Xi���yٳa⡎d�����qP��ѧ\*>Z-T����N�}v�HR����u�����D�KF�	�p�zJ��&���>���nIO��4v���"k&�����w�Ә!.7]Zc;K
F��Ul^��M���붒�ɨ��[�3/-� 	.�Ѩ��M;���$W[���;@��@k��l����5���:�ڊ�6b�ՕyBF������ֺ���t�R�g4�����MS�p�M��m�yo�?9�C�
���Ь�*�4K�Z�Ż(,R���ni�j�3��XR���=�X���[�@~s�'����oT�Wv�6��yA�Ǔ�(�,���1/¥��t����#���/i�i��S��M�+/�,�3'�0'��e�It�{�v:oU�뾬dڔ7E�J�h�}��a�8�$�ebx�k�Zԩ�W=��sm_������Ļh�[+w��sYd]_uf�+��+G�?\݄s`.Ў��|oKf��-D_R׆�9-��鎂驴/�Dc����y�r��]@�U�D��)�M�n��Cq��]"7�v0M�8��$.�w�Fvv���4OS��5jU�j3�3n�Jơ����、p̕f����X�t�,#���D*���ڰ�X���7+���~��{���H��L�I�x7?udjk�(�L��lxᒠ�+7jpQԔ����ʮ��mn�]���,�g]�e�"Z_%3��ok|�sle��(F�öݽ�Lֈ1��H�L�TG*stv6�R1�t�TR�����(��2�Ph<�m YuQ����m�@⮩ێgn�w���;oK���i�MK���|�j�}ʮ"�ۜ�����Ӯ�9�h�G;2t��f(���u�aG�F��~�+k��v]x�=���"�\"E�=ۡe	��^D��5�iƃ���kߧ�:���3���^z��g��u�@�os�
/���_Eω�5�����z��U��:FQ�N��Q��W��������(Q�%I�w��s]y��֚�a,B�N南�	�p��7�(�1i]�13?|�=��|�0����k8���M��]��?Ƒ��U־��Rf|n�rM���^��Lh�O8��ڱp��8 uފ�v���:�)��X�6#��:u��f�Q�P��d�[6��o�W-J�����)�R�{��s��U-]���ד^kd��o+�ظ�y��!l�zg���`s�au����f�y�О��o�@�pO-�C��m�οR���j_����MS�B:m���d��ex^�9��P��rv*�'�u�갸W���<�MP�U9��Z��2*D1�	:��xت��=�ܠp;5�J
5Br,zu���8@�=+Dy����[[���'Ҥe�%l�>������	��۰��E��}�-��!�YL*�u����\��o�:�~P���~Y���u�f�E�Q�똫�v�z��Z&���{k�,���)7�؍�͍��V��5�˚�<Naol�I}���n�%�Eh���&���]���q��
����,o��3_��}����;�����}D�57';��'!q�(��}��wZ ��+����c휩����"@~&o���3Z��\����k,�j��=/����d������T�;���3�)��.a������_�k�&���оb|���<�
��]0s���S�9�幛-K,h�g"nc���gd������x̝�5�= ��鎒β���A��?O	�?��
��2�)}/I��	^#pv�gFGX�V�7�g>c؝kب���d��8(��,<A��$���$ʪ��J}n��,ry��{������n�Tbo)-�\g��ZQ͸JL��y�Ƭ�w�B# ���#ѝD?UBm~"&1S��.$۪c� ہ8j�Gb�"]
�7���T��}(���������"�;ޮA�����+�ꇷh�dzv*�a����)/fgr%���,z{z棕�َ��W���]n�д��;Vy���(d�">~ۨ�>�Z��Ù��_�:l�m��S��dOlx�*ˮ(w�{0�m����
0X��Y�9ܑ��ͧrlZzM�[�Oe�������s/E�ӣ����#]�Ҍ8���J/�/��&M�Z1�%���J�ŭ��R���w]j�<H|x֔�3�tǕ��8�٦�(N՛�*eci�y���έMu8A9Tl^���z�q�{s���B�w��W�t9^��;��0f�{�J�\,��[��Aj�a�/�t���ȱ�ꪚSR�t�P.������h*i�?	��-z}I󽌍���̂�t����l��P��!ysyT�����?A�f�j����7�����B��o�쎿1H���{���޵x�JoK���P���YC;�R�20o
��gPX5����		?L��l���!�Q��W��	$
�[�V^w��E��3�Z��pu�1O����x��{��C.����՞뢸s�b�[����;+��|@�ɀd�]Ǯ��gg�/v*P�⸙�H�4�#ާVA\��]u�\P�R����y�O�
�VyV�ȅ9V���������TO	w�Q�Ɍ��ǩ�w{Ȉ1I�,���-�=�>ȭ��3K"�d�by�9\�X�)ط�X��3�G����X�������<�B��Jw���w��dS��_
��o�˕�f�D���Uv	�����?����4�&#cݴ�)�2_���O�L��T�1�9j�'ǔ����{����0j���5�c�Æˡ�"�bYv��3�t��>�S`נ���}
����)����l����m�ىduR�H]����+i���v
��PFq�v�7�q�n�uu#�mid5�8�]^����c� �+]�\
#l6+u�٪�>��Ie���*���$9ś�[�"��	u���G��i��9�2���x��CgXvs�N��ʲ�q�Q����ߢ��wY7�*����z ��Գ˽X�D�zJ�cd��g//�Wo�(��ks�i���=M�ݍ��g�'����iD��u����F(s��,XDo���~=<���m��bzc�#i�b���`.R)MnmX�u1����mH���R��A�0�}
�}��M��s�����gG����ْ�E�V+��z�����dɉT���3�3y�����KQ&X�&~��%������R| 5;Jv�n�QE�c>��vs9�_��o�*X�Q�\y�^7W�]
}��vM�Yo��~�E�����D*�nպO��>
3�p$\���㏍�}�F��}�(}@��w�h7z�������Zg�f�X�p��2l^���hB��FP��M9��X1�z1����4�kۛ��l;f��ʻz.�=��v��i��]Uof����@�R�$W��*Yڌ{+����r��{O�|uЎ���Լ7�~�y�Ǆ:�|���tn�]C��^;{�ҞpSzz��r��������!S|lW{Qղ���Y[	�����R&DE��(iw#p滙�#=�=�Fڧ��`��B�OR�_���)y�tf�\hٷ�;jQ��z�ɨԹv�҉ւ��3Y��#�Z�(��ú�'X�S��&8�ZC%v�o��:�# f;�d�y��G+fD��C]i�H�a̐�[ad���5���a]j�b�g��y�=r��ct0���Ymڇqfec�Tm:��ӥ�KG,ló��#��9�O8	�U����+�?m���;�u�]'7������ܽ��oF[9�Mh^���̦Yv��ܧ�����`Wv:�J~iu�}�;,�&��:fǈ�O$ߧ���~�on|���s��65ȹ>W���y7�E\<����6�3���a#5."������+{�"~��e����`�V��g���݂j(S�_����w�WP�ŝ�GK/���y||��0 �q.�x�Y吣g:�X��?����9�@�Jyޅ98=v�������޹ŢoW��FH�L:6�Iz���z��R��6��g��1���m�I�{;��f��s^�7�t��M)������I=�JY�;T�_1{�. �陷Α�=z�r�b�ޤ��z,����0����\�,��Z��ߖy�a�x�	yI�����Mu-�z������S9s�=�-f��>�;K�/�-���znL�#.a�X�kZ�mQ��<�ވ*�$}1y6&)d���z�{ܣw=��:����FWC�j���i<.?���PV\*�	�n�svs�Mr�܆E�����X;_�vs�D�֥�0�&�@e`�<ێ<Y݉f�ۮ�][��b�و��SW;^�;ϋ��t��k������JI��wTR��Tj��]�e��x�������px6�=5�����Q�"���я �~�O�x�x"��V��x���4+X�@R�#�s4��}�WX��`�������&�]6�����_{.�o��>C��sf�O�黉k�,���J�\����yz9��u���+�[��1$k�7>���u6������jⶳ��Q[��^K�t|#2�ž,΃��L*є���|{A��<M\h�N7�&틡O������L�@�+ӾMs[y�V�ug�z':��+�:@���^ˋ�#�ݟEh]���n����K��ef�YS�m*Ke��ُQ��6��j��|��Ħj�3�tv}�򬷲���ǪH�����oƄ8-~J�~s�CD�����<wZ��^�^/1��.����`���?�ʂ)�@g-�o5d�ӆ�65|^�[�����C�v�����ǖ�����ȹ����g�c!D��ɼ�UVa�j���+\��8GD���3�خ����V�M	 ��SB���ԵS�'Ex]���!����t�3���M��Q��f��;.Ń�W����c�.��<�"d�M/h���F���o�"Y����8VwX*�+z���5冪�7��W�ݲ��EdU����yw۴��Cym�%��!�B�PKZ�qћܷ:��\B=jGxM=�iO�2������dz�^�[ٝ�.���.�����P�Ҽ�T�!ۍev�����h�7Ofo�C��VV�+1����zN��jY��Q��/���RZd�P!^Ȭgsr���uf�
;n��>�p7f|@���d_a ���3~��c�^CH�����]�Fѫe�z��4`ҋ�	�.*�C�?V�.�	u���U�f*+Ty�ћp\�{��8��Y�u�������@���ȵ�.���ճÌ�T��F��W�?i�28;�8�^}�o�!I7h�=�΄٧<cӚ��+N⛊��.��M}>������\3�h癸�lݜ����"�

�����3������~.����N�C��>�lG�����d��cmYɿ{����qy��!�7>Ƶ
���7׵юb��=$jA�Wr�U����y!HUۆ�[�8uq))�������N�u}e��C}����d>w���6��y�� ge����n��Z�\+�s��)w�wu���#�6Ʉ��ft�}91��=ri�}�7N�6+� T�~a%�3���ǝ�'��<0eF3oq� )G���'8�F�?�,��G]i��?<�((pv�ök�?s �["�۬B�����.z�&]q/@۬cr.w�7@59�|z9Ji��η��8��N�nk޴�N׸��c������PTtS�GV��2�`K_���8v=��n	}Uyb`��3�]ɩ�uTv{ ET��Y&6�)�
w��͎�{)w*b7F����
nvV}�E�{��Zx���LlM�P��b�K�\D��9^�w���Ǣ}�RVRD!���J��|%���"w0�҃��=�遷���,�T�H�>�X�!����W��FgW���Ӽ�ҭe2�)���x�ҿ��;s���U����{<�5�u�[�V��$h�[B�Gu��d5�sL��Q>s�8Bf�zN�6ݫ���^�kd��T[�R���1u5!�J��[��"ά��(1n
�q��p�r6^��x�{��/Z�i"�Σβ=�X3Y#223��@��r��@����N}���0Ma�1PB��ɻ��p�ʽ��}�i�GL�z�������10�ФT�x�=�0�W�f������ᙫv�ځ��PV.s:c��/�\��g�<�b��a�@�<����21E�m��5Mv�8��РOk�(����k��R~���'w}�ik�e��]u�����SOn��>��������� �*>�u��P}�Q8���P�D�p�q, ��,���K�+�[�G쁋i���R�ӊٷ�
��*d�X�Xg��/t�̵�~�e^�.⢮;���m\gw�v�Mf�J�(sȬ�6odW��dӂ�h-.b\�v��Q�ռ���k��o8h�-4��9E��j4������Qqz(�䤥%}8��3�����Ot�=1���Y�8��p���j^��ؤLp�-��/^D��3\YQ__l�V:_M<bz�o�傻g��EۇKW�2!=��9�n%2�wD>����	���w��� LU0��)��y[>��2[�ՒY{���mT�V���}A�uG�H��yy>O������&i�+d�Wd�]���.M�:v�QдuO��;�k�ʺ��s�&*\D�;�Ș�LՔktm����k�}�_�a���0�%��97X{�T>�@���axp���b�S��ͯ��j��2t�/c�69��Q�c�]ǵ���P�t.�/]�փ<(FsV}��;�gnRU��@g)��P���|u�Pr��Jua�²Od�ڋ�2�3�t�F%~
�Y�O�=���$��jx�,�5mJ���U������Lo��.cs���=�)-���(�|��%�*�VT�y����͚�ʾ�3�gwU���;y]��_��K��Or�\m���ٗ�'����s���\��������o���3A�UHR��pz����z�����eB����ǽ��A�f�с`����� 4#��@��cҠI"���(e�zp��c������=�}!x.!�,9�����0�:����	َssߐRJ�Q�+={�/It%�sC:K�C��0_+wwed��] �y�omeo3��v��^O03^��,ھ�;�Ie��p������B���T�Bo��ee�C�ʳ��۩�����-�!�<�ժ�����un�H}�2b*�e�!H�}���J���a��}^Mn��Z��/#Ja �{"v���UZ����=7�_�Ƿ�mDg$�1M���}]�}V����t��ӣ��q@��3�vfᯖ8�o�d��!��;}��>�b����}�ޤ���!�%P�^�GA��+Y��xU�;��
�i�V� J�Q&����w[n�G�v��*�8�;�fi9��r(�!FƽQ���)��{���+0}*ߖe}V�5M�NZW�ʾ`����L�ɨ�U�����.�)WT��S*�<�Z��������c�&���y�Z?nW�Y��*����뵺G�x:�ϣ�1��ռ��:��t^�(��t#5�Ru~�4 �h�,�-���f��`��`���|.�����k9.�S�7�a?NfLˊ��z��Jn{���|��#�Vw�.`^���Ru���|'�
3n@銍{���9j���oS�[���{�g]ܯ��Гf��ԍ@(��?d����IQP���� ��=z��k�v��)Լzρ��ȷ�*�3��l��z��y���|#"�=�)]5O'�U`4�ّ:��h�8�P0�MA���H,�PP�+�I:y�U��h�^��E!�ER�)4v��䵶�։X���{Ў/rf����o�A�[�Z��a��ȅa����okQ�V)mǽׯ+ �J�ֱI�jU��5)���Oua�v;�*�\6���]<:b�6��f2��5��\���A,Z�ޥ�]��F'bc��v��s�Sx��.�����፻Ψ��hf�w�Οe>�WU��T�ᙋ\A�5Βkgc��x�1`�T�}�TEV���޹u+x���/7��88R��k/�م�
����jC
��;t��m�]]J#�v�&�\2���w�9�{I��f�W;�ҟ�Z�.�^�a,�+�l��9_GW,�m����ton�B��<�\�FM���~��]��o�3nZW�0h�ޓo�iGSʅ��SsN�s��k�;3�ߟ��V�C���V3X����2��:44��ҕ���]vȳ4���3"���(�f�UK��	���yV+�n��y�����>�$�����gYre�Z7�5r�I���"��q�t�.�8���X�/#!<m�>K9��V�;�5��\�Sw77�Q�:�B��Le�ɄJ��p�\���wv&���fء˪��B���#�k�D+,m�k����CWf��H�n�_R�?^���0G@���|�#�T{�4KȬh����5e��]� �|k"���W���r�n���&�|O(Z���I��Z����Op��ъ�o��։.�z�훼I�	���]M�@]���C��{�ui쫝h��r�m��YAwRZ�t�f�y#�x���w�!�A�YZ�
��)�e�v4]NV��T���h<�Z����t�����]�m's��Ή�n��O{7�8
1,8i�v*ڮ���j��h��/	s�}^̕yX��P/P���b
�M�-��&�����@��F^�!��h���ۇ�Kp��ۡn�<�i��䌤8������OE�4��+-�����<�����T�5:�w ����L��}�T�,d���АjL�8��Z4�4���lsh�&g�_Q�6�	@�9:�NĤtV�+U�U�Р�\��>`p��	�M͂<v��%�w>��}y��Vӥ�.�@99���g�ͫ������;m��79�c%�/�����3+,As�)���K�o=Bv۾YD�M:��V��+,S{՝�K��̣�����/�f�ce`�Mjcu�Me�<+E��]P�]�_�]����K����M���i�]]�mg]��Vǩ�⼥������stG+���Ɯ�M+���GC�Ht7�ɤ:L�ݤ�VS��K������6֠�[ �P�[U��$�� �š�˱sOc�'
�aF��;}�Q�N��ڲ��-Tr���ۼ{u�QH�y8�m՞�:��ý��\�9O�pgo�MoG׽ϖ
Nf�{ٶ���R(�z�x���u�E��e�5X��R;=��E��@C�ә�'owc4��Nv�!�|��G����ܛ���^p�T�[x��Hї�z,�Oʖ^Iͻ�n\��F���Y��{�z5j��k�LS������#�У!����c_7�/U�<:��H{��F������9JXu��0����tǌ�fM&GC��w��W7Q~��i���x�>�R4�;=
�!���=�G�����YYz�d٠PE��똼���=�b3�OhuXW�jޤ��z(OLEC�&$��y��p������}����k�yj5�K�a�U�TOF(ye)��ʨy�Ā�)�u���ã;�lmZ!������>T��>V|.,E!> ��pb:~����N��c���F�x�lՌYj/�dyw�	�����яu�5�`����.���~]{}�`ݣ��Kk�MZ�al��y��d��s
����u��z�	Χ�N�-A�������Bų]WO���z���q\%�� �,IF�_\�J��O��3i�q�fz��ݕۓ�֋4Л.
d���WYyf���r3o~GUҜڋx$�.v:�nD/e��}a>[d���%��h�v�q�F��/��Ak�� �W��n�K���m�a�D�P��ɝ���Z}���Z58V8ê�n���n��nwl?�u�7���*wI=^�q#tH���i��[nn��Mv��Uƿ_.��V˞����{�W�x��7�W]�N�M�wP)}��{95�":f��mb*���LWo���s��s&+{��I�����t��Z�T��_ �x�]#g+���N���ж~��)�y;��_C�x�o�3�m���>�,�G�򸀽�[o6s=��(���v���9��c��<z���&$����R��~�����g��t�Q��y	�s��O^:��:�]IC�6��)����C���ϕ���ߙ�a��O�{T�n�w�i�;s9qkL�B���������s�6�Dh3bp�`�Um7�}`#ו�����ȵ����-}Sxu��R�V������q��Q�Ή��~��)���w��|Vk��_�E�Ne��Ϝ�1s�'�/�r%�*ߥd?F��Yr�'浈��ɽ�蕎��>��7<�|�f}��穚�����.��.κ8�M�U	MV!�F��y�Xc*�rR�t3��l^W ���/l�֑i��lj6�6�Q#nI�;��&��x����ƛ|��w��9ʕ�U�ݧ�L��|���!k^1:�<�z:���m7ć8�INe��;{b�^Z7�O����辯m��xe�N��YK���W��Y�R�N�<�S-�VF܂�&�\���z-����;��אY'�U�$u�7�&��=�=y~y�5��F�p�����1o^z�r�h��
(���sE��\<�6�Lz��2DØɆJ�E*�����<�V@��%��Y�Ǧ[�4�F������y;�31c��_I�AW��kk!'����xgg�v�Y󚽧��$��*~�){�ȯ9����ck��ߚq��]�r�H�["�Z:?*�c☃�\���J�*�>K}^��j���𲛨�w�H�}�,�4hs�W>��c�Y2��8؉��$e��xG��h�6GR�s���uc@�6m\��хχ�lq!����>\*�-�[�6Në�JL`	��W��ۑ#�8Y,�^$�w�䆙�K�|`mBP5�'w>:8����v{5��.�E�`�`��V�y�Y>Y��U 3yH_g*�I9 �r�`l*���y�0D�Kؒ�YV�^�W�ꁉ�2�{����ɡµS�;��\�(Jk���ލ�:�+���P�j���P��v�YQ�P�	,'�K\2�L�\��u��^8�J{�f�J6;�ےq��.Ҵae����ѧJb��u"�>�,��)�rdI&vp�W�#z���x��>P�zG
7ި�x���X��⼹�A~��0}|wP,��������;[����c�;�LLPMB�$��g^�Sȯc2�<��R�����L���1s��p������L^�h*k����"��~j�jN3��ݘnh��^�MR��{��x��O7�?z|����ϯU��� ��}]r+���I+�k�1�w��.����ғ�c*�=�n��5p]���W�W�E��`P��_�:~{W@����F����2��qz(�_�9��5�v&!��fo���U�i��O��u�J
���??z�ljZ��J�ULl����f�tN�ɝy�̊+�>ӣ�;ܮ�nl�2�'��>�{ؐ�);ZiAdYO��93��fb�tlG��+A� 1�Z��b_l�H��A������ZV gT�=F�y�����ӭ�%����w!����3���{�3�&cG��V`�6��˗<�_��2�:5���̞&��b��Q�GM���+���<~������Ā�]=@�1�i0�Ӑ�j�Yfvc��8�]CMחE0��]nv�2�*d�٢�=�c���@^����aj�[�( 8��c��1uqMr��:�nGӯ�[Ys��%�,n�Y7ڥ�*��Za�^�v�Y�2�����-�ϒ���l;��z�j��뒭Rp=�q�
w��O��9^�5]|�w���v>��v�#lH3�v���N��-�Gw�i-�"}Nޯw�H�g�؂�>��/w!�r՟<CQ��i���(F��鈙�����Ҍ���Ll�\�k�*�xcq����D�9#��Gp��U���ӳ{�lfKfn���ck�O��*���C�i^�IQx��fr^a��:������x���r|z�T�{<y+xw\���_�X�:�3�Y"�z�L�8�S�5Q��>T�7���;�O��o}�[��C�8�Z��ys�z�A5Y�DG��q��
��C+qA�����O����*wH�|#�&�mL����,�}�V|5/?+�;!��۶��Wj&
^7	��
lV���Qu�`"Oe%��>��^�U��M�eCbxS�|������o�*�~�{&��c�tTo+��J�?T�>�T�1�ţ�P�\�����_bkQ⾊�[���}��;��zk�|��M��_,ڎ!��AT#h�������F�0"���;0�����l���n8/"'��B'���R��#
uڍBM\�l�qo$Kֈ����tn���J���!K8���7�^�կ[����aRܾ���0�7�e��i5Y�4NQ췥�؎��m��{����6H9�z2�s=zAՋW�΃QAX<��1�ט)
{��g}f3~��v��`�-M�"�_�t��	O@U�Y�Ħ�]W�*����L7�qkG���m�t���}���a���%���*_eh�%�t��%�P�I2�N�ǌ���i]X����W\�K�Lzw�G�׼���n��}el�Z_t~���<��93�2ͦ��v�ϋ��uݟ_�y�|�ܓ��8ٹ���@��0Fz��aA!��Q��o*������g��(W�
����$IQ�BR�?�.;V���F?3����[�8l?���ǵ��ۂu5�p�u�s0s�:�ut�&�a_5�Ɏ��9��0S,C�	����A�:������z��5ܪV�ƨ�P�a�ړ��`>��L�������)Q�Rw�t4nf���7}�5������J�D��K{�;�Ƃ�GqG��hm��­�����߲�'�9Mpw�И��,�ޫ/�L�Y+2�'��v����5�-R�y(�!�E�`a�)muj�4�����T�Ƴ&]:�s�^Z�����vr���tkmPhL�݄)v��n��q5)�=M1\���{�n�{�Ӡ�L��{F�+�F8����p�g1_,o����B��O1h"7�5f>ὼ��u»�Q��5�q�j���D�轕1WY���jY9���{>��	1�E,�3��i����5�b�����7h�~遥*�̋>u�zb��MM��vv��1:=+��p��cԏ��;�p��/q6�6=!��c~mR"�cv����{��^�bB�=GJ!�ѾGF\����Nu+�Q���ܿ}kG�^%���Jr��dM�8�zn����5�G�v��ލf��y9��;3��W���n���ј�y�u,�Qm�ee��0�?p%��݇T2�P^�X���e�Y4a�3��dO�����k�C�c�So���F;!٪�XhYfM���u�<�@�t�3�]�ך�>��1/t��v	���}�>=�͍~��F˅�~��v%��I�jғ��{����88���L�ە[��¯�!̈,�"��x��8w+�͉�G��E��m��u�.@��O8��ǠW+{����������3 �J ���5{sT����W��2G_Ȓ'��Nm'��s��ۼ%���.�gM����vW~���8�!&�eI�d���ҍ�M��ѴuPPw����*Hyr�뺕ݜ��q�j�N���]�%~���:����ܷZgYOF��)l�)��`��u[-+���(�tںos?v2�e�Im�����ƾ�2�<)���X��:��]߼v�6�Ur��fݬw|�n~�j�/��U��e�ٸN7]����	D���nX�^^���Hf�����k�w:����S��ը��װ*�_f��g�/^
�5��\~�<7����K�-�����%���wmy�$��G����-�����|O�8�D�ʠ�$`�{G�w!#�F�Z����t8����N�œ�ж�[������W��Cȥ�����V����13�����m�>�{����r+�x��es�֏���K�Y�VK��4����?��U<��i�=iIx���Ã�l�&�T��2���`4�4�}�z��>�����f9�Y�Q�&�ؿ���ʜ{c��\��7M}ۃr���Yf�;7wW�Uݛz2*�|�J�K���;P�r�>���׾�ü��*j�s�����Р�Ԗ2m���B��L�3v �~�d]a�{o}Ȱk�.�U#@��O��^���!ࡻ�j	;UC�[<���F��P������*#,�j�<3��n:GEO�Fǅ���m߰���f���)՛��f�������N��;fjlS�n����&��Bڎ�p�V{:hB�(;�\����em���L�R��U��1G�O���m�Ӊ�}�ۺ���5P�M�=)TZĝ}�$��be�����bk��s�f�1<���H�C�{��K���%���i>U���ɵ{��sI�����|��y�<7<�]H�r����|i�P:����R$���P�߬jo�:kŗO�s�\B�@|�b�&�u	F�Cpb|�x
�w��S'޴�7v͡��!����φ��-^e��r�u?n�6:�d��c�q��/f��V��u��~�� >kB�����߬So*fdW7n�s�w=�3P[ʷ%���Tm�%Q�p��Ǻ���>���mZ{�i.�0�)��ie�O�ǘ�U�WR�^û��3ё���jg�LUp��6�ł��3�c7gL�l�����sq^U��>��^L�p��9�7d�G9�"��p%�^��{�(p�絛;F��I�L�����/�m�8
 3���'ڼ�~̳���4�z�t�%֟|��08�ԧ��F�k���p��eǷ�LոK-I;��QـLum{�Y�jł�Ũ%���{F>�u�Փ�kI�u=�\�yE4��l���M]ʯ�:��Xx�lt�vK�A��M'�X�|�}��oe�ȫ����+����P��N�RoeL�����vh��ɩ˴A��'�ٙ�:�x�N�J�h��j��[�-VL�Mgf�������׭�cҲ]����=�ˍ�+}:���ӛ��	uڶ�]���V��x6n
1�����Sw�n��Q�feujՂ�9=�[egt���W��G=�ܶ�wC������՘������PNK�V�����T_�dǯ�\)��ڼ��Y|򔵚�mV#�(�"w�m���#U���w����\�SL�_NuÏR?0��U;5��_��A���z����k+7��0%�x���,N��\�YCJ�ުt���5S��/jMG�Y��ri�����c��$�0VR~uKEi~ݫ��9����Q]����,���:��
vj�u�x���<3)����6�R�湨w#��xl���б�����vB�SO����Dh� �oS.`)����"��{(X�$Io.�6��.�+pP���|T��+�j�����*�ծ�)f?�+�!�����Wѥ�,h��H�U�(,3�1R�p������&~Nr����8���"c�E\��VȠ�o/FF�Mj��������7�J��'�1��7ޣZk<�j��^:b�/�W�i]vs�zJx�M(۽��,�e*hg�.��=!�)�� T����=}���T&��H��8���+�[���w��c�&���6�/4^�
��j��H I	
j������V�K�8̪�c+rW�����ǁ��-�k�� ĭ9۲��#*Cy��i���W&Y1Ti�P��}�Yӎ����{�V���I6��u�Y窮���������]tAbP2��8T���	������Hr�ް��7�!
�;ة��G��J|/^�s��^��ܜP�Ɛvi�j���MK�Ui^n	ul�	�ê����t��3K╕H�����s�m)�j�Q�fu:k%L���p��P��;5��GOb\���h�ub�]�L݉�K&�K)�$։��9c)�Q%p}�j�5����
�_*_���-NKQ�8N�af�i{)���S�p�h����G9�gV�Նk����z���5�wqC�sBNRs�ͣ�+iͥ�^�a=(]m�a^�T�X;\��,6���	��܂�S�{�����*Z�S9�s��gLgU��op9Qސ�ao%�b�/�g���t���t #���-�<��rb�9Q޸e�)X���U�q�=WV�&fYYn%�IDcг�ֺV����[2�C��8t+��z�ru�S+�jv��GS`�;^
ɐQ3s�<*�����Oe;f-���l�2e�ue�F�u�I�U��q�a�b�YZ�u����E�J�I�^�6�X9j�<���ۑT(��-�O]�00�)��1]	m�ݹ;�x��������4o:��㚕��Zt:o�F��q'�x��N�n��R5��F�1�W���4�u$�|n�z�j���E��_�uO?j]��zM}$�t��m�$01���R;�I�O>_=g_t��{���A]�7$��N�)+;�0� �g.L�=��5.n\ݣ�B����JC�۾3	�e.Zյ\��S��i�/�o�o��al�i�t�17���9]�]��s�U�4���MKp�y\g�p��M��NE���Z)Y֧�槸]�@S�:ܴ!�MF��Tv�.��.���\ u� �T�w{Vxd+{��(..����4��Q��{j����!YnWY�+�Kz�|
�DÊ5���r����]H�`;@N�qÿ���%+l�1=9x^5/��騎�ّs��.�������7K=��c�	wg=����q�H��j���q�m 7�sc�,��N֑��޾�ĩA{�*�.�^�fR�E;ߵ��s�F��S�� �)c��q��3}�-���;��%ʙ��D�r����lEvuw<{nM���w���h���48�{Ċ�[��,���[���[���M�l����w�{Ws=���nHҨuj�k01�����a]{�S�5u��W%v ]F�>Aw+�(88X��d�E,�-s�m�+$=ܯ3����3�3�������b.��F�lZ�nL���DS UܳjAή�nMsf�rf�w��$��uyep����93&R?���-fe��p��5�rK�7m��(*��������I[�KQ�u�YN�u.n��ٹ]��{���Ŧ�]\���S���x��ʻ��G��V���*�Rܬ���[�v���m[�b�	8{q��tX�X:?�%EDa
|�<ݘ����7��/O�M<��B�ƍ�?�3�z�[OE�qK����g�<������]nO���0����u��{�l�:��jF�x7\s1��%\$���g���s�	�R7�y�%�-�����dz������I�s�RY��P C�OLwR�[87ww�$|��X&���yī
/۬����x&����HW^{�����9¡
<��O����~a���
^(k���(��s�ǰ�L'�r#E�CN;�*:�@�Hz��sW袽s���DY�x]��шГ�DU㺯��j�  �(�H�ڶ����s�Q��U��}�4L���#|��V�����֊��lX��-Ï޿� $�q���H�ߐ��ViTv�}RH��s������m�eZ62v�O�΃����0�G�-���5K��B�.�9c�RU�W���İ<rV���~ɉ�����zS��M��%U��=t3^���{[��k/DBDWMߟ�t���X�wUb�!Q-8���g��{�(�19�����i�v�k�R���� ����?�|EW)�l�`����w&λ8yXٕ��u���J�ho씟nrũ={�9�]pDp8�A��Őq-�M�,ʰ:����S���O���A���{Bx��- ͬd���8;��j�2�wj�Qc;�uJ�|�q)�c�0qNж
��k�S�z�P�ﵐ�u�B�S����g�;Bzf�+�c!�j�S���B�F�8����e��~��}��Ktf-�K�ve��-T�J#��� y�Z����˭#7]8+�_�sܘ�F�y�u'�w��GRѧN�*��ǧCтCp�4g 973�ez.��L�!	e�?��Զ�1�(���;�7Q������ץT
�{!����N�ɣǦ`��[ї��KN��� |t�`�P�h��]R+���J��˄�Ʈ�.l�Mֻ`��X�ou�:V׻ �,�:����$�iޥ�Uqy��5���nѡf��b�o���͠���~jf�k3����~�;��Ш�n�\�,��C߽��s5fe�C����@�>�����}�qj�)���)M��2�z8oTC'����7�U;?;���6�?-���n�DD���1$�'a�J�M��5��:�^Lfr �{f�E�&:�M��N�R������>��X��k]z�����%Dd�O�A6[��xq9�N���������Ul�e�ر�,}cq���!�:�"hD�A�}�3>���^�$k�;v��N�I4��~�Nd>��'�`o��	��a;�\�
���٬I��WN����0,>��1VxE�����2~mBS}�j>ݺcf�>'&�Pb��t]�q����cn�ʱQG�a᧞v+�(��ꗉYga���̡V����
�˒���Z8��҅@���+��ȥuz�2�C�9;Ԕ���|�J`EH���2گ�M���U};>��V��_/�\gF�:�ON�l�yA�T�+�SG<�E{��A�p���o�w^�p�m���&��d��*�����1�"�3ջ���]�J�V K�T����,*/��C�"�lNt=i-2jVW������f����B�^�f��|�4���X'����GҾ]{��*+A�b%$�܃ۆ��]I�[���P$�Q�o[ϝΪ��\�V*B���P���Xm�?>>�������7b�륳��p����L��vT"�x��+��M|&?彁{��Y���,]�Kt\�����՘����_� ����귧�j��F�Kl�>K���'�&�{�d{�'2��¡�?	K��g~Y��uDr�q��z>��3�x���D.��-�x�썃7�_{��Z�;�����s��������ܫ끦xOL3����������4C�>��77� �9VY�+'���L�9&vv�pI�����?���ǥ
�^�qE���|���=���X���ͳ���kaW�^՚I�xy �9�5��[�1>C��Wf�D���Զ^ؗ?o��c���;Dr��.�9D�ůq�PW��erMI�G�k�4�1l�ή�ƣ��ABُ9�����AiQ�("dGq�v�
\\w�6�<����������'�]�r����gG�B+ꩃ�,�#�MץnE�&�nɋ���zw��|�$P~́���dk~����9|6Ue�I�@c�]?nl����g|�1�!�3��L<�(���U!%�*��n�~?�~7�6W��0W}�������թ�s������I�}�r��h�]"��/h{��GO$<�06�ˆ �i���ܬ�� ��>2�"�za�~y�� C�*jc|�bT�*�����.���~�0�0S&㋳�y�9��-��|G,�O�LȆ�9xE���F�h�Fey7F2g��})��z�p56��>ή��%�ն����C�	���b��#��e;ƹ���l�n3�zR�_�v�[���래�vd[l*#=�k.�S�P1���k��Uf��aR<|!��gq��z
�
��R=h	L����q��Nڜ��o�z���E%��4�P�-��0@��;�A�S���?$�ݻ���ֲz�z���Y��>_�0�4.�����FEݮ�1���xLi�"R8L��}�lV��|�
�1���P��dO���Ԇw��e���J[$y?����������}�8��껚1�^LT36��c�^d�5n��ȩ��6(�($�T��b���6�o�O�J��vf�DV�:ɀV�MV�J��e.�Ǻ��uX�-���Ή_������{"|;S<Z;@-�ݬk���6WD�9ٻ�._q�����>�� ��iW$��gu�Q]`d��!��zB���9	HR��5*g�7�ȹ�.�L?V�Z)XN-ᷔ�$t�����m�ge�f`��z�TCu�Ig4�L�'��Ve����7��u��|* ���w��D��YÓ[���gE�u��q�!�ٽ�u'eʳ�U����3I����C�s�̑�0Ӂ3��O��ϒ��LayaRE�y���zU�&J�68u�y��=6H�L�]|)֟�¯�0��><�M轿��� �j�	�k�mN%�����2��}��A3P^n�A��f��c��@rҝU���z2�r�ӥ���9��.$�&M��+�I�+g�ި��'hB��G��M��v�/�ўܖ����3C�R������|�	��Gde&r�M���z[�*@[�W;qc&j$ 2��qǷ��R��5�툤��ax�u_�*����:3=&�U�&��hq�E��P��a��A��;�i6.�dyy����}g�](C�B��{}�*�����_���_l5-~V�f�J��H%�è	��[!l������s��T'�W
��Y+�8h�u�.j	��#\)n�T��M�h8%�\8I΀$����Hd`Gz^@�z %z�[��{����͒Sy� N���Buvr,����*"N�"{8)��?r
�iM����#��"����0�{[V�A웗�
\����3A�ﶻ�$l��R�}��"3�+KVDәY����,Q�y�VM�OFC	�v��vE�$[���r�����v~���
>㾭��/v�Y���Jua|a[�'�*��C�S�硳g�ݴ�^o�-�22�V����W���yK��T��n_aa��,$
\X�l2TC���s�r��Ϭ�<�ԅeʿ�b���K1��`}I:�ѕ1��q|��$�!0	6!�SYT�Tu�/�2���� ���fI� �${ɨ����)TC� tTg)��V���"o�!I��,EdvSm$Q��[��(�P�w��z�,��]��������h�CϷ@{C���&�zQFL<�3 D�����>q�0R"��Ȼ!��ȡgu�Č��\�M�g@$�͏z��lĲ�ȥ#O����uY˩��-k{�isM�V����Q��a�e�(BH��f:ԝ-1@���h� Eː��x�B��j-(ǹyA��@"�� ���Nlb��3)���j<(�J
u�ج X,0VQ�=�v�1@xit��0^凔^Mw�DH�/Z����dUj|�G���Y���Aϥ���l5���*�h�D�Yɜ� H+R%��C	8r��$J�p�M`H:�}�P�粲�8�"�"[�MyĖx�U�k��j�[�%����l/:�[�`�*�!���L]Q�mI!bQ�>~3�w�t��Iq�̸� '�4`��XY��g�,	�d"+��#��b�`@���A�GK	��e�&I�8hM�o��PU���y�����Y�^�+ď�B;��Vŧk?%���?� �뻉�vD�1�G�x�]�k���41�2K;�)x�����k�����뤕�o���e��-�����sVP�,�2䮽䖶�����\i$l��3�on]���76��d5­n-�"'_�,��Q�@��i�dy�&E��\�6n@�Qk�Iu�v	kӠ�pR�'��2�k�6E4F�#���5�= J� �"8��w_#!.�u�88r�z��[�*^�5.��kn8�-���32��̝bob�<���4�������W@��� f�,8��"m�]݀�"�=M�(���%�r(Mu@EȂ�xa���b�'�	����f�qGQdY�	h0a�Gz����!G(�8r���,�'�N�?Ci;�2B���������۾EwEݔ/'d�q���f焻�[����,��br�DC���S��#I�@E�Hp��"ψ�|�d��$�;h��y12�.��/�E�d+lyY�8���+M�z����h�E�@@x�#�� �"��0҆��{��⯩�= x% ��H
�z9�Y���{[
���E�`T��4t�V}��Vx�r�`r��#�:�z�C[��ix�����<��x���vÖ��(�fy	�+\�Ҏ���D�;X��$d�<XxԢ�n �g$Q1'
"�r�	v$W>�6�"4��a��Ť�5�� ������z���g�i� @H�q^<ϡ���ͰJ-�Ľ��8l"����G�A�3�����&�&0����'~���X5�wg}[%��ʏ�>Fw{�m "qu
����5�E��ˏP�6T'�.D3��A1�B�f�F	+�1��>�1%��ʶ%��U��f�@+Lf�P�� Y۰��|I��Ԉb�JC%c��������wEc1��M���֊�܁���jvg��[��`v}�y��,b���+�ܾ���p�лb�?H$�h���Lk+�`KȔ��+�H��N�^䙂[�<�8R+��[�::[�OR����Z(���y��@R O�,��.s��i	3�x�?��w���+n���|#��N�Ypl�Q7�����ր��:�6���zk!���� �V�[&�Ki2����t8�+`���K"�έU����T���g�®���k,�׷s�hW�,�4�{��k�S5���q:P��B C,@��2hi�NT�xL����%�ζL��: �=�j-��d�,��<�p��$��I�@�ϣ���Lٶ�c� E%Û�.Xz�G�A�@��&����u�ٙ7*q��Y+����7"bǈJ]ݖ�ŖES$jf~JX.�`K9��8��ԧ��f�V>r|2$!R��#�+��R�����9����0�2��A�8��p��ÄY	hPXvyS#����Y\]�� �dp�\�A�o��m8Z�:vWɂ�[��$<���65F]s�0&��L�� ���["���$+������o�J� ���,�� O���.CUy�15���4k/��e��F�n�@��✒�*ᅐ(��@1���4��OǮ�@���G[����Ĭ &�͈(��*��DKAu�G<��:aM���awL@�f�=N�D(a��a�JX�.�W�N ����t|��@�vr����8g"�EX-N&�kUi�� OR��&����rK{v���@!2�L3� =�U �������N��Z�38���G$��2��v䰉L3����ͬ��^ �9r��-o��vR�c6��<��;|��<�/>T���T**�X� ����VR��X3���l*m�[�#�����ɸ��$��w�^�����Ʃ��]�8�����2%�aF)N޾��{�]�h8�Z�{�.I��.7V�w�}�Y����7�K`#ū��B��18/`4p,|CbN:�SE�� ��C��=*@��to�0�3^L�i��Z�6�狱��2^��b,���g*)΄\�<X)K*��Qf�m�%��-�z��D2BqZZEk�A�i��"H!��"Kq�oWet�P��N�@���Ÿ��}9�k��(�@m���X���4�C�`��ˢF������{�4�,堚aŸ�ϋ�̲��l�i
6\KȒ<G.��=qY��A��uv,��A�5�ȷ�n4���8[J.��j�v-�\���D�$M�DA���l0�<��rMH�-���^����2��E��YWW�( �@'�r�� ���g��K"b� �@6r�$v�$"�Z=h3�==$6S5�>L��Ah-�������Nb�����r�KrB��`F!�a��.B6a�EC���h,ʪ��5u�!��oi�e !E�d��$" }vO�P���c��1�{e�~,��Mk��adBL4�,(�%�#Ň�S2���dF��ɪ��ް-�� �R(P6E�(e]��<[�A!����D�L������7|~�T_���1s]��H4��[�Af����XH�aD����eŇ����\�� ����a��@���8��T F���a�� X6r�a��VX�T��F��I����ᨷ�I5��@�\0�!9b��ɼX;5S�.�@/�Ē�ũ8F����Ap5ڈ9�����]����7r�3&��E����ds͘�츱C��^�q� v��vj2��E���ޔ��ܧ �[�4�4Q(���>L*j@�(�7���X�����o@��b1f�hf�a3��C�V�xfU/Z���bן��{�"̿V��ɋ��YH�+I��(��V^Stk&���A��2�b����xr��3��JɓY&'U���)2�b�	}�=r�>�)k�[ƻ�5e��J��T�]R�vJ[}�{ P�K3���'\�;�d]D����Y��"0��ےͤ�#�Z*gL�O�ja|���0�.����`h�7Z�<O��4�Š�PZ���g�8q�����o�X6J[�`,�XAr���ܖb|CKZK0Lu�ه)[��	�@ Qf��P	�P[�7�x0�L:l8X03���O���^���)�˕�s/��6� �m�,��a�DZ6�,�R �J�ae���`�/� 
�d� �	�S-��CHWt3N�gat�}I��K2�W�瞼��J�g%�"��u�a�h�� A�5Dǔ�q%�K6�n>�-������'��C,�U��L����Z�0H Y �����ŀ��ۃ�������{{�P���Ka�'� ȴ$Q ��d8��MC�K �XP"���0���$�:���`Ņ�"[O��Q�o�,�1I��,�)��b'6�0�&��d7�	��F{��7&�S�_:����g.�@���^w]�H,�2�v �m:@�\��&�BHZ��=S�P�ȁ�7C$ =B�	 IfdF$��6ZQ`�Y<X 6y ��k��.6�,�����5�Y����� Rm�G��Jt�qf�@ثP X
�Ť��C,�a��5�8���r 4��x�� 1,	`�XF��l,��!�<R��t]�K�+缔Tϯ�9�aŤ�4�f)ó3�k,�$0X�" E�qa�θYf a`��mI��c� rj 5�k,aܙ��,����mVR턓���Y�XR���ae���X�ü�5 %�� �� S0�M��0r�X39.�a��fY�l C9!���}p�Ř!��o3\�rD��#�z$�M�3x�E�"�Y���� �8�0D0�fr!��w$ .�5N­#*Vc�s�U<���I��� �����f����� f` ��0`�1�� ��� � �� ؀�f] ��3'��0  �!� ������0ffo�� �3ff�݃ ���߾������`�33g�	������wC��`���333fo���3337��=� �3ff����0ffo����w�0`ߒ30f�\+�0`�33h0ffo�� ����A�f�����O���y!� ����@`�33y�����0����f0ffn�l���h_�v0ffg�>P��8�337�$X0��������PVI��B1T�&��� ��Ͻ��/����f�   �G��Q��Ғ�m��X�ԅA{��D^�щH���q�+lE�jUM����Q-1���V�h��v�D�ے�nb��4�O�����9k�L�V�'fUIt�ƕ�Z���ֺ�*�h��뻫`�l��JUU6ԥӹ]�U������T����ѺТ������(����&�����'YUJkJ֥IS�N�٭���Q�����Z��"�.v��❫Q%r��5��P)v�B�Ҵ�:�5F�h�on��
���)JS��@>@  �ހy  >� r@��_ke�gv�sU�F��֕���9-m6��w�;��U=��<=o{^����{�z�)��ь�;��l��Ur{j��2��ʄ�Ro��0���Wp`[�i	�zڭ�[J�mNG8�޹�٢�֯s\oc��=�cNt *��N��Gf
�����
���oaנ���Uyw�QvӼ�������U��l*(��@{��[oG��ڧ���=�����mݵM��{t�
�OF�k�cA�=�SN�mG��k`��z���]���SL�F�y���ͦ���U2V`z=��]�J��R��:h�%����d����m��v7�v��`���T�U�ۺ¨i�=�U�5�73��r�=��1��0��&�*�9�\:Pv\zs��p�*�	)�ۺڽ�u��Nuz4:c#� ��{��޺���p��G�v��Wl��W��[�펯���f� m��Wa�����hԽ�:��Kf�V�S���v� �f�k�;��[��R=��e7w
���tث7w(��z�yWe����a��۠{ܝ6��8�EgvP*���l'��T���%X4i���*���(�(
�yA� ��Y{�����ǡ�)�v���v�mV,kY�v�\�	�J�s�R��pX ��B�h�ݮ�]C��l����ڬ1-W[F�J6n�3��z׶4^��x�r[j��� ��+��7gZ��:�����h=S�a��J���n�z�ݳ�����{�SeVON�[hn�A<U�w;��k�V����vB�5���4	4�\�7�WlX��h=SռD^�����'����׮��z͵����:�z���8���MKVuw[[���n�]m[kf�u�K�n{oc=6�]�{j�7�  *{L���* 4  �  EO�0�T�	��с0 Ii�4�1Oj�AOPڍ=LGꞧ���EO�A%J�a	��&�L�~����   C@ �T�4h     :��{���~�_��ez4�-s��g{k�X֒��.:I�4��M��`��oK�c�e~@(������*�q0��(*�DZ��z~�S� ������EUt�E*���;�����#PE9A �E�/��@D� H����!P@/P�*^
!P�QE�j
��!x%��TT�%���-K��@A-�E�*� -��T��+h��V�U*(TR� �D� �((Zh-@J� ��%⍠
� �E[D��D�R��)h%D�@P�E�A@m
��*-EF� D�"�����PV�5�!P���Z	P*-A��T*A�T J�ȍ���h�"���#QR����QA@VA*"�T�Z"!x#x������(���PEV��A� 
�h Tm��h K@���-���Ͱ�C�r�<�;�,gyr 3,Su�kR���֖v�-Z+��2��-V� �-k�c�1���wE� ���m���1�t�kB����L�r��eb��o`D��'gw3��w�\��uqNI��`��Q���x=��tO@Y�س)�{����g��A��Y��������=���u��,~� 48�����9ga��] �4��݊<Lff�ݎ�)^��2��䤈���ٶ 1Rb�Yk� �g_��̹��-����)%- �9l�5�"�.%O��]$�*!�:����:P5�Y�(p��-�)�cXA 0��ʔ;�F�ZN�����=5Ķ�)�jЗF����k�e6�BE�t��h�].n�~�z-XF�#KP�VL�YwLS�V`�T��q��[�Y�`и�R�@6g*�Jyg)̤�0
�-7����	2kfB��z@���e�Y[��M��021Oݸ:�y���h�#�(�%?�DIt�Z�i�[��g%>�}�նMΏ�������ԲpGhape���*x��Y�lQ��#�I������W�i�۲�ʝs0���V*ʔ)c����*]�� �f��E�+DMxIȝ]E;Cv���Z���Hrgx��Ab���������"�G5���6-�6��g2X����BӃ*�Y�/-6�n�.Z�D��!��<���e���m�0=��)WuiѮQ6ء;Dg+w��l�YL�o��5����3:3NZ�
��n+�,eYH��+7�p�]�]��ѹKB��	cXz5&�P#��Է���Vh��$�pj��5��1h��i�ЕK�LB�x���@��5)�([�e��V�D����4/��c��I�$KJt3������ẌYX���ܽ���(u��6Ȑ��ʁ$X�oRÒ�L$�<��W���]2m��<j�u���	M�Ϟ�(W���.�o+�+�R�4={���x�u�|�ޥ��%�If���&�B�8�T�a�]{�-���L\Dqݴ�Nѩ�R� �qH$��L-e &j_J��W4nc=h��e	���0�H���0s[�D7�"4��"��j�Y��S���V�Vs�P���KDo"�����ƫL4ӝi9Wv�j䵗�J�ft��w.��Pi��r���J��7� X�-
�<��c�$!:�hvp�پ��oj�2��kҢ%�Z��>W9�o#��}�-Ί�-WC�B�����2���]�{XTрYyz��.=ݑ;� E�����
������Y��c
������_  ��ܭx68i�8�]O�{���~�C�._���ۑj�!ۼ#n	���t��.t��9ٽlҫSY�r�[�:���)ٷk�S����Q�-�b�Ẹ�[F���A�y�Kߗ�y�W�76�a��eB�����B���;�B�e�*�Zّ$M��SZ�qȢ�
�ŋTl�R��f �8���Z����F��HL���+�!�V��U��S�,�ǔ��h��	�!�-����� i�/��3)����ׄ����{bmL��U x���%!b=��}�ϟ<Q<7�V�I��FV$��)][�`e�_�+C,ˬ���ǹ��V��X8��Bֱ�t��Y�Eru�o0f, ��6���s�h�s	a$p��w����R��f��Gr��c��q m��P�|����Rn��J�
�Ys�m,4��m�S�Ѯ�Er��&�#�&��
���%�v�l,NdJ�o����j��@�>�ڔ���N�����W��F�̰5ɘdڷ��j^��:n���I&V�.z�9U�c�e�L��ɴ%d��֐Km~-<DZE�nXІT�TL,6��ĵ��E��^�Y��g]��6LTvӺl�C.�G�8�h �C(��E�:ܒܶZ��Yhn!&0�f�5L� 4�y�dd�:�=�P8ɤ��V�i��t�!���3�;�Q%;8-�r�Q�n�Jb�.�/�/���y3bQxZ��1�,���¹;GZn
#^u�nPG��:�w��f��Ӳz�";�̡L<r�/P6��Z��.���M�񞔽`t�w<[�f
[,`�O:Y��m[�Az��"���5�F������@"�d��C�[h��wr��j����m���ͷ&;B�����s �Ĺ�b��ƺks*��g]�紅��Z�M�<$'�
������T{m[��q`�Tþs��B��z��7WFbw��1�UPH�F��Ǉt+*�m�.��%E���V�J�"d���*]i�K��i9v�쟱Q�r�Ɖ�14n�c�NSoA
�T�:���$��f��F�J�b8U��e����Z�J�b�~��y�	��JèSmna�7��~}����#2���(�n`/�,�K�����L�֍*,4��ν��G�.��K���66(`ݗt�vXWYp=��Q��܏j�'�$(����1s���p��=W����oEފo���hP9d�"��mb�{j�c�0�6��S�dIQ{�U�� �^�K�N�M�N�b��Y�T�.^�Ed"�фk+M���WܷX����GU�j�+r�hr��n��Wu��J̛E�J�j9W�z`�u=;![p٩�����!�nYy���̬��U֞M;J��K����1���J:���=�c�sM8�	�$]x��/Q�\�.���[�eNʀD���>�0�]f�J#E�ջQk	��$��X�+PǮn,-�mڠ�v*jVV�\X��.�]�B��;
�N.m�(sBe�uX���^l��٘l�R��b[�$���X E���i֦�v�͚�u\4&m�����n�圧p�rb�{vb9}C޳|��l���ʌ�,A
�xf�,�ظ�bX˫8�?��T���N�i�1uN�YhY
k%�F\��E�,� J�B�FN#�5"�s��n�^�.�g����Oe9M�f���jF۾[��<���kR��J��Ι�t6e
״�Η-:PV�n ,�D\T��qs�,��DW������(���f��C*�#l�:�o�j-��p�(��2��I"��5r�6���tޙa�u�P�Dҫ9]k�.;���/�v����]�G)�o��4�f�[�O�D�Z�E�g1 yR�B��94���H��eܮ�d�XpY�wu����$��o:������]nm��5ƫxa��(��՚�K�wðp���!�j�|%Ue����G38NI�����ɍ�h�wM��]�w7�i��l�P���ަ+�h(�]h�\a��[+�mJJ�'{jo	��82'��ɧby�ޜ_���(���J<�q[C�'P�A	���Xٟ�SB�]
[��GN'�3�.��Nm�Dv�CU�-_Rx#En<g��+��ݔ"����ohг��vS��Edl�-uW�ld�>��)b[�.��Ļ�[u��OEi�j������A:�R�����aj�ž���$n;:ݡ����u�r�s��*C��0q�e�*+�N�	=ڷ�3�z�l����ʏ�Ԑ[��f�<�u�\����	:M�][��f�"\b�X�t#]+_uu2��7e2đGl'�mV{��4^����Vf�l�!��5C+�&�t�(���f谺[y��x�Yɏ�v��Ͷi��0N����)��vS�w�s2���88f�Ύ���ժ�n����Fڗ���I�@)'��WjI^�J�a��C0��ȉy�p��Gk�����oY�whA7@f+�ae]4�n�.�Z�����ym�wy�P-m�iV���Z�q�ϻ��a�qԾ#[{�tV6����z2� 0�P:�e4o�ٜU���E��䡘<�	��\�Y��I
 �E��kq/��1��J���# ��ᘓy /TC���%ً��7��"��nB+�[ȹ��wP����ݭu7XƀP5;-<Z���*��K��N�Ȟ�_'�XՉR�{YYX�����Ƹ>�6ˍk�
9�Φ��&gD��uYU���g7E:�����ՠga�m�����-�V��W� /hG�S<o�5V]����ެ꺻�%m�.��B;�B�73����5n�Y�D"��(@���L�͚W/�w�8Ez�}pس�a��ո�0��>y��n�n���aVh��4�&�%��Jt2(LI��~���Cf�%�ِnfkO\���(�DNQܔ�w�K7[�O��']͈z�K���%�h�Z�92�ۂKL�t�ػy=���"��w�[WY-gWn�0��dP9rK�ST���`�R��R�&�Q«K�t���λRAQi;1$iM3&�7PE�-�]YO5m��ckv<a�NڱQ��ՎHhdY�eL}ϡ��l��hb�`v�3mmEIWG�b��ͯ���X�
�,s��<z��h���;Y�x�&��1)��Ja�[���ʋ#�Ĭˢ��3*b�h��\Z��;Xl��M�֪a���RH��d6[3te�����;�r�T+NH���8��A#�f-;
�ϩek�y�-�նM�alf�l�Ҕ]�f�Y�
�W���_͉�b�R����2l��Z�Ȫc�(IGv�0wi�9�F��B�J��ij��fS��[�#��
	����ު���m$ZT&�&�"^��ى�����a���E�w%'.����|]k�v��<�S�q�z5Z��SHaܼ1FI�B�%���X'�Ǎ�D�h,M�W�ue'	R��]nָ�����Ę��wWK[�_�����g���8��3�����H��ֺ6R��ػo�uhV�j���5�\Mn�o�\^L�-�����,��(eh���������KQ4����=U�(^� �4J�6�RZv,�6t�u�&�rp:����#�M��_����&c/!o��Ȯ��"%��b���R��ZOZW����&���2Gj�8�h�6��JRݍ*�yJ��j�ZږU�M��r���`�V�$4������6��;*�2k��$����^]ꅘEV�RF���o-�
S���z��ɼ�6 U�͊�m5�Le,g4��")Qp�*��I�ÈY5t��^�gcSbO������-���3J���m�	��~�-���FU���i�hQȒZ8%9�5҇A�F�kZ(��:4�J�r��i�hY�an^�ݣ�c�P�HQ�ƒi.��ew� ��c�C��&�F<ոa'Y��xD��v��f��0���S,���Ȅ���K}�&c�A�����J8�@�EVXv)_N��c�/n�쎵�ұ{�hj(&v+[WX%��ff��U]��@![
'����oi`=Q��`Z�T����N�:�
�{�,^�R��ղ�X�O;f�,�iM8@�+�,a�5x�m)+]�L�N8�͐M��� ��+��xRv�ʵn
��Ѵu$�۠1�]��U�a�F�sD��bj����f�w�����S��I�)��XQ�3+r�i�����M������TJ����R�ia4�z���H)�˨������!9�cU�5Zt�n�ٹf_���1yY!MZ	ʜw�{��^"͵k�]�tm�B_�nAu$�����Ө�$��[�b�ʥ�����"Ӥ�7�D�4
�% %�6���oR�&V��&9Q�%-�CKf]�q�KA�Y��J��7�Q\���V�+��ܜ��h��ڑ���^�����ˡlf�ѥ����еcp�5�8��/ZNܫo\�
�+c�p�]7��v��8i%���)֭a�4�5�-�X�8�(�Q�˴3N�t�4Dݸ�S3(C���AJY��"_�9����Ǯ���V�ű%��m�i�4Cr�֗���k�U�
ʾ�>JLh�1���^�wRhJ���7�
0�Jx�u�
��鸅Lv��T|����R&ݙ�k��yL�R=%kzS�����	�9���Ҥ_9Ss�';;�ͫ,�7[o([��Y��8+ӄc����
���3\�xʛvbWy	r�
��_�vK�7l��,��u%��7mJ�7wK�4]b��Ve���QP��]��`��+��,PW	P�L����x��qn�un+NZ���G+rG�� $���e�Z�.=��z���~xd���7"Q@�*�d�c)f��G3��x���5 �'-9қȲ�2���3��h�g[�I=pՓ��U��<ĖLŏ��$�8��e��p��xi�kH�D��"ne�j��ն\���[�s�=�i4�(�$���*w@
�IL�sBѲ������@�f�/	�Q��t��D)��Z�#�'b�
��]̌��.�Z��v��g�y�5�i�ė^#�J�hpulT�H(V�j�,T����@�S�a_�aY�4��Lp��]�u�a�����V���p"3yR��V�*��`7T�i�M;�:`]�C(�며gp��/@�wٸ8��[��� N���̛(a��v��ćjVھ�����"^�3w86�7���8Fܫm�5ݪR����u�J�T�
�t�������*1R�r�d�ˑP��^���s�����Zl3tev*YC#R������*��դ�[]#%at�Oӧe&z�
A����FN'+�i�LF��d�D=E.6*X�h�o�q����mv� ;�Y�C2�\[���9-w����Ν���'V��!.�Z4EA4��Zkfޠܸ(l�L�B��4���ޑʵ�ۻ��D�1\��7�T�fl��֊n���~�M͂��w����`	V�l7;(���c���7�kc��p�( ��-)��T4�a+,U5,���4�m��.�^E	�#A�
����)�k�Cb�"���-�6�CM�y�K��K1��+-o���o*	{����)t�Y:�j�p����w��zY��F��W��$�)KQ&n��'�Y���������~�#�����8�pg�$�I*&�W��_���}���6_M��a�.� 6�ɻ���Z�N�3��$\�k�H�I�#}�oa��-��K�m�#}��oyn�="Q$�;��W�f� )Y�[���������Ϥ�����G�H���9�fff�f.�19�t}$�����7�F�II#}$lt���7�H�IΒk�#}$�����7�F�H�I#�$o������7�AI#}$o������G�H�I�R7�H�I�#}RF�F7�$}$�ԀS�ZYa�P�D�YaEl��+����H9+�H괈@�9�%��I'��%�@	$VIlt�Im�����$�[mn�l��Y+���0!BZݰ��-���U%,uP!Ie��"l	*m���)C�S3$�F���ZvJKc��KhZܡk�7dI ��m�j��D:�9��{}ܔ��	:�m�Pa��V�m�J���{�	��N����'��� � 
����9u\�C�蛲�Mu�W�V�Kvb0�V�>��r�_K����ED��3S�P`ʣ�D�}�.dy���>-�y�=u��L��r�`��Z5w�to\�IꞺ�|�'&ۗN�_/���L�7PMĮ3���1Wu�)3��X��<lU�V������ŹC��k��� ���Y=�}�93�G	2ʤ�+U��2��2�f9�>Dm=oE��>F�\�ӕ܎T�����B��e@ә����"S���QY�ho�ĭ�o#
3StI�ɹ:�qhUX�巢�X���wB����Х�e�:��:��B+�E�ۉMF���	�+��6�����9��Vf��9��؅�3�V�"����	��ֹղ34���u��+UA��^)2غ�5	GI���K��b�撅���v"��,��#=Cm)�s���a"01��\���-��wr�L�����Sq��X��)�X��W^���.
,#��/�Ns"����bh^���x�������bjpwjT�w�t��g�ܗy[\���M�������Tza-ƗV�� ���,!a�*�>�hS�e'\yW\���J�S��nl��X%.P���l�Zu�:͹P�S(*Ք.��,J���V��g+:]��.H��g�*��@�i"ӌm��~��JYA�9}� �Ll[+���ӓ��ͮ�5V�N�Q�tF�{��%���#g4��*�"Wn�U�u�r�A��Ao�-\����]��́Z��sɉ	i.I���}[��]��6��v���=��[��Jp�t��}Y���M��R�v��h�%�7-JQ;�4]�[�,\��<L�j"7rӒ���l7љZyws�9nL5~s;������*7^�6�P5i_%��m�.�����4M/&�x	�k�qԳP���5��@l����k!maG�wV�3k�q{A��t�KR_B4Z�ʽ��T�!�yBμ�jq�v�)����V�g53҃& �����sKN��g)�Wa:yE�(;}]ْ9l���J���T��� ʺ�4�ӷ�q�6��yii�/�~y�v.*l���tګ�'R�H`�t������g�h�.2�p��J�Ã�%�Z7��1�Pp����l�f��w�Q�ݵkNe_p�V%xb��T�9WT�kVeo"��k�������H�
R��|�<��JY+��v��2�S�.�,��W
+2��{�ա2�I��g�E�6t!�����o�F���+�N�w_J�($C���\=g�7J�E���1���*��؞]����6��G������fӕP����|�	RܺTn�i���:[��w�^���̼�͹�?;���q�ɛSXڿk���ƥ.W���3�������0�"�l���]�x5�u��BJ�NE�{�����i�!���t�\�:�1�&���?e�z�3���v`K3��+ 6K��p;R��8�����k�t�ɢ�þ�At���1a��KSr�դ���ս{���T��VE��&j�㘹�u�~uf�l,['�0� ��&7�a��͊X�W'~U�c��6�A�9֣t�յ<��WG���8��;6�S.n��{)~��E	�Z�B��kVJ3���*n�D��Tf�0:���{��׊�q ��-���jn֥z�q�J���@�#���5���Q��St)O+�6ifI�G�W��oE���;g�xc�JOE�n9N�A8Hٽ%s�1Ǟ
�יy�f�)^��z��v��4=�TW��Y�A�
�YvJ�r��:��Xx��bB�]�;ˬ
�v�Wf@�#S��|�Y��l��Dv�һI�|��l�u�6u˷��7O�A����E¤%�:����h��iy [�x��"�a��ʛ�q�ے�y-�Y�v�ĝg[v*-�GE�{GX�0���$۫�4xtf6����84Mr�u�
hob"���i��.�gRX��C��"��|/��t�'ۜi��sz�[���-W�]䟗<��ΰ�%���-� �˗��'����ٗ%[�����*�����ͤ�ܘ� ﮲��dg݌Vt76A����1��JM���NeKQ�5�Yx�@{o+�[���#�p�*]��H��h��uݒa/�EM;�~��*�ml{aNwnJ*�Z?��:�ue�MU|�3n�'Dƻ�c�Z�ð�6�h����"����[��,�kEm\�+Mj°Ff��}�!�m�Z{�lm�GVe+��0{��5��%��rbw*`��T�Q��O�ۙ{�k�V�>�$턵�&-Pkz%���;d=��OV
<��i�Ao3��ו��H��@�VjȢ��|�"��M�q˾y�H)�����6�|U�@\��)B6�婊6�:܋v�P���vnmЖ'&a@���x#����饊^ؐ���ʺ�ܳ�C^�Z�Ԙ)��n_V��+��ĕ
Y;�em`ᨗI�F<��Tr��+g-�u���^��%V����J��i��=�L��˯���oJ�w]�{�@O�D��D�c�uj'F�7�o�umEN�]�SbC�tn�Hf�Ȧ
�b�,^�n�~�5��	�xN]}����y����,�h��U�D�֌�w����,xr���+O(��ǎ��[t�ފ�)���ދ�e	�]�1\��Y�f�(ˤ\Rޛ6�fZ����q2�����.Q �*6D6�B�,��)Y%+�� ��9̖k4XF�TYK/.�ݺ�*�P�����MQ;��
Ӱ>��sj	�t�!�d��]��Aacj�y����T�i���Z��uL�$�q�Z��$>KI�# ���?p���F�)�0��GoZ�1Y�"Mۍkk2��	��޵s]9��m�!�[�� Ǡ�WLp�/X.V��P��ٮ�`-=%`:���1$�O0b���h;�¯B�ma9W(�謃����B�W=�ٷO���U�RuP�%Z)l��}�Z���|y8ڻ�H����_1�r��Bp���J2�Z�-˜�:�ǲ��6�hQP�2i)��S\��l��#B�@E�.�Mۻ�q뮱�L;�W��=w\w<qҕ�=�,*�u��2�1��� ���љ[�&��uӼRM���eb��m�á��͋e����Ĺ�8,��bl�f�˭xjs�CYӜh��$[r�B��������vϫOӈ�>�%b ތ̱[I6�������0	j|��j𹗰��c��-nj����b��SN�U��aM��Ӵ�${qU�����?9��� ��(Һ85�]ʻ�0b��qN3 ��}*���R�ڳQѻ�7~�S��Ub�H���G�׬���z�aA���eѹ@-y�q�;����fڬ�J��~v5iS(��ƱU׏��>G$���Ɛ������cv�$�mm����3A��d�u�Fn��{�,�8�7��5��,�ܩ����yk�MV��z��v#�$qUX^^��*ZZU��.���YW���K�,���֘�h9��ni;/�[3Yy�L�ik��S
�)Km�ZCC[B*	�u��,	�ϥN7{Ka���(�x�j<���C�Ӷ����a��f�;%U�r,� �	���"(^G����������h�G2~Cq(���/Λj�B�@�Sh��(�fVFl��Ln�c(��E0�],:mi�j�h��b�#U�~���),*�ә44ꑚ5gd�P�bHe�"�	q(��wcl�I*R�N�τYu�x���UV��\�+;n?�@�쒈	a��J!7H49t!D ݊�J�m
���2��)��'{^��E�ޫ�%瘎I��W�@������ "i�5Ez�@����/8RQ��˄1��f&�h��Q2�Jh��fe-��X�[X	�PF��rj׳���@�o,X�}��l�Y4�����U���?	�U��w��vk��O�_#嚽�\���t`�eNDI�r~�s�"*���t-��f�]�D�sZ� ʔ�,�Ԍ�@�p]P�B��s"de^��p:������%��ٹ�e�8�7�>��H`L��vG=m2���
8���,Js�D�R:��"��oX�it�&���ĺ�(�hl��f-m�Z�h�$|�fD��ZJ9җa���3�C\�m�v�V��g�v�o]��0컣/Z:��sټ����	@��O{k�X��p�yq#����!Ѯ70�V=��?��e�A/&bzE"(�V�� UӼ5���<�ҤX!��ӑ���Ř��s�1!�o$�ő�����+���s����72"᥂���f�U�,��d�4� ���G9�M�Y�y2ଳW(����3�&�7eꑅtP���b�gf�g���(�i\�ꝡ���"�:�ԓC�N���q=�/�wn�]��� �9b���3�������NO=kf�@Mл�8��:kC����t ��Ӑ�b�C1��D��V��Rk������j��^˯ ���[	rB(�_$]!��ab��J���S�m�x7�O�r��4��F�45Q���M\�'�a�w�k�X�r������U�'�X�	H&Q�7�FI;XŻ!Cd�H�o+���`WZ�u�U�h��U�F_��B�l�	+b�8���.����fp�^���b�g��fvox��Z�'!�;H�2�]�U����U;_�+�E ��Z7ULRU�T炬��yd2��8�쨪����iI(2�r�p�v��l��e䚦� �h�u��5;-��v4^*/�`vx��_�e�@e9����U��S:��t�1���'�,0�-�F: ك;=�����b��QI���.����S7E]Ca�D@J��i��9�cڦ,dɬ��>,T�]�%S?���^\슻��b.f�m%LQ� #C
Ģ��9�)IF%Q�N��Q$��.E��
oxՏ�e�x �EC�d�!�.�a ��$�y�B�"k��nH1'�pNeE`x���#.�B��QSϪ�d�<m�EI�2I��Ƭ��\*J"�����U��[=r��oF�:Zyd*v�0�q�K,�+�U	Fv�*���#}x�`��B!�	#���G�t<�l���+O���I��.�<�e�\⭖�r����"0X3�e�PO�WnK����k�� .t��dbu̂W`6��%�<�����p5eu��:5�G+E�kg$iX� �}�{ƛEa��J��^�_���ۨE�3��δ��ݑ�O��6_�ˤX�=V{@m���.~�6�f�4D&�g2�$��e�K�U)aR:�Թ*�(���u�K��:�1*r�+	0�?��6븱@Vt�B�喚ˤ�t�Z+z;�;J�o{�f��>[�k��V�̥�v�A����u�J��z��%fkN�ɇ�����A�9�t�Ȗ�եՈf����]��H=�:�+���;)�W�Ĳ)2x�8��v�*q&�S%�q�4-r���t*���dT�&�
��rX0�����ʛIU�-��4N�k�+Y��Ti�O9]#Ϥ�Φ��;�p��q&�H��f��vk�s�Ò}w��R�Kg����H��1*?Ė��	AKMl�L1;&VU�L��<��ՏB��i�V�O� ��E�ю8Ņ\��J�ڣ���f*���b�:�wFS*�jڬ�i���ѩe�,"�Z
��X9,��`Nk��x=�o�v�#a`���9��݌4����)Rp�Ş��e�S���V�ӛ��;1"�0��_��.��}����i6���|V0��\%����$0~��J`y�����p�k�XO��B�D
T2�8�˚Ǆ=r4�
��T�@�m�B�:`q�7W�eW�n��]�ˊ�� Vi��E�-�j��Ӥ�%)������Ws����XV��5���������1����������Jt�T����BV��)u�Ah�,�څoDFw����xf�8�q�����;n�� �T�NXǓw,Vn��e�"6�<�urP�R�,kά�I�6Ch��1��$`K��&���(��Q����`�l��-��J}3X<����b�0P�5&�vR
�8Ѓ����k{Oo{��X�u,��J�;�+0���	��T[�V�R�Ɨ"����]k�3@l�ޜ�����$���JAI�רm�\|/�˧���fL��{���;��t۝��?&���m��vvJڎ<e\�hJ˝W�"Z�u
]�f��WD:<��ܦɕ�U+g;U|�p�S���FY����j��)��֚���G�"�*�z�ஶ]�5��ƛPs[������nS�����/e�{n<S8���'�ͻq�P��d�;4�G��R�8�ͳg��rT��}f���x	Kq;�r����@U� ���5�7A0�������Ϛ(������~�D2����O�̩2��Nw��~s�ߧ����^`np���H����G�6�KU�����
J�n�hXܖ�(�nm���[%v���mm[�M�p�,(㩦��F׍�o��<-d(����3�Z �E��'��̨v]k>�+���>>�B���F�/&\Ƿ�\p�;b�d��S�R�hKrxRl1du7��f,�'j��4�����yW�H���D�R�Ʊpw��ƸR�g���:�Y�<���[�3ju�i�D��R�������0����8���RWX-]\���g]�,u��P4n���,%
7+0��V��~�|��)iԷ2VbՑ�(L���$"���@�!R��K�Ys�"��aN�*�\zU��N� ��d�rVmC|��I��y �*�!�+ʼi:j�OH���)�=��5Y)�_i0�b���\qYB�	�D�+�Y�H��'�.�\��%�1ց-CW�X�4,B[�"IO�FP���w��j wc������RR�?�d����L�UznP�Ѯ�R���?�[#-ne�R�MR�� =�a����khN�u,�,1�sN&�j%��q��N5����&�qـӉ�t��������D��~������:j�e�#zǕmm9�,ǒ(���&�&����ۗӜ�j؛C�ՇI2:i׻����C$�N�_Y�j��M�	RU"�6l9S%��l�Q?�SH�U����n-nD#�18Ս�Uk.,˓y�2<Q�Bi�ܖ������U=V+��7%����ML��]n���LX��z��*�K3D�3���&��E�^`L�|�z�؄����X��m�[˕7Ƭ�U�qWm�i�=i�;��kU�T���a��V��9��.�I����5B�6�	�u\o�)ae�㙭kT">E��np�Y¶����������i�/�H.�U|�L�{�tB�k��i968��g4^�k���q�j�9ɋ�MJk�N���L^�k����EEBA���p�:�~�_���i�JKD�aY]r��l��r,�i�9�����Q�K�L6��]6���.�?gs�B#��tZ�4�j!Yd"?�! e/�O�`��-���6�\ ��Sn`�����̥���#�q�D��d���'�DƤ�S����1�/:�B�}:ؕ� �VX���B�t1FЧ-�f^r|� ���"�0�;�OO��rdC��ǀ%V�T+.��pRl�!7kg����f��&��N������*-^�� V��K�Y�}��o���9�u�wT��o��������xg��� ������[�{f1]a��QCֽཻ�޵]��v��[EH�'�X�e�������,�����/=ń�>뫦�-os���^c�S�W�e�cö�l��y�#�Q�Ұ<*���)Jx��]��"��E�L+��y��<�k��)�k(�ȼ����䆭_���dZ�}���k}���*��Y�A��x}Y�n��|R�	� �4E�;�C����U�	���t���_w9�R�}g��s�o5^�Z�	��.@�������ʣ���+���Z۝�율�(?r�FlC�X�/9.FzIaJ� @�a6
mx����7�C刞���!�T �Lny1^-'���yiҼ2��>�Wt��\�뫂��Em�@���I�_��\��I�`�����fB����3$����HK�zd����j� �����~��^.�v�\��ފ-3B<��*=���b�p0�n<��K����XD蝪�\;�\��\���r�����gS#4NL�v�#�����'!4��
�Dg-��n�i�1y����?hT8���~�{�ӽ��eb��\؁��!��C<�x�U���8�� |��[�N�(�׎���*��n*�j.�Jl/C���F=�%e�Zj��
���Ǖ�8��4���B��8lY'p��n��;�^xg�y�|F1dகˤ*V�&����N�G�%��`۪�T��T�A��'�LOCwu汍xVyS�E�'��׳1oF��ṋ�_U�Y;(��]��	[�����5x����*|�?N�����庨�71T��W�P�*�ti��h��!�#g�K���;��Ǹ�[EM�3��{��(�]�D!L��|�3����г�uX	~S�C�4U���э$٬⳹�TDբ��44�����cB�-*������3��~H�0�D�e����pU]�g�G���r�i�F�~3	�k�w)Z�0t��6^O���N����r9�(Q���*�Tj=!�
�,{�h[���D���r��櫧�"���^����PS�EV��2+>������o��\�����Vh2dzMd���+%�R��z��][Av����vJ*�V��.����N�W�	��T��ʷv�o�1��x;LG��I�7�x.��ƶϸ���.:�I�zr�a�!���S�.��;�)�s8�$������p�Xz�w��1��R��U���]z��Dj���*��� ����S�%g��P�<�ܰg�} ـ�k\x�翂�c�B��D��_��t˫���G�x$}w3ǉhP�8�ů=�{���0?��^-�'�=a��a�;0��J(F�Q+��zʌ��-.�s{�s�C��c�H*<^7�^��I.�,H_�����D,y�|�����R��3���p�~�(!��#��-�����)СǏ����S-��y�VK����av{_�b��zI,���uo}s�Z����g��!'�$��А�3!�x�q��e�I��3]y�r�������o���|qꬉ_XDź��*�Y�S;�����W&�$�g��LM�и����&yU��&^���<��Bm���L;��@Ƴޡ��}p:~�d� S�Ή5­�ڍn��/�H�xT����i����yƬQ���e1I�nޣ�E�pR^��"��g��<ŗB���G���ן�<��Z'��а)��<7]h�TһM��瑡��;i1m��g�mF73�됡	��k�>�����Ā���c���^�2����L�{r�{
Ͻ6���N1z�Ѫ}��KL�Do��J����c�8ɝ�Ⴜ��#^��ΨQ��b��54zl���=sUv�+�Tv�dT4�ą�Z>^���T��ouy���a3r���yd���s��N�����;��nf�mK�p�\`���"��^<��+�$X%�%c'��v4���[�S�V}��0�{�M�Ḙ���'g����{p�Q�u5��kE3��.O
�Z@N+޿j��bms��^�#�K�)�~�$d(K��P�#�j�}�i-���~�d�ͳZ'�{0QO"��l�&N�{�ã�W�K�z�?sU4��H��j�A;�DW�����g�Y�E��j.��|��Bno=���g���炠�Dg���ԯ��c�.�{@�������9�w<��A�f���IY�-�L�w+��;��G,��;[x�={��[�'�_���NG�,�z�"C�_2���g�?	�n�j
�׺���u{wc�q���{=qa�I����N���p*��!gڐ*�v���(;ڝER+E���������w��C4�)#eP����"
��L�I��6k��	���L�C/,��v�����nL�x�A.��}	(j�`���ș[`�TW�F3>�e�dnV��A�8�b��\��r�Q�_i�>rՑG��(���_-��-�ys�iV�S1K��J��E��<�
-�d���*V�5ktv5�O=�A�zL��p�.a����D:`\*VKs^>[��`𩦻g�&�f��ZB���^w����'{�l�rŜ�ה����$�\��ڒ��;��h�?��F:��N?="���.� n�����_���q =�s�7�q��Cζs�u��wvk��YX"`Sfeo��;��p"�R#x�l��'=��X�9?_-�~�:>\{��`)���;�^Wf�o;�>��g-��R.��@~
��@[,?vup&�b�z���#����-�Y�I�K���s=2weu��in�>�Y�3P���J:��v���{_�U��C��{{z�g]���;>#�^����D=��xp��C�+���n�~�-��I7�y˞X�Xf7�;�`�:I�P�\*'�����hz�ᵲߦ.@��X�W�b"m�=�
��0���*O���vAf���\�
��R�Ȭ�n���c���8�v�q��ز��?zj �;sˏ������V����v|���뻒罽YU�x�Y�pn��W����ӵ�
@�Z+�3���4.��b���Wya~]%?m�Z��;�S�x{�W_Dl�<��-���θ,ؒǝ��t^�tr�f#Y}�3�-r��4�^�Rm1&f���_QW�;��v^��GEL]�M�`*�����]`�N8����<�����b���·�)��B�����L�����Iו������=K���럮�ӳ�Rl�OG;��Fݭ�o����=h_�P@��t��/{�{�:�
-���v��u�q��Ҡ�+5����[ �W��^��:�{޶̹�ӛ���Uklz�է����>��0[��|nB�l����W�ׅ1Ox�F5N�v�Rz��o��;�ᗾ[��iXU�=���[���֝���9�y緳�b�x[��{q��z\����[�"���T�Ȋ��������|�K\E����Z�
U�{%)x��Av�Rڡ�]ln�=S�G�س ��v������A6�����|�F��]�x�!X+��
`�R�cV�����۫G\�n׫)Z׉B�%��Ay� ����;�d��~a�=�����ayY���h_�RnT���*�w����:p����^�F�7괼5Y�P��z�cs��ϲi}�]�r�<-K��\nT��C����-O7�6c�T��Z4.��8RR�y�7Y�@'.�:䜮�gL���rE��1��;�	[�����B��J;6�����,4��짋v�yW�+����N�Hp�>��g#��y<��Cy����B���٫���b(����p5�+��b�ޕ���	����Q�9��z$����	4p�q�m��Yw��r�h����^my�����g�م���ľ����A1�� �D\��g�84g�����=��l��JQ.�5Åb2�t�=m��Y͵N<�P>��ZDz��`�^�&`<�%��^�TB����t1(A�ξ�^��J�z~���e\�q�f/�2�&������e��z,�ٖ}I-��q��:ج�+��[=q�u��f��e����QY~�!��wS��_7X2h��j��嫃޷���Lx%I��eZ����7=ru(�^c��l��NU��`{�|kkĊ���lm>t�ܗ�}��o�1�}��Q�+�6<=���cKP��9T�`�-�^UĬ~ɉ~L����5��_��
���p��U|UwyB��+����Wi�pfڿS�p��a�L�����W
���Ey�Qt�4P�������Lh���)zY�8����k��^�/f��L���^�c�U�#y�+�c�v������|����������҄.�Qs��2s�9ɵ�xE�^Nfvzv��Q�;�4^��u���8G�`ܭ�V�����M���^��]��F�s+1!)�Λ��H��ȁ�x�X,�A�=�Ԡ��]�N�J͟+8PC�K���yi�y��y/?4�d��b����U���Y����R�d�x�Z�;�׃�1t^
a���T!86���P|��a���u��N�����ڸj4�i�ɚ��ء�%�r��ǳ}"�W���r����3Sǋ�)ژp]��p�!S�<g�����ש�ϵ�������G�'��^�>�V�L���k]�V��Oa��d>Ky9w��9��_�����d��fQ�@��V/I=�O3~���J �*�?����d^�c���+=q���ށ�ٜ�Ѹ{��胣��v�`���Ü���P�;e ɠ�	�c���b�Wa*y%�d�����n��y[����3��rU�$;@{=Ix�<}|�gf�I;�=�ݓk�b���.�^��]��}z2���pۊ�8K	Asޣr�M�=�G$D���+/2Zd��A~Tb��׬m��T�~삄�mt���kxM��ج��ɑڻ1�B�~�;}������T���2�+Cb�l��
��N躥=��k�ry���a얶VC�v;�����;SqX;��k��ǑX�<��$�X�v�z*��UJ,Q�Rmd�(�fu��檀L����%�|� �r�ˆ�!�(j�wwR�hla. Ln�/�Eسa��U:�P
�8$�h�&Չ؈�	��d���
�م
���� ��S�Q����$�*B�qS�����h�CJ����r�J�#�H�N�@�'/e�Ӎ� V��?����(é�T��[�2.MV�-0&%�T���=�X�:�-^���ۺ�޵�-ۊ�?�1K�&�
�2���$z( ���(�c�3f�K��8�L�<jw�~�wjW����n^3��g����B�����Z���w����!��G����A_q�C�V(/X��=���Ds��;{Iq3��豞��O\���o܃>4E�6
}�+�F�7�{�������w�||=Թ����F�	NZ�����ܻ��LsB y�{HYY���|̯-�6}C}2��򴂰`۞�$��K��Q�G�7Ԩ6�m�(q�૞��Yk֟7a'/9�,� �K�u_�Ƶ\��ãō�x+��j���`b��C�+�+���T�uCd�<���[�>!�!�w{�7�ܺb�w�v�j�Ec����E}�c�!��*�K��s3}(��ҩ�rԹC�~�JS���<uyf�<'�*{Y4�<l�p�ؤ���w�׈����� !�FSp�W2g�0*�h	
��ow=�d] σ9k�7����j�W8�D��X.%�en�	�eВ��2jt�'�0����۹�u�-9ҖS��*����8.��B廾]v5Ҵ��q��L̮��uu���1B����eF8v_��w��n�w�]�:�'�s�z[ڿv(��ݧv;�-���y��/1ɞ��)q��fn*l�m�Ο�����p�l,僆�Z q��v��Y�{�<]�{z4(�ܴ}�%��phu�龻�?d�x;V���l{��"���u�ª����{e �;�O&��b����8K�Rx1fz��K-ͷ�ٯ{����6�
����+��@6צf��m��iY�~��?Y-�)� ��a*��*S��]���������ݎU���.}���'Q3�Ƣq��׸����7�<֊4?GEo����aοrx{Ӽ';����2��<\&ln)��`�3#��Ь!*n֎����I\��>�-"�^u��~B�(iѸ�~s=Ae�)�sO�4FҼC�H����I؄�Wv��vEl�+�٦��<)��U����^��e"{�\6���4�Xw�iG�G���{��3����0w��ݲ_F= ^���s����ãaՌ�C���yH����M�utD������׫��}H-D�Z~�T���>(c)"?�"2�����I$ �-3�I&��m����:HZ��ǵ�ZV��o�F�r�ۙ�04��?jX�n��9X�aeӢԏ��6�4k�N�"��(zi���[��fJ.��__)���¤����m\��5��\�Y��ui+��A��]��AsEȱ^͜5RWQ]����������N������o��Y����@L�56���1ڼ����U��'���)��F4�n�Z�94�@�iV�TZx彮���s�:�{�\��F� NX<.w3���3����E�,s�Z�R�<e�8�C��u޷M	t�r�g�.���D4���~+<e��"Q�����[[q��(�ơ��I�J�4�@l���ɥ��Ճ��-Եdٛ7�t��f���襼5t�^bY��)�֋We�]�wh���e�9��f�^�.%u���O'WvN�������;�s�� �]���٥z��f�&�7���S=�8�
O��Y¶�X;�NG��J���1�5��
�ݖ鰈kN)�����Ѭi/��D
����m��:�C��30u��9�J�"3�ns}C��0���w.wYr��Z�nvڮ������W%0ı��X�$�����o�v5=��A&�tJ�eK�ެɛ��m�Tn���#��n!��P�-v,ٮ*�°��%n����L�t��C���uHc3�/�]�0�Z͕y�u<��^�ˍ#"]}y�KyYl=1����OR��[���y£|{7J��]�q�& +���A�S�`�+�^���ܑ�Ъ�nuD\��f&��J�7Qٹt�����l��;�.;�Y�VyV�έ5�X�]M�1�V(��i���-��v���.��S��ܯ�@�U�l�CV.�ݠi .�v���ʙi(p�o�j���1�Jl`"G^�+�<�Z���r��Y�H9�P��1�a���
P��n�lԚ��9�����x.�%D��8E����Xti�Q���`�*~��(�x;��������>��
�c�s�u��*�oȰ��̝�4��:��ޮiG�m�p�{�.�q�o;�%
�ׇ��1g0E��'6��
�
j��-mL���Ea#�q�rHC;���@�0�%q�om�w>��?L#��ʄ��u�кgIp��e1��R��]��ٛt3EҬ
8�u9VR<f�_eVw?�I���Y�"2T@����I��#CCH�~�`"�� =L����?R��E �#L�RDcG!	�� a IV�2��2�)�� F�8�QY�1z��|����+�� �� �޹���$D�`N0�!G܃"�"�%6#��˘dB#�B0��4�0��,��F ���`�|�3Ρ�L Le|c����3�Ie�"���3s�|cL3�teg�����$������@�(�FH�m���n�(��̚1}�8��F '��,@�Ge��2~� ���$��8��ŵ &��7}/�u�7��fPex� �F�2@��L�� x�ny�0,�;�(Ƀ*!b # �|C1f!"H�8@�N���+�b�ȓ%
1&$���`b>1����# ���S_}�b�ܝ�E��ۻܪϨܖRФ�9(�vT�k����0��~k�j?��j<��U x�1?Qc� �F� ���H� �6Y�@d���O��,�DПz����f�]��$G�"!�D� �0��!��H�F 2:ߐ��ş_ؼ@�ȉ�.$�֡�� F8�j	�@YM�
#��
,�}���C1� ��7'w�yU2�� q |QG�*T ����@
�5�`O��0�I���Y��T�g�ޗu��L�D2@�	1O�4a�c)E�!����q�b�j1x���|��iFm �	��!�`|a����~1`_�ńYc�jH�P<EHa3���N��wo�]Wc�0�H��|G�E�	��W��3�4%��ɆE�$�f>^�&!�DQ�����0���Q~@Q�D � ��f&:вY��4��҈f��I�@��]�ӽ�\K�Rs����	���X ��"$�iB:P�J l�p(��,Z@�@J]�%ݸ�4`(�<b�dE�3J#l�D�a>(�ok��/)��R����
�N $ �5u�cD��gG�H�#��;4��$р4��A!4�M|gBA Eg�<h�K@c�'|�(����!1F4� �'�}B(�&�f:@��v���H� ���Ĉ7��+���d�u�3wW쭰iO�5n�[�˨��,�YW���)�uZ�E��U���ͬ�; ���V랕��A��NdeOK�\oY�o9��#��<v��fT-l���^9�I���)�Ůν�ETĘ�!�)	<`I��գ�F�d3`"<�U��rð(�If2P@�� LGmL�1Gו0��HӖ��FD2"����4����>��_��8=���rB�`jXD"0�Y�P�,Y�H�0"Z� Lz���@DY $��@�,��٢���ş��)VI,X�\��#��s�%���]v�	��m��/��K�q�_���ߐ�p�Y�0(�����an�Bf	y&Tx�"L�q���(��J�� #j��1�!���"�	2E�k�;;կ�>�Wu���08��F:TI�	�u � O��,���D#���h1������!����l��� L�B5ƚ0$�(�R�a0#�_��t�1�K0(��ޱ:�����B[ޝ��0 Q��Q�!�D�1�؆bZ	~"�_!J	@�kd ?!�C Y� �!F"Ȣ�����ᑏD�	%}K�~._�j�_n�w�	��0��t����g�&nܮ Q��Ia���f<@g1�h��"��(���������C"}R#�aF!@�	6c�EGF�|F�����O��MDKf�������(�(a�1��Y�C�`#���� q���$ �=�	���q�y���	1�D=��t�`3DWە��S�hΈ� 	�ő�g������ݘ���$�#����ה&>��p�1��H������Q�f`x�?��a�Dx��P$��"F(� ���@��2sx��LGyC kQ�F���y��W�I*u�1�A c� A� # ː8�$@�@F�m�3],�%�_� @��� ���E��@Q��`Ncd��)hI��ʈ�0� N��HJsP����f�W��<F�^@@�n)��DGyF�D∍0��f��$�1�� �(g���i�Ꮘ�&�����Yև�x�1&)|&@00�(�~@<PLB8`fZ����U�u�s^*Wȍ9��>bq_*�}dv�5���dZI#E��C�}O�_d����VJ�5��u02H���1�˯ϐ�W�C�Cb��v�%/LW\�������˒��X�!ucu�l4�{ ��"��q̃ �F���9�dXT	@N���
���n�:�R�e�rյ����!,�,�X����-ՙ[�L��:9'�yb����Mc��h�Z5'�;Z{�`����+�*侫s#ғ^�x�#��ʝ��q9�i�fdFQ9Q?�]}i!��+�9�$|t�@_y�� �"�0�KAj� �@a�)0 �L�G���1�@$W"G|��-_O�����0� ]�b1~h #GԠIf-�3XKԘ����s�}d��7<�$� a��|�@�$��pF $8hr�G�@��s/��"�Q�����9�wI@F�#��0�D#$#��Q�dx�� V����2H~ 3��s�<.�?N:�f�� I��VLx�� H��#J0$4 Y�W� "1�!�)�&<c7x�d�D7����H�M��/�*kCh�M��>]r>!rD2�C����⼧O9��ުO|@�W��n4�/��+A������M�rs��>}>P�t�<lEE�+���r��WNĚ�̩�U�m�F���Sp�2��>gE�훋�� �ϞHҫQ��Y>����K^Su��.�Ò���N����w
#��X�C���\>9���S����y=��W����\�~?���ΞcQ���_������x(�ĕ�������Ҋ�ު�DMM�&��=�碴�@fOU>�ͨ��@tם��=�'��b�OtK�#�aU�U�۹���`���<1��|�b�쉳���O�
�H5E�h�T��ck�_�i����̂���Y_o]�XO�B�c֚�V}y���5{m�x�5�7fڄ!��h��j�F�������ϯ�}�����ߧM�Ib1w��[C�2�Rn�w���^�_[�k��Yޟ=�b�^ĉ]��:�Sc+)i[	h�nVǪ]n-��j�;��Z�j��B���S�ng����(i��P�B̴Y��,f[|	����,U7iu�)L}�#j��� 4��d�zGY���e.9�j���nz��u7�G����{"�����Ѵc���׹�\Xb��bQ$��uZ;�rE�L�0ѿ!s)Я5X�O=���W�\��)xty��b%��ڃlsk��}�=��yR�������o�
<ˣQ$i�"�+ľ�N�4]�ſ�惟qoј��~�p�y����Gz%ʠ�����N���*�k���eϟxd�,�lm}5��4�Κ��;� c��o�w�1�:*��\MG�io����!�	���1�ܾ�3+���ENBg+�Uy�kc:y��J�Ż%}M����ZDÅ~�>L�����i6��9o��.��XT��,��Z2���s$y�����\�]���'�RI���Q'�T��_�ۍ�S�C�;�}�s�Ļ�Qq=�5Dk��^:��[)_�ʉ���f>��ע�p�S3w�z/�=��S��'����"7�I��"EvZ6*+��{�6�M��c�S9���J`�Y�ڍ�M'����Ol�� '�s�����qخu�G��p"{���~Y(��8�J,��u�2�i!5���cR��>6�a��Y5��f��V35��Ol��M���uT3�V��ރYtz�'{z�ت-����JjA߳����sCC�;����4BQ}�E���o�(�{!�]����Q�]��t��"��r��ux8V���61���̢�64���C�xS�e�R�,}ũ���%!a�Z�@:���>�蒊�LIb`�zbb�Z�Fƥ��*��J%����d���,�n�A�˲�.}4\�9���T)jڹ�*��qW�����^X�ǽ��F8a��L(�ׁ?�4$����~Z�{,/��"�a�xg�/!��"��W��UHv{�kO wf�P��U�hdo�+S�CO�5�O�;h��=�02ג�K�����.F�AVC�*���TD���+�R�G������g�&8#6�5�\E^3�s���Q:�V�:4�y����m[ Nt��e��Fxi�>!]J�y�M��z)7��i�%f�3Gl9a����,>/�P�˹��R�9J��s#f�NI`{"<��ɚ�Y�~���;���r�JNr�8�X��.��0��;����=t��&�n�`�~�/e^�����vS~��:>XU���P������3���^KỌ�l�HOIq��fV�VC�C�&c��j�a��z�/�|!N�/>�Ȅxl7:c)����|+�F�զs��S��N���"_^�1�`�x����mN��4����n���i�+vu'����S����spa=s�Gh��n��M�z�"ʨ�"�I�΄V�mn��d�,�B��g�噶����|tAb{�_��wg��kj��VZ��L�\��y���8q�=�^̙F����>�ng�\�qLsw�apr\�,�����y��]����3A�.}fϩڝ���6�W��K�]���}��Fl�.;��4�M��� �+��\����}N3_e"�OZ:~����sպv����j��U��0��ɪG0O�?lN�(=�_ݞ"��x��!_U�'��
�w��y��If�ʾ��_*�U��(��W
��}���WN�
$�h2lt�� �B�R���j�`�W���/h2����~����8R{��*E];=r{�=��ا��T7d�u��G���Z����6�ݼ��RrfV�Es2��ӟ�E�J}��~	�����'Ӷ�\��/�{��/a����ػ�|�<��QW��m�0	��g��S�-s¾BӐ�ur���z���Ex��\��=V�t�0<�	�`� ��jv��z�	��3�9gd�A�{����s��r~�*2���\Q�K�&r"���jy��󮬉����U��d����h�K�9�E�&�-�z�bCHc_yf�}�v	d�vbV|7D��W��Ow|Vc�����L���bc��{��2�md��r\]d�>���k�ȶ7����7���jы�i��e=�1ǎ���]��,�Y.�fw��o!O0eۮ�J�GJhW��G$I�-s���U���'�kf��|�-�~�!Q #u�G)��h�]�lh�m��\�r\u$�R�0q:I�JiT(�7��76�hL��ͤ�Ih��f6���F ��sr���m��Ygs�ȫS�9H��i]�fs��WL���
�d�,�k��q��񷖦M̸ʿ����==���(+/�@�����c�X�;��wF�SU���E��D��޾����S���j_M�6em��4�"T��w��X�Y�7����;m�Y�t��b���k�?#��Oyh۹c=��X���ћr{�UK�kꏭ�SN�բ�!�S�	�����3Ҙ�t����,i��e�1Wh$�C#����!hǳ�K��j>-E	2��Eto���u8<*d���v�q���@!���Eu���&��eOy�"��}$9p�ێ<h�P�[��B����1��]���h�D���B��ZD���@?w�u3.dȒN?�W��\���{�;��8�P�Em��[3�r'�a�T�2�{1X>��\��[��T�tNdQ�S����ɏ.���:����̔�rJ����ܳ�$�S�Tv�ׯ0�SV#"t��w�~<������QI�5)���8�NMh�+����ʲv}ӆ��GX\E��y�]�����Q�;^KD4������
R���z�r���������P0��%#x+�����RvP5s+-����Z������Ogۚ4�X2���} +@.�N�{�b.��W�DK��z������iP�
�RóѾp�O3.TCˌ��"��q'd���F/��\lڡ1�vX�RH9��μv�����Cwd��
�K���̌�Z����\3�����л��B޼�E�KY�˺~x�����:�鿄�T֢8���WV=׊�q�ݷ��]<S����+�mp ��%�zw�K��vT��Xx�/m�Ux>�
WP���əQ:c��3�����=��=1��?����F?ϧ����~��'��?vF��NUM8XQ4VU�|�V��sR��\��ľ"�琚�M���6O��.':^�N�j�bv"-�+�3&vC���UeRļy?t#��X���r�s1�B�TW��QОdQ�vY��7�MGB�A|������-�mR��s~~VlJ����>�,5��H���Č���z'H�U���lQ��dw�ߗU'/��w^�h��~��"'�����&p�`a�xs��O��Nh{��c�Utlߖ����d�{��W'�V%��S^i1��4����
�A��l"I�( &�M}gkwײ��άTߐ<�j^{D�;��k���K{^;C2D�oT+��scNz�wO�v�m�>���zOg'S}�O�s��
���?�(��	����
o�+0���#*�+�ؽ�VZ-}��5�>~_u�P��XCذ��2�����exZ�������Ӈ���V���Ok�}O�7#�o��Y��}��_~'F��������:o��ӵ�.+�h/�Q���L�C�mY�A���q��!X��"/��P��aT;�~ꓡ�F�qn-�]�Δ�*�G�Mw��u`�Zհ�����s@qo����=����q���K
�}:��8����aVxMU�؆�^�����%{����K�Iw�/f�J?W�3�v:;0x����0��	��/P��.�Ӽu{x7�P2z|�*$��gb-���/&����B+�牃S�H�/%x
���^^0"ȳ�u�;���`T&;�Jɰ"3�!�[��8����^F�%g/M��rޭ�q3�h�f�dgqVs�T��4ugmA��{>�6K�[~���@�kҞ��lj���v����vH36K���br�����W�VӶ;���?J�4����ƞ��]hk�e�h�d:�6�:j)9������GE��Q�k-.eoԤ�c�쑛4�,Y�%�__� {�����1���~�>�/ cPsU����������>܈q��y�YV8G�3\)�F�Z�P���3e���/�����ղE�D��ss�_��錥�J��9A�q����~1�l���f��jV���ְ��&�_T�5�)����t���%��`i�qC��\Ϸ��+ � �t-
�*_�U��[��+�*E��"����#�R]���'��[i��>2-��>� ��3I�nb�|������k����|7�YßP&�g�R>o�b��uy�H��v<k�SnV����w&��/xc뺳2�jg�ٳz���n�|:��
X5�#u��mݻ遞�]�klq���Xx�ۋ{�2�in�5���ۭJ��3c��(��Q�M�Ӎqg�J' �<>��޿LB����~6����(�U�����]C�f�׷'���}q��9��P̱ޟHѮ�"b���P��@/��H<���毙�1^_�$�^08�m
do#L�*nԚ�H�T�g7h�Ѐ|�����o��9��N�����>�[�������<s����ï�G���2�&�P�𨳴Y�9�v�x��E}��?<o�a��K���׆�=�39��ez�L�"R{հ;�ts�t'.�vX���:��q<�����BZ!��J_F���`ǌק�\T�7-��M�Q\;���*��%�]:�!��n�ܔ'|���U�٫���e���&(}˩���]���vgĬ�fS`��U}ܻqn��â_P��_ڹ������7 ���t����N���G�o��!�8�^켷{��=X��W\ϻga!���x���1q��&���i�}�L+�t=L;��2gU(	ˠ�t̖$�����~�@e�Ee@�8)}Z����_�F�w�'�\V�}:�C�w{�����m�<��!���ìt3}=�a�CzS�aB`�!��� � __��{;���7sDN�AQ-.�Q�T��ua�������Mp⭍:���K�VX�wF�a^�6:阷��K�u)N�;D\�ʂ�f<�v��7�".��֔��Zp&,�v��t.��%Cq)?szu��4S���r"f�:ۻ�br���r�';�)p��!��}"[��v�<��H��;�dҝ�W�m!D��d P��վ؛�W��ht�2��F�	WF�n��X{��C��tGZA!M�sx�\3�lm�֯tݕ;DN��6w��@��:Zd\�� C��\/?p4)N<����R5v�Z��I�Kް4
�m�m.��^�]Xn2\���j��&-����0L/z[��Jb�D.�i��8�v��7�;�]=�� �^��8�.��	��yv/�x��쇦�AQ^̫T���ލ�	�fܸ��[)��r�ͳWZ����d�ޒY ~��
0�Y�Ӽ&�V˹�}�jE�#�b��"�;7��]�'%,��]h��T��3��ȥ�yj�P�Y4
nL��"].���L��o]B�Y���ȫ�t[s	��ȩ���K��]�W�=�E���w͹ǲ1Q����O.h�y�l@^����Ռ�ܜ�>q�ј�}��iQ)fA���z�����Z���hk�n�=�8#*
�K����{{�s��S�z��d��M��a��v�` ��м�U��t�l:�����E�݄_D��vV�I��Ղ{=��K�sҎ�s)��le�ᛄ&nN��$o3�s�l����Xm�(�A��d���T��1[I$"p	aK(�d�AT}�s%�" �QV�+@D�O��SY���E��P�d0�c�m�5)�j� N[B�V�`>�/�V�N[7�RC�q9�V�pz^�j�`�8�ظpiͽǒk�s�e��o�L��ٍ#u�m>޽؈rޤ�X��j�d�{��
� ^���,��;��u�)�4HheL�ږ�r0R�Q��mD�4u�P�],O���Re��+���|��:O! �'�i�]Zt�C9{u�q]c���I-�y`�;^@p�B�S��iL�<V-���UѮ�p��S�K	r�h#|dH�˥N�e#m`Qg=�Dep|����� Br-2:����yi�Y��?hըQw�#�]��]ે?iB�������M����R����vF���(�o�6���Ig:��U�t��j`���j7��ҋT��ݙ��g�e֝j��r<�0�v�[>8�6խA˰*JjBr�tؖ�;¨
P)���"�rJ�I�]�j�++�'@�Mj!�v�E.����ơ-�:��)�M�]�	�]�|t`+�*�qoK�����6�mr��$z}0|�^�(����K�.q�X�e�ظ�U�^5�2�j�OZ�:��Qg�W�Qh��0������z�v�6�q� A� b���شf*֛�{�����'ծN���HT�ˍ7Lu�#4�(���Ec�YjH��aMұNS���rB|7����:ɳ9�q��Wl߁��Ց�y|vooD�h�lᗨ�B"J4ҽ����m	�g�3I�d(&`�ҽ��W3ي��!�d*+��sgfz�JU�ȗ3s�f��
]�2���J����I�Y�s���W
���j��ۚ�Q�#:�|��uf�Fn��m&f�k2���Q,˙b�Qi%��^�w �,9Z6�M����/�|2Z�X��!<I�H�M%I����lS�a���]q.x��z~I�y ��ڞ�j�t���̸��Tt�0ś��Ɖ�d�Zx߅m��K9��ǎ�HD�	�f!�e��v�Զ;-��ݑ�����g�i5T�0F<oO�D���)�(;����OOZ�ʸ�:�-ڳLF�Ԋ�����݉�ˎ�+�ێ��Y78W��HBs"w/=�����pw��گ��Ah�n�U���3��G��Kײ�g��C�k/O���=kʬ����fL�#��Ige��v�:��t;�sF��+��DFP�c�)�x��k|����v�z�&>��Ǉ��ԅ�̈�I6h4ĩ�|�r���Yb���t׭�6����k~r�q\���nYQ��'"g�H�#��ײl�ٵDGvK���~Hu-��vꬮ	���y�u��{�d@{�X�b����tѬ+>�]jrY9xf�u���D�;�����78E��3PjM��STE5,z��@���ֽ�������u9v��qN��f�z&!=<����?�>����Pk��<�f �2�Yy�c�D���C`j�J���������G�+p��z���o×���(Pc��}�4e4�^5��ns�3�.����r��O�@l(Ǫ�o���z�u��X�ğ}6@?p�j�~�2����#DR0�Dc-D��a��Ў��l��"-�T7�z5�C1����`�������wI&w$�$�Z�Ր�`�!gTӻ����#�s��V`*;r��0���w2;�"��9�hw�f����wmv��t0pU�V 6�ܬ���j�dc��:���՚�9�%Z{��6�����̩lۓ��h�r���1��skm�ba.���o�lЭ�:�T� 5����z��;�|��H_&���,e���.��̲�b��̗�ѿ1�e:���u��}�O�˿��쾮̺#u��y^��<cgf��z�����U�=�;��+�I�О�����F���:���bݹ��o2�]{�}�b=�����{������y䖇d@��o���ǲ_�fq��v��ݶ�~~�Qߚ-4OVi��8\����B�M���v�����#a2:���NI����H�]'Χʈ���G��q�N�z��x->�[[�a�˙��|b�/�l�f�<}�/�&���YBq��Lz��ۍvm��>��^*��|�/}��}�q>������7����WS��TU��]�D=�E�Ry���>?`%�t�Z��}'�k�-�Y��������ӽ��DB8���+%���B��UE�L?Š��hH*&Id��G쿹���Q���|!����y��P�W_I�����eŭ]�~�3�<v	����O���j��[�q�]���|/�fT�@��Y��C���������ɠ��|��1@y]��0�A��d�
��F�~闼�s;��֧��/�a��Yn����sQ}(I�C��;�e���#�����w�����^���5�<~�!�#��ތ"��9�3yX��:�!��GwC�w�	�QR7(G�D��k�L@�f�2����k"������e48���`67E�2�>U���fW
A�ֹW#�+�]Қ(V�Яn'!Xv�D�h�ٛב����m�j��e��U���l�ᒣB���Ҋ�D�Zn�n��}w]_pAz�r��-F���� �Z�g�1���G��2�_�=�f ˣQ��7�
�d>^�`���)[��ؼ��3���Au�������ً�eAT2V����9/�h|[�u%V?b�B?��������������y46��=�t����,���&!\�=���R���R_+bU�xa�~�7ƺ::-N_	�J,w/�z.t(�ٝ��F��6�%�����eЎ���WD�+4��M(J�<x��7<�u�ա(���ῳiB��"���2*k����-���B~����L]�����v�M
�d��h�F^�8���՚CAv<s,�{��#fz.p��T�hEǢ�a��{ ��V��1�x/	��_p.2�[j��Wk����@A�ޫ.����#v{+�׺B}�L6�����*�{�5,̛V���`^�X�}G�<QVa�B]���YV�t]�f����������OU����k��^����/�3վ��"�(,x�o`�X\0�/g��hIh�2��}x���tJu�c�:s�U�\}���׍z�k��/+�y�׷���)����#��4Fr��3�U�0X�n�T�W�{�xْP���q���|���0�����G�5�nv�K�^�Y�����'��/h>���v(�� ��n����[2WKn�Fz�	Zڑ�v,s��tI�qh��͝��xgN�e�(�eI 	�ý��k�������i��e��	]Q��*�Wc��7l�c޻��3������"ܺۧ��.�>�� =Њ�^��.=�ql���e��۞v���Rz��_h�Tȟ`و������O��̫�5�5>_{Z��r@�9�?O�
�5f{�P�P���ш(��C'�+��J� �21Hb����FK��b��0%�4_䇫����}OH*���Vq�!L+h+ۜ~X��d�ڜ�=����w�юU3��������_k@� �}�S`)��yD�yXyo��":����(�����YD���t�Q#�[�c���ׁ��F��l3xM<U�P�<Ve���\�[P1�F�J0�#�nǑ4�^���	��⚏�:��n�Y3]����	�w
�3K��֕y��z���w�Tk�@U9��њE��#�%�O
`��U�{���g�˟;��
oT��m��� ���0��%ݟ�e��ƶv�ё�������Gw-C�.��С� &��T}z�!���3�
I�W�����́�<��,(�t�O�!�>���"U0����Ԛ��|gy��7X�=[�b;���zfx5b��Jc^�� �x>���m���ǻW�Wk|y�v�gn����a,���VS���1<C��l;䢫R�JR��^�훵�f�Ѭ��ؔ��|M�e�R6嵃-���wј!� ݩZ�����a��~�we��,��6Oe�(A�.��;uE��ԕ�i"�3&`��J��X�WQkŔ8����H�cad��L�cȲ������S1���r�,��Tt8���V��7�f�(i����	���܍׈dLo+q�D�v�'�'��#y3�����x��
.;)ߴ��|�y�1Q����Ϣ��Mz�
S�l���hӵ�*n|c|8��_j��u����V.<��  �̑8�0cz�KN�N�n5h�-�3�P�4�]�>寽��Ǝ���}q�(���mR�:��|�%���'{&��q��y��}P����]%�q��F��$�}�j]��"ch.�^���~V<�#�?mߺ&$x�D���c�Vn���u�GD�gO+����M���\K�9�$[��]���������������z�[�ͷ\d���Y���7�M?+���%�u��g�F�l-!�3�{��\�W��w�=Q�.�C�#���)�fRfK���vϾjL����"���xM$Vx�.�w���u�w��<�Խ��,��Ef�¾K6�(V��®�qdS���Wﾾ�ҭy�(�H�4Y�Œƌ��+�m��������+VC�ҽ3z��2�ï���*j&�(�E���G{=G�#��۸�3�>Y[���Ծ��\Ñ|bs��>_x7%w��g����M��F���ˠ\�0qHK�;����|�/�MY���������ǔ�}oJ�M�ۼ�3�39p��ŵ�W�U�ץ����o��e["���gv�R���̸��jp��%l��1g+C�I��u󛁣7�u���5��_="��S�Ǜ1<����V��ӝ.����y���g.�~����0�f_s�6�m��p��|�c����%�5���T4���na�q�kg��������yY����Q��F]Q�s鈂��W���r��=�oÙJ��Y٥7�G�a�_G�C7���ĸ'uG�+�6�{;t��#=�b$R�8��# (��~��W�Rq^^�����.��)������)�;�rfa��܊�Yx��^	W>-�<���)�,�%��d���_HvJ%����<���`V;��G�Y,�\A��w>�G�	qU�������UӠ�k�y����QQҦWM���o/`v���쨸�ٌD�}���.�:j(���6�c$�����[dX����ۛ�u�Fb�?W�:��ὔѪ�w���N϶�~��HU����{�̵m?^g��:pU�[ײ��ٿK.��@O�l�]m��U��r4D^9}"�T�͊]���//3׎h��-�_s�-a�իxfl������LT�ͭ��f�U�J=��O�㪤�V�{$�Z��sax7��{�:i�� �^'��~���雷wu��9:���*=M�vx���0��/�b�$<7b����*�%�H�">��K}V�⡇*�O��K��j�[B�ɏ1�&s�2�(˱��g�no�E0%�M�Z�\�s]�yv��f�h�wVRh���{����}��:�4�"�t�p~,�Ϸ��RR�飝V-���2}�d��Y��Js!I3m��!>�k�)tz����>�S�"��B�yqk���S�~���/��Y���ۺ����g��LR�51�����S��;�*���y.�UG
ij�x��m��:v�"g���S�s����|��*��Y���?,�"�Aj�9N?�g�L��^?w��y�u�!�1ۆ��F;"M�ag�
��d���wA:z^?�>������}$9�rk^���k��=hk���6Mr���9��C�����/����:���R^se^�@ǥ��zv@��:`IoЇ�����,o2�NS��ڈ��V��%�V���:��9h�;��U-V/w��11Y]�ٛ���y��U�1�;7��������H��gҋ���"��p�krj$:غS�&{*���q۸�{�=����W�;.�kMSy��}z�+	g*�f��ϝ�=��o}��f�l/(�SP��-4(DHAq�>��nS@gkc�ح���\{��P1ގ�zo�q]s�_��"ld7����}~������_IU���X|;�b�L*w|�����}2��'�-6:h<�-�F�G�~T`��Y�#yrb[z]A[Ox�����Jc�-i��l�+��Wm���sa�4^�����]�0w�6K����7�¬0�۫iR/��I�![�^^���S[��,�uf�43��(b���d�o=w�u1�.�	�1V<�z������X96x{�g������f\�C��(��rUA��j��d���k,m1G$�J��׮ �B��2��SmSR��zÞ������=���/v��g�h�.�냦v�o���CK�F��c�Z8_��׌���{�2������Q���|�&���~(1�����)r�
	�t�ˮ����=�x�֙����#�����|E�.(��p��H��3�+����+�q<��E�ȋQ�6��н���Z��"��C�����F����fk��
������,c����Z�&_E{��\WO
��!��<ǒ8�Ԥ��H�t꛼���,�,�37э^�����f����G�=�#H����@m�7W<>׃�x�� `�U`��٧�����%��{�.���E>�O��ɀI�t��@�}����S�]{cH�8�i�����c�!K�h��1U�65߬Ρ>icB�{��3Omm�q��R����ׇ�[���ǃ�Ů/�Hwr��Qw�~�����Xť��T3��w�<X����bʷ���!:������˨v`FE�ڕ��.뙏b¸�j��3�s�b[z��X�O�J6�2Am�ժ�8�f�UakC���5�U��O
B��Bi):�2@-��ߜ������8��ǃ!�eL�l�I�TS�a�C�c��0 �B0�/�ӎb��+CD	]S�4rR�#F8�������}VF* #��������`�;�X�#���E:I�g���
�Q�n�*�1�+/�=^��q�5����c>�wk�%�������֫Ҙ�������r�K�,�_O�;U?����*�p�#���gĤ*�x=��.�������j�sS=�p���E^6����4��ĽM��7޽S������/�^[9+/�K!�/36_c����G�k��K��Y������ߧ$<�c>�c����^��6vr���HO�+��v�sh�^~m���-�Z�;����U�|�B��@?A�!�*��L��d>)��/h�>î|�f�dB�a��US}���8�C����<�:G���潝��r}gbT'��Ӻ�m�@��q��>�y�����f�#�.͉�O�*�-H���F���G��7��1��n�3�[���5\��V��b�ˑ}D�k�j{'CW��{#$E��=�TzI\ͭ�&��ȅm�RJ�^1��XeX�L���ɖYo���G|rov��}pm��s§���mW�U�魲�_k�4sK���XSy�����ߪ_���L��\+�����њ(l������J�Ė~w����!��fg�XWx�ؖ�7ӑvj8���8��-i�˲(�zZ@<�3/q�Q�V�_jQ��aM�X�Jw�R{�Ζ
Y�۝�I]Dd��}G����yؑe�F�V�9%�ӳks{��=g�j�wնymN]�^=յ�ymp�R��:�������x�_!5�����\c��3OҤ�a��&ߺ�A������B�;���ܧ_��v	�����ΐW�WmE���b>j��C�����Xr�OҾ���r��5�To��e̪�t<p���D��.c��U�����=.�%G�TyB<��V�!C��n��@�yS���ׁ+ًù�n(R��3��^��g���p=uT�}@]�iL�13*Pfm[<3�E���z�A�OS�tC��\lp�����I�z�Lk>�G��z��l.�QZ&}MHT0Mo���Z���8a_����=!�|[�'�Z��u���#�Ta)�kS����ϯߌk6�S�?�N��E]կ(��]=^���["rϪǎ\�vU�phu2�myy�xG�y����l��n�:��)���po=�:O�F��~���|�5�ZF�3m򜙛7�+j"���Ց�LL�U/*�|�O�{)�e*m���lS��������ܦ�O,�7W�]?n�����g��GϾ��m�B���З�苘�?+u�S�l��d@���=������ �,�]����C�wY-��(r=�^fF�r���r�t�:2Q�;Z5
�:�;���
r���W�$6���N�����v��I�8_qa�Vn*�/��Nn8RT�]ZWU�=�C�}�>��1�8��P��r�h=n&���Q�!Df�cc&&l�O��ذ	���'�p�ҭ��\��wϱ�+{f�:�\.��������|�K��+d��P�V�ҽZ��C��JM�����L�3��X�V0�Md����vX1WMe�>#�I�c�*ZZk�Ҡ7��diJ���If��+E�Į�Μ�޸9aT�b�u�qX$�×5��]y@ܻ�{�� @�=`Ό�(�ݦN�ѡ��{���n�n�9�E{��!Dp;ݰ���͜�r��zd�0(�aK����x+bv(�.��Wӛ��U�V��᪞Wd�3��;�&���aߕ��c�d)������Ҹ�N�͓�B�oj�������+�i��/�u�qu�C�%pA��-��b��M�(:�o,Wb@1ۚ�&��ȷ&���%I��6T���$���Y�7��Z�Ր��ĕ��/\�G:�j9������ۛ��Lb.r	�	uuٻ�P�ֵ�fs�x�-Q������i>��s���,Ùu�l���R�d֑
�4��2�]�R�5h��v���XOP��Y�g�����#�.�2	����}}5: xNvB�0���&T�x�=�v|�kJ�t��83����rI;�IZ�Ǯ�^���X���ɦ;w��M�].�&���8�dWd{8v6U���U��vi���R���3)���Q��(��vM����k����FC��D�i�Y�/z`m�X��	�����ܹ�ܱnN6���er#�A�w[�6	��Ym�qU���/�fuvIv�z�pO�u��,(���Z��s��ݎ�ٱ��g][+�XT��*ܾT/��q����#���h�Ӿ�q����w��)N�Rb��γ��B��r�����+&��!��F+zu��3�\��(��Qv�#�*>ףU���,I��EcD�r<�$��y�M�h�*�~?���Ǻ�e�=u E9��{�3�����b#����־T���|��į8�k�3����֎�W�ߘ�.�r.^n�w�~��Y�Kg�����ֹnUn��9<G�<�g��zu��a�0���i*�{�M��_\�U<w��]S������fL�U7���[���n����ӽ��\.3�5	w2N�����)"ǹ��۸�0yb^^��R�3[�2��'��{�|��Ƿ��;�c��ʷ��Y�C�m�Kê'Q`�>��H���ǣw�7�\�::8.v(l����R�G�� ����=��dj�V��v��P�$��L�����Í������Y	���sr�i��Ծ�k�ZP"�z������).F�T�W��Jx���=9S���AS��0����:����6����H�,Ltz��䈫���=�i��	������ߣ����f��+,oVf ړ]���y�_9ı{��.���H�6=׾����V��t�f>�% �5+4�HgV�?}�[F���~߾������ ��^�?<�$O��bJW��w�fdG�����:���Y�c#`cg���6������wn'f�@ܨ�j�%g(��<xPos~�O��z�����p�C��Zc��`	�e?%b��;�l�mfzc���~��'[ ���g��'s�ь�G��ɔ�M]KX�|$��uWvkB�e��b=%:xO[�x������x1�`�y9Q�>����̚�<��O�͊�z�k�M/�¹�J;�
�>���+� 5�I���*�>�`O^F�-q��v����G�-�b�jAa����!�:g�R��]U����LAw��ތԺϯ=�hp1�WT�Q�e�L�lr�m�G�S�8��BG�h�O8-E�׽eϼ"��z7}n�u����gb�'�*����~�+��~~��'ë�[���^�Fٓ�]���:���{��B��K�w��Y��[��y��fh���>����d��:�{}����XA�F�W��M�{#�����~�v�����ݙ�1���}�Nk�ɟth�"}�kU8��x��f��8�߽�m�G`�R+��;k���WQc�%s�����)x���t+�=~��c�7�g�L���u�~ʱX���gG�9���q�w���L��Ng_�?�7���׷�8�z�B���t�^�����W�=���A{}�]y]��s'�T���)�+u2/Fn_I�����5V/Md���_�h�����V.����=4u�}t1�n>���ٞ��L�Mpq��i
Q,���."<b���ώ�:9*i���'�8��	���)U��9+KTN����5��dv;�N�ڹ��ܠEc���KX`LѓV[F�UiWV��i�m4��1�U-�Ǣ�14���C�w^&'��|��ܭ�ޣWLt��.S��l99�'��Xd8�@�ة4�������$�cr9~"#��rXv*���i� V�+�Y�Y����oZ�� �U7&Dm���g"�H&eTM��Y�wPKE�([�
F
t2!H�6����ԭl���i#�p�������N{�_���|�9����cؾ�k��c�*�j��;
�zj���+w����+�����M�L��dަ.��^��
�_e^h鄌S��~ܙ�*/�m�{�/�w���K��1N�Tmn��$I��3޼�
y�#=e�������`�so k�I^��:�qp�_,��>8��RwO��Ъ�+	Ƀ��g���	�vn�w����S^�IY-4��\?���3��%a�gW�r�y@2��>����Clg���%&y`>s���3o���)}(����q��(J���jy[DP>�1gw{�>�5�C�!u��E����I��%?��Uf]wtCooU���c7q�(�s��Е=Mc1$���V��O΁���k��$_�α
f�EF���F�󏬴~7�8�����W�c�c�\�����x�����P�c���=왂�S�vo��G�%Y#�W犗H1�	�*Q��*�I6)��_v��3�J��̭�}Ҽ޺���rp�G~�fA��gh�_�mM��
o��ٹ�G����w����F�7s-e[�>1�W?8��zZsh�A#0A�ZS����Xwq���J�f��x`�3z�f�w��ǷJ� T�����䓺��k*Z@���y	W�W��q���L=}��y�]�=�JRO��/�S�$�Ҳ��)�vi��@r:�6�9���4<��]��(e����~�y�M��v
���	nc��}[4+���YW�U�7�H�1�Ucz��`txǓ��=|@>�9�oOF��Cx��Ϻ>lX�>�=$8�MN�����]�kB)�݆�C�M(o��^o��_�:=z<;����wq��t���lȀR���8p)zq������&(���_�=_
� l=^�O�~����~d���}މYS~FJ�z�d��u������2���#F]F
�Dt�����pL�"�p��������Ŵ��{���4�!]5d;��彻�>k��]�­�wѮ��;�L^Kz��~�P�nd��,<t5"e�N�L��7t�U��K�n��Wr�KP*�!	m���i�Lz���u}'"_��Ԍ�-���y�:��=���P�G�к��O2���}�=�Wx|ڮ��������诇v����H�޾�+��T{�LG�mA$4BE��Ȼv�m�:�����b�F}�;2A�[4��{��(}�<��(����,�{KLE��U��;�E�gb'�ה�
iɍ����/�}��S`g�'�WΖ�T�V?g����y;�MR��^�!jӴ1�����m+���Y��ڬ/�%��b��>stݞ@�Z�����j�����V(�
�-�ƙF!�&�d�Eڒ��K�yg�n�R���;<�_U���N�}~��c�Z'� �5�t�95��}$72x�D�7�<��5X=a��T�b��C�GH�녜|�a�x�|�����o�}ګ�=�/�C�u旅�����K�9��=����F��Q�Yj�ר�������lZϒ����ꍳ��]^ȣs�~wg��� ��SM(_}��L /�b5�Dm����c�G��J�v�S)�]�M���,7��ǎm�w���1KP����G?���$a�"/���������J]VG4/�vQ���u�����o���(k�eT��뭨���揷[v�����4p釚���O��Mx���~<mV���a�p�邫��i��OR��;�X����<�j��_B�����/N��>�j�w�i�ߩ��@nκc��	�bGm`��Dv;��w2��v���5*��Nb�ۇ�[:s�T}�P"�A�=��f�|m�/�9���W�����tl;�EK�X�/��p�y������J~#�;)}Q�w3¸���I�O��������d���Vϼ�J#���F�n:.:7�� o�ٔR�|r瘩�T3]3~�[vʟ��c�5F�����z�z_��N�ЭJr�{��k-
�q>�}Ւ�)e�,��
dK�� [��nW0����")��{�����6���1ɚ�\�Xfʰ�l�Gv�jv;+)V�^O}���m��βЋmI���&2M @r
׿^�� K9l�CP
���z��8"v �����Mo<�Ǧ&�����u��X���WFY��jy5^���8��N6�;��>���^��1Nb웉9=�<��;�rP�we�c\trV�t��~�~�Oݩe>O�����zLW��5��Ż>��0�犵���q���|T��۔�]�\����Y� �Ok��z|�P���G��FpxH�J���7#�VY?(?kN��gzy�0hy����uW���d���ە�׬oť�\�}�����k�u97G�))��]}u�S�m:�Y_��n��G�|w��$��}�s�1/2B�˟eZ�s<<UK�q��E{���Q���%?��{���Ow�c��o�yoJ�J���S嚍�`.ӛ�#L	��e�<,��3f{{�w���1�����a��Us2<���!7��sg�f��T����{�=X�j6$B���-U6��ފ����[��;����gfEG1a
W\����|M/P1�?\)�5�=�͌���	u�����@ƹr�7N��X�"(ቷ�s�\���Q��ﱏ顊am�T���$�_g���2�3�B� ���JV90-�s��eݼ"n�yk�gc�r{K�M�ӌ�j�e�Iy �6,��H5���`'qܬQλ�Ԉ�HT=t�n �v��z��+�u��G&��f��=���r�q����c�U�u�YJ��v�u�̂�[ehd���6���-����ʀQ��d��]�/2��n�SQ�[��N7��	0�b�8��<��YA��af����H6�F���1	7�w����m�Z�%b��C!k^�_j�,1������\�j���ra����G��a���*���غ�����͆]�����z����A���=��~���}'��a�8c\үu-��#"=t	�pg�Z O�)v���ྻ+�|F����cL>�$�����s���3ٛ������8Wi�Y/.}��ϊ���`N-���!�}����ˑ?�ߺ���}����EW�`ɊB�ߢ:�՟�N~�Ms�xJ5���Ԏv3uH\�_�ݏWF�t��o��ϻ�~�7�w�/�U`�ϼ�:�݋��mѭ�K��q�=�(��}1E���0 �_]n��\�_���)�	���}ul���p{��(m*_�4<�O o�e?*i���v��5�"+Ɲ�V�t����X�����=w�U�l~��7F~��VIZ`28R	iJ�a���&�µd�7��dE_]]V��SK;4]l��*�:Vw�����J�!����h2�	{2�Y+����L�<@�də�?u�µ�}[JOt$�ݫ�)��D.�M�Fˏd觕�ENǌ��c�|��VkX�f˔��QA{�z��<��j�U��B��d٢9M�jXZ���ɱ����;�R�\����Z�.���J�ifӒɲk�|yZǲ�W2�	����rT�S6�s�`�+3toJ���/�a��-�E��n��Ϝk�I�~�TW
��m��0������B� \���랯��R�W�<X:�]b��TL\򉺛ښ��ėt�1��zk��T���~n��|82���;~l�'X~�gʅ��[�>���7R�c��&bO��� �ji�%ۿ4R�۷�赔����Lٶz}0�df�VϰFll�?�B�@����K�#���f��k��^燻��W@@Ϋc�D�<{r}=6���-��{^p+�+*~��l�>��viL��'��������]�x9�֟��15ҝ׳�n�_y*�5�y8�����vyL����Ѣ�a]ÕYbu[,�ت��9_�]�c㶏���'?E":�U���?O�V��Dd����RD�鄌�82鮸bn���ka�|� JWBk���=@Q����c��왣D|��7]�������+}�֮��}r^^Cu��>V�YUJ{�}.��w��G�kP9B_�o�ɫ�[>�Ma�=��Z�Wڮ�����]��/��3ٱ{jh��T��!�����B<v��]p��w�"��+&�jjߕH��7/����}��°XX�\)7PO��}N�],wG; �Ff��ѦF����v�-��-*���V�X�(nYn�K�y�6��L)�vj�;��!k&�⻉�	w�|�6Sޗ��!*d�a�όwo5W��qǌp���,��W����{�z'�gc϶��~%�c&�Fx�K��=j����ᕊ�޻�}�0�<2�����h���2;���%���Z���>��|���r`���*�<�T/s&c��`��t���J�^@."
�̜��yÄz~8�A�s)�,��g�P��$SN��� ��f��V�~�^��ʅ���W���L�j�E_g��*�hء�=oO[�lO
^?88D��<i��Hf�\4i6?����~HCL�����tLv;�����Q���u�����C2�dpǵ��x��=<��oM�ݷ�����}K	����Ѣ���&�7�n���V8}�﫸wc��vD�L?]5�UH����_{���ELI �$�V�����pI"�C�K�z��{q��O���Ɔ8���R���\5���R�0,ĩ���[��hϹo���6��L����k�|/c+�\���&�����I2��T<z~t����]*��زy�VU���ys4�*���� ��a��p|�+ۥ�S4^^&cԽuƈ?y��-)��dTyp��v���ze)~w��_�5���7T{�.{o�L�)���S(7ݏ��&�.�kf�Au��WmȄ����j�UU�W2&��7�7Ta͕ζ���G�o��m��0i�-j3�'v+�oI8~N���}w��)w{|�S��d{"I 䑗"g�q�C�S����f���F;�M	�7N�3�ȭ���_�����^\M8���7�\jVu:���W;�՗m���c��	�=W���`&��g.߳*�R�GZu���S��*"H>��c��8���;ck�o�.N]I^��t�g9��v;�PH��w���3�0j����6x�\�׫M�7>;q$�Z;��>9~1w�����E�8�9��c�*�:����M�~;�ϕ���w�@�b�T�K�{F��󜏥�4�Jǜ0kx0$�JAO'/-���=�dkNl0R�ފ����V�s�s��¯7�;����
8�>S������a�m�������"z�K'˳����Bx�����Ĺ}Hz�W����j�h&�oM��.'�&�ʠ�p�鱗Uq���>��=�K��&�ʀ�3��>{4���R�pF~�<�eeN8ݞ,�n�g���|u�zS �@o��{���@zp�;��4���`q+���':��O���k�[�fx�R��舍���y����y�av�O3�3�����/�NIގ'��g��^����ޫG)I��\�P�Lq ��)���\�)vŢ�/E������.Ď�N�d�2hBVu4%uםy�-'V���o4�5w��&CʊI�jF1�vm��r�eu��4�mͱ�5u9��>��<�,���ՏΓ|�X�R7a♋^�Y9՝���V���}�$��m���˨�7m�-����fS0���������ƺ��ĎSy�d�I�S��v4"g?h��(��͇W�ЭZ�1@�@ �p9�]�	޶� y�9k���0S�vS�NU:$U]�Ǩܣ��d&R%�*	��ݷJS��Ě:
�Pr��'�=[7{.������ �Ý��T�l̩�����ڧ�IdC4 .�n��*�l��O˶��L��`����8��q��99;q;�]�bsf�]�vAv���j�I�hoCBb
�Y�b�Z���v��o_^������$\_H�Kq+g�p�&����QSU�ƾڳ	�-�]�b1G],l:sgv\�!ՠu^q�;�Im���,���g�o]�Uz%5�i-�[��e䳀][h��*��ǎ�p�
��c�� ��\|��R�o/�U���u;N�QI�#�O��)��k�k����kPZ��b��=K�R���ZP�9)x�1���p�3���5�L��N�*���5u�*�{n���
�1@�w����*��.�9��4tsX�RN� 2F��2�n����oY��yI7@�
C&7�ss��n�d�ջ{j$�dT�2閕tP��u�ݳ�m���؆Zۖ�-������ˉ����ߙ%,ǧ�2^ ͶP�u$R����P�!ߥ�bư��E)�6<eV�c��6Z�5��]X����{���[2pUi��/F&'r*�%�TX�N���Z�����f�����N���]>܌���y��ZN,���{q�(;uk����e�+�����v,�jo@��d�$�,R���|,m�"��S�����4"ڬ�9$�m�7a[�B�2�*�vӽwυ&��=%�� ��;0	x��5��7O�SU��\m\`;�°� F��Jez�]]��d��w0#�3�Ui`~S7�%@)m�7)���]�U���jW�n��7�}nP��
 �O6K _k)�|��4�D��2�*�7S1Qj�u�L��O�*69G!�[`�V)�":���'�<����6��4ja�n�n�vה%*/�B�i��+a��H�@O���݇�U['c�o��c���*�&�d�HhM�{+z^U�h��m4,C���p4Z4�����I�+��u�d ݌���Rk�{+�����w���׆���|TPm��8@=i9p��S�oqX�PR�6��i����I�$��̒g��2(L�RT�rY�}��ub�A�㘬���d�Y�V%J�
�V�ܪ�OCX����OgS�,�ID��X"$
�]3bˍ.s2������8�dH-%	2-�Ei�D������m�k�̑�u��,��	����MA-XG}�^��G����WE�D�,�P Č ̋P�S��y�WZ�q����u���@ڑ85��[w
rZ!����Ue�ao���9�7V�T�s0P[lU1��uᎸ�Ax&��	Q��R�t�ED�a0_�8����)+$���Rej�6���G?w�P�H�LB��A��Z�i�ۭ&e���EwF��e1��_�-�E�)���F����M���,ff7m�0�"tԳ�vr����E�5�Z7�S;Vc��DL�ZG&����:�׃�����f%UE�T����L<�,��L���3N�6َ5�D�?d��<fEA؋�F�j�[�ڷ{�x&�kjߺ��)�V
����m�L���S)��	��3氏s����G;3��?�߮���gVF��n��d59������:��ެ��^��y֓Wz��ۢ*.~�L�叫L�f����]�5`5=�>糕$P�rxo��/�'��>���u&��]�����yPJ�Ѯ�9ԫ���v�^]�NH��5{�v�~����q0'	=t|������s�;��wg[�Af���1%/��F/SČ�w*�����o=]kٚ�Aw�t�2[Ƞ⻮�qX�p��L�eE}l{w���移�L:�S�/�|��31�X�n���s���c'T��,��#ϓ�&6MF�ղ�����;��9ʚ�v�5����<�]��7�v���7cg�WV�}���{�18�2��U��wW�j}m-HEn?h��P0Ӛ��eԖ���1�>Vje��N��?��[T������) +�4*��J傱�$J������!���o��%}�>� }G&�zW~��N��-䲾lܣ�织?(�^�39X<(��W���{V���h�S&��Ϥ�pu;�����f����s4�����mA�_� 9�K�����I�~�`�;&�7wԈ����h
}��\T:�l�k���#�ob8D�hKk{��t�MW���N	i�1n��Aω�wk^����ٸum�qᓱC�<m��:7h��"��sW{��#���}��<����A��/��ډ��k� 4Ֆ���ȱ������+�Ѱ�=�K3wk������ƺ�"d�"^G��=�tZK�3l�Q�#��z�^��Vj�=6�a	�^l���ni ��pYy_q�W}�R���x�?X���4���ҥP#*w�f��y�]�J�F\xVH�gd�|6:.�ǋ��G�d)<�E�z*���6[n��`�x��>w�x��}�6������X�=��Q1�է�:
���q�
���������Ot}t��+�510�?+�̼�1	���˗B����G'�s˭�A,Ա��Ɛ\s���]\���>��V&���G��b���DQQ�S�ϳm�r7q��*���򙊕���o�Ǯs8]�<7ؤ2���t5z`����V5u%�& +"�}2Y��^����)f���,]>����\��z�x}��fe�p~Q�L��\LZg6��y�&�����^����g�7#F�zO�u7]�,uz�]]��X{n��D�s������ M�]��a�W����A&o6fk]�1��;�δ�P5^�5���	���w�J�bJugto"�yB_	�����=k���w+�yMj���0�UT�a�/�C G,�&�of�P]�㥬f�;h��=`���BE��U&�v<��=6Mn�a�Jc�^N���[]�ʫ�5P�4����9~�d" �H�d�h�"�DG����y����}�:�厴�ohr�����p��YS����V�=�7�������G;s��=��"3p훭�����yn��`=�S����&���|�z�+� �N#�}�����j�T��z'm�O:��T���Vʇ���=�οB�ͩ^O~�����i�5�f���
ђ*�#I���@�O�B��~�esrŪM���K,h�>�S�'��p��sl|��^hĶ�f��{��fF�	�1sB��Wӝ8�=E+�{�{�e8y^��Dx��m֏��;	��������>˿&���o.\Ǖ���{GF�3K��݌�ڼ�C��SG�ժ=��E�4���#�ק�
X�ˮ���u�0�nz����� ��m7��z*�=��|$��mGT���	�����=�	������*;�����A+��{�����i��;������\�+:[�39ޤ��/CJ�D7>z�'����U���D:쯋�}R�����>O-����)S�O��QS����ݩ��ͫ������{u�2�������yK5�)�ʼ��
��=����:�)79��2����]�	��p���<�������(6�vn��u������5S]M<m��K�F�≞X����sg{U���B7�ON�~��;sڐ��U�y�����:l� �`���ۖ����?���/���{)����$��9�[|�]^�lYSQ�����-nn��Ř� ����yݚ����1U�R�|`Bv������
�K�R�ǧ&�l�У�:]���En[�8���$����2���`z��Yn�]��E�[��g��mp�ϤM���`������Y��o�ݣ߾HA�x�{B��R>�"|��z�;���v_{ئO��ݚ�k���bV1�|k�ܚ�5������^��?z+g��z���r*>��ۥn�{�}�>72lº�S+���>���/#q���T���Y�{���#hK^q��t��;�^���9se�t�)�8�?W��V�'=��8O��j8�!�"��$�!�^^��M;��p��@���0�%����׺�Gx�߯�투U�����|��;�^�F�L�۹x>P��S��n��I�]��^1~E�P"2$#[Dwbn�f�����\�^���<���s�x��I�����C����=u�e{=�q��\��Ks��e����9���R���*%��WW�}L�<�X�1���I�Ƽ �߽�-
���*�W5�T������u�7�{���W����r\����3�-̺p���o�ʰJo�P�{7�J���I`������KW��l-��v���qX�a.r�9go췡a-�2j� �U�()���Q~��ѧ������m��d�1��X��V8أ)Ŋf���r�\��WJ�VH�э��-����hߘ�B$�2a@�t2p��~N;�y����U����v�X��8$���g�D$�D�L(����u�}ׄ_j�=p��r�R�ŝ�>L<�V}��竷�r���隊�G!��)K��~3h|jV@P����Axj�ǐ8�{<��nq����"%1Q�UG��h�ԍWU�ل�=CƝ����j,�)^�N��� t���{��
UZ��o����}s��^��;����T��s�V���]z/��G'�Q�B`��b����Cݙ2�k������4�)�
�Og{I��:�CƘ�1k�][6O������fp�^�1�C�۝}Z�QԕS˾f����])]놝ڕ���"�?�)WYp4��Q�O�'��W�z�a�}<����5�9q)��&h3~���/� Y�r@�����gԻ��Ů�ȹ��oG�k�h	�$"��EꙏJ��M賞�(�[�)#���u�w�g^�MVE'3"*����8�F�u��A2@CB�Z���Ǉ��s������Y��9��ڮ�\�y3�����;Y~�ϵA����1����?<���ȍ���| y+�{>̯��w�B�|u�f`�=n�p��C�;X�V������U�Α%_�.�>�uԭ��l�:r���\V4m!�7��#�gp[��b=�V�����.��n�.sMҮn���v�gS;�����u.D�;+�w8�Zj1{���ɪ>CI�ݱ�Ƿ�r;"��]���W����|V���6��~ �o3�Y�=5���s3˂����ڸ�z�A�Ӫ�ڻ�{H�^�Z��v�ҁ{U�n<�c��JGqUt���p�dM���?1y��q���R��?\lh%�>'��8�Emb�l�ș=��x�#�?cwj��Iu�5+����=S�Vc�W`�����ra(|�E�Ϻ7���Շz����v٥�w��>��Kc�)�L� �Grk�;�C���-GLb�_[O#e�7��S�J�6�����p�8}�����u�S��̅���L�c�/5gF�J�sW��'�U+"VY[��#C���3s!+j��M�R�H	-�ۡ�����Z���>~7�u�^�^n<��?{A"�X/��0���x]�d ����o"+J�G�솏��	k��8��<\9I���9����#�@}'�+8�F�z�k/f:ɪǛ]�J�2=.��7P;Tz��̋����P�{����k]���8oʋ����T�~>w��T|M�=F����=Ӳc-;����2|�-�w���nMF:~�?��
0%�v���2�h�;�O�)�2J(_�����Zom�U�ז$0��6�J��=�b������)��8�mu�0lt{vՍ�hd �$�{�=��df�K+��g��|+Y�~b��57�v*c�5LN*�8}�����}|���Ξ��&A��{|��pgn��s.�sj{��Z�K0y�ꏅ��]rv7J	��sx�P��;��s�0s1��:�O��N�8����*��"����ýd�h]v��:��m�0��+s���oO���3yd�9>s������t̙���S#<v�g�"��pz'sˮ{�Ǎ!���}7�=��-o��T��g.o�t�-�-q8�#��Ԗg�%�qѷ�j���?|N������.6/0���L֔�����=k;��f��=��������c����=���v)��N蜈9�2����2��ns��崅T�c�$i��Y�þO9j_�(|W��R?�A����\�8z��=#+�I�8%�H~+��W�g7������O��Z|`���&c&`e��M��H������r��"eO#>p�սP����S���$��O�����q7qO�R�1�
}��cn8p&P�۱����0���c�2��٧���GU��k��3y����ވ��1'��+=g=.�b5�?r��'�+�D�˫��*naVm"B9W?�N�^�<����X":��;fq�-��_N�u����8F���e]c܊�� �a,�ַx`4�1-Q6�\u{�����[����4��}o�d���_C���
R|}ٽ>�V�	�;�Y$��A���_L]sh��xH��gxtE�����פ^yW�N���޴�g#�����<���]�E��-�3ِrC�{h��'Eb��BQ�r�V�;D�|�2´�N�D�-�.'I���1��	X6�+�u߱8���lom��י����r���c�Z�5���9YP�=�yrr(V���P@w��v�ȵ>{;�^}�e�/=&UJ��]�i<��&ƪ�ΨC{����/J�tXb���X��W���G_gc�S�Χ>��E*�+�&K3���1}�׶=�Ç^�3>02��9�\���Η�9���<٫~� ��~G����}�f/&�����F�t#+��ϓ���u;�����5�]���d������N�N��{4�:�kW�9^����;X�R����oy�B�����\�y{|�2�d�Z�T�&��m{0�]T��_-����3s�����H8��3�m��K�Ql��(����*w �fU*as�Y��3�݂��V��G�M@�8*�o-}�B'2j.=�=�~��3*(u8�b�>�a�h6�����j�W+}W��"����gJ��OW.��+�{�#�;���[�k�}��x(���}��S�գ��gQ��5��2�!D��j������s���E�9�9��y���x213B�m��d��x,^+�u�&�ט}�,�rEk!��&YcS�q�/�a4�K]Ʊ�؛n	2�[F7i�eCqϽd�=��Z����+jɿ6 �J��x7=s�<��U�X�-%
�e�������bR�El\�9�� �~7���k�}Yƭ�>�=��/1�����ۊ��"�c�욤	j{�{ս�����;8�`�e>����͖	P7ti��LlTV )�v_��t%��9D��pcݰ=#Q��w�ۍU�����1�Gɤ�B8t���-W�[U��u�&c�8o� T�E�|d��x�}$Ϯ<ܣ�-����ʇ����,{i}�Q!Ξ���]m����/s��}����>Ʀ��A��S��b�ܱ��G���\��2}0i����d�����&���s'q�b�uȺ�)g��'=q�%�|��g9�y����G��y��lXAM1&���ڢ�f��ȸ�����5��y�@� �R3�����);��s��2|Y14�=�X�A�D���k��ޢ��[��a�^vN����W�=��2!���r�$��qwΡ�*��c�Ò7b�[Q'�I�G`�h	�I�TSY%B�G��t����ݯ	��UO$j��מ��^���+�3�9��]Nn���1�:���wO7��0n��Z졪3�v?4>L��������췏0������-��9y�{�*����aŷqН}Cm��C�8�b��a�y���U�%Zʷu�R;���o;�ԩf8�z2�㻹��j��o?M�Gk���S�l]r���6�c.L�ampi��ÏoW19]����>n�Oa{��}~��U��s{�'r}���;gb����� �}H�`����O�Eį0X��)H���hz�X�˪����X��)\���F5�ܐ'���DF�/T*~�*'��V(%B&c
�1љv���rL�vW�:��.��>��
jf��;��I�'܂t�jw����&�݇	tP��ɵ^ʉ�Do��b���UaOoo������?n��y�3I3&E��:s�>��ʔi��/���^�$d�p��:�{;d�ɕ�^ep>���@,�A�uq��]�ď�v�9��]�-��af��eX�i�I\˺ Q @�!I� A>�'� 6���u�S	�~ܪ������{�M������[��TX�/����=�9J����C��e�Si��Gd	�Tt�њ9�n��0y��o��~p�N���L	ltEx��efn�j"V����Ӊa���ޣN�D����{��k�g6+�������n�0�/՛�BqP�,��5�s�h�aCÐ�6뽟lH��G[�C�t�K��o챕3��WjK����PVV�݊�'t]�5���&�bʘ/&���,p����P�r��2 {��-��T�r������ܓ�{i�|�^tÕ�iky��=M�^�}��P�ld3�Ⱥ����;�7��d�Tɒ�:�z�t���/�Cg�Q���а4Q���\�]+S:�|�p�gIF�����V��1�	.2I.�Vn�'�BC'����]��%����[LH��#y�p�S;�Y�5����[Mݮ��v�v�t-��� �+v���=j3x�to�w�^�kb�na���X������Xr����S�^_C�4�#}O��nS JQ�Q���މ$�7���D�:��S����\z�Z2�R�q��d�����rU/�9[j]"Ż�ݚ�jo%�(�Cj0$���l�c�;�6�� �I"wa��8�с���f�Kmp�����,�8-~vȱu_EN�� o͇m��V�oQ��௩mΎvV�����Y�i���b���c}��Ҥ/�m���V�۸�O�1_�nѐ7(�w���;�J�5ν�nM�I�Q���V��V�9?�����e<�B��5v��ŶH��귁+}w�|)��ҏ93���xh��]��%���x8r�kC"�
���wEo�{7h��XP����L.|�3��pd��M�tX7ηJ��Y}L.ʐ���d䊠��K�}�}Hܚw�1�$7�����o�}#�N�f��V]��Q5&����7�������o
��]_M�ūغ��]�'y��c�Y��oVp�6}�ibldYY���ۚ2��r%��ǮK��j�'dӟ����O��&���n�vR
��{W��Zna�?sֶ���KZ�����
�x��V,hX�����Fa�ⱷD�R�cjڄQ�r�����\Ix�2��u���9��53���4cGh���VA�f��� �ƥ�˕�B�&���90���q�C��(`	Yޥ�݆��W��j�?u�������h�|�$䫆,��2G���4ƼG��aOf�.���7]tؔr	o��tKb��3�jm�롋)k�\��]j�r�vqɼE��(ۋ''�:;'i���ж6�,��|#��Ͼ�x�#��W9�y��1���&$g������@��B��w�B��G�y䐮+�=j�����}�;�.�����nE}쾹��a��Q>�Z9G�O۾���O:&
)MV޽�)ÊW�n%N�ӏAo��]&hg\����r��>�RW0:Ǜ\=��gW�����̿��$^�'�r�)-�C�_}�ٹ��5��ξ�?u�ޙ+���P6{��o_]��K���Q��S�͘(ZGg�7km�b������$����l���"ff��R��������^}{�}yn�^M%�U�j�no���O��5�1w�^�T/�_�g��YVր8�������=-��ϯ��{1N��'�ؗ�&�*�~�ێ��玀7.'E���b�j���F��ϥD{��f��qx]���2d��;��^m�rS��2Ϋ���騧�J�����1���wS�wOU}�$�X��AlZ����Tk�u��Gݔ;;gh�oVne�K��{���CZ/��U��m��@�+�u������U�(�/dױ^w���9%���ʢ|K�� �ugth��z�[*�8Ĕ� ��^���`��4Onq4��c�a�[ ޝ�WG���6����x˷sUXNpy�*���v�Y��b��؛B�z�4@��:㱛�ϩ�^4�|�!���1y���>]=l�c���/�=�֍�s����w�Й��B�ڞ[^�����z��2ǿ?���kk��U@��^r�MX&�vS�����s? $�gr�S��!�jEen�g��z�72*!"�4�Vn����n�E�O��y�����1���v�i	P�0�pY��ͽ���{�OMl3쭂���x!�<�l��/F��}���8*k�+s�����^L��%0���r���R�㸩�w=�;���q(
�&���s�Y1�*V�8�Վ\��뉓�o3)7	dգJY�>�����F-�:��O]G,���:�����U�t��b��hc��I�V���H��B��W^����n�j�z{���Í�~��"�J�+v~���%K��쭥N�P�ʿ����g��F���챾��E�z�d�x��ixfH���+�h�Ut�J�T6jR�7��}�{�+�@PH��4~��}��Zp���Ϩ��TU݂��Y3o0�o�h5n�ꌪ *˙~��;�P�󝛧��+�EAɕ�f��MpejކME�Rv����`�jq��X�:�T��+�p��-�W�p�
gM�
9x��uz��0�D��e�&� K`�gSz;�7����@��dS	�	I�j2[YU p�-[u�ۡ�ؚ��wH�,�uUs*$M�n|H�(*&.ffa��d3B�(�U�N�[z�AxS���`�x��\{�o�X�q5��R��"4�cQ�4�4��a>@�aH��_�<�
�Bzi$���4 e����N��}7��h_z��
�5�eSǦw�
on��Z����Ǿ�g5���U�7^`S��ơ�7j��*��0{� J���"G�x>yң#��Uэ0���@�}t��x�"��������\&5i#ס�=�¶�b]]�o<ɝ)O�פ�TCN*g,{-����bm�{d��λ-6�G�e�S�fp�gc>ɨ�㋷)� Bxm�h�z,�q訣�Oٙ���ʵW��K��"h�����o�[ ޥ��g�{��K.�^�P3����v-���W^xRT����{�M»�t6te߯�Us��uOY�����U5B���0 T��R��Ƌ�*�����|q��u����G���y�5Y�W`����t$��s��U+E��"�ߤO���U���a�xN��$6&S@�nW��k�8WƓ����B7kk�:�]��������� Ul�����T�a�B)�9wՑ*2	n���l��ڷ�a�5;'�¥�Y٤����R�c�^��2K��Oy���w�WH��}��ufnw���:E��v���/�`��?Ӧ���W���˭�F��U{���1(^ͧZqgVV
�o��u��X�F��E��q�,��:z����.��+��¸qѹw�R��&���I���[Z����%[����!)��|�g��=;~7����goO��'��<�=}�W���W|���)�2��E����&�ZDz"N%�.�/v)Ы{�}~}�n�eZ𫹪�eD�)W��v9y�/m�~���I&6�*��=�jۭ"x*/�F쿢z�ÿ/�����v�b�w���)��DG+>M	�ڄh�ZOy�f�'��fϻ�RC����)W��v���;@�ys��g눗�d�SwB�<�Q쒷|n����,�
7�p�j�̫�������&��ן1�˹�����y��&�����رH�jA�[��O���X�R4)��$&:wH�+0�?~��ml����/,������t_w̻�u�3N<J57ʳԺ���'s�=]�W-��};^؛Uy���T�g��{J����vp-!M���e�4|��{��y��5/w�T���*�W {;=����	�쪦E}3��[#��5y�_>x��r8��}���:+xO�MU����Qu��#���f�u�@��p��
��$���ws(��6��Y\�Պ1!b�Q"L���	y�{vch�Wz%��^;���u�p��E���H&�x�lwX7�UZig�n��Żhdq��Co��ɷ}�MwjT&� ����ͼL��W��=��:�lj�SO�9�������0%zO.���w�gq�^OR�t��O}���x:���gz3ƌ5�7)��Y����ؽ�&z��c��6�.+�ǹ�*���o�O���x�-��VE������;��Z���{�v���Ty�������������F��|"X:.-d�h�ӏ��VZ�{Q��v,�p��UZ=��6OJE�?���{��a%N�<����'Z�=px�u_�?�&��{[Qۉ9���G�V�l�O���D�ˀ���~}mO����"*9ݯ�����}V@�Fo]��YpW�ʬ��WVeJ{{��+�)�W��{\�s�y4bk+3��ң�j�8&{%���R����{���Y��~�]N"T�[~�mZ\��n����{Lyݠ�2c9�{VN@ځu[���,����G��*t��>)AW�S�/�y9�͸��dׄ�m�z�y��yf���t}��k����X���V8�/�=�9�gVU��Zh�������e��]�g8U�j([�P?�W�<�e�_�\V��u��]	u�Y�����:�1�jSS�����Ⲋ��E��ν2v6�F�kM�wr�����I]6�F\N���n��cw=�)��+[�0m2���m��<�:B���̡���*�ݯ�j�o�v�c��)Ǖ�y_U?LMw��4GQ;�e�=���WN��w|g��#�$��4.o�77�פZ��W��nv^^���ҡ���}�K����y���������?bB�S����e;_�7�e�\!-e(�ePad$���$k�}��8	ϔ�GS�v��z�RJobS��
����ّ����ws��x|��E͕y��җ�N�����~^��.={�c�(�n}�����tz�_g��s���iv���I9��uu����B�8;�D
7y�R����_ض��}�"#�<�1���l�]������c<��ɔ2f���N28O?v�>���֘�=6�LQM��w�1�|Yݽ��g��TC~�������_|;�zxeT[ƞ���1���U눪�����s�˺�����+�v�k��e_��w���~�0���~��d;ȳV��fmR�?6��>��`科��w��xԿ���q�'M�a���g��w`&*��h��9Vo:��M��W�o�ْ<����ic�Ǉ}��T->���O�o@���)=>��K�7;E��y}2����M��y��H��TZl�ُdR�C��µ�\����o����u��fS�V�V��D�C��c0aG���]���k���*�vLE]��GZ��V�Alh]�5�t�g�qg�ݭ��j����-�
2ۭw���FӴ�Z0�;.�?."�fL�:hu��(�@@��Q�\�L�LmN�O��u���kmR�e�j�P@<2���,�S�&�X���B�d�u�,ݚ&:�(28�����-.2��YI�X7����HE��Ql6��8?����>2��l�HU�JlS;��w�}���;��Ǆ\�#W(7@;���o�(f�22���磐Y�ވ�0D�q�)s��r����VwO�[*�_�Flu�2�����1���ۭRn�Ю �Dߺ�Y��^��]+K^bߏ�u�n�^����<�ND۵2=�����fg��F{�]������5�g�+�K:���q�~��b�_y䝔�&�N?��K�bF���ܖ�j���4�@�{ڽaEϗ>.-��FG*�˄�qj^r�Cr�{2}xEXڌ�x�idl
_k�~wf��"c�'�f�Z����IܩH������ܭW^���y�潖}���8����@%�K��ʥ=;4n�3�ʬ�68)�n ���ئmb���:���5g�+��J*X�����-�(�7-�h���/Mz�����Wl���3���F���3���A������NjN8�q����L���Ki/f�����xoS�c߹\���#\�O����g�4��Hd:����}�U���q/<�M2�є�����j�r�Qɤ>2�owo��g<�������Wn=���kyc��Vu��hT=h��8�9u9u���,VN�i�㹋->;{��2MR�q�O�\�.�,9�@}G�z�qt�q�x�R������*�S�8���?w{y1F���W7�=T`��$�����Rj������N}�N��.�k����� �ȈhJ���	U���p	ӷXg�U�c����<�xAW���&vws�f����k6���y�D��Z��}����Sc<�<��ڗ5M�L�t"}n�}#vvY�0*7�3�l�IQ�N��|��I��3'}Gr�V)s��%��vO����ܨ)�ޡ~��n�oz���9�u�r���"�/���ޮzc�t��˔�2��m$�qx��]�/%�&Uk�;]��7Pi��\����D�h�~_���R�u���N�����ӏ$�_Nl����.֒���<vRv����7�rR��6 �{v�onED']�TzD��oω�OΞFn�Q~�cG7r�۞:2T_|v}k�ϕ)h��s�	�Ә9��^�[�s����L��1mIU��-پ;ٮ;��ѹ["�k�J1v�(;�y����o]m�S�#�Z��ؓ�v|��OH�!9W�f���:�	C9U����fn1��*�<�I��ǂ�ABؽ��]]�dx�r3;�ock��`�ۏ7�u��.��\��g�4���u�X��wD=7����~N�3�ЎVcu{Ls3�����|\�g�+�ĩ����p��	h�Ry�c�)���9�z�蘼(ϡ�c�d���-T��ԟ*yS�s�('����Cw�z�=Y9����ҥ�>8��1�%@���q�`�ydD�zȐ��;�{�SϽv;�w�w0D���0w�w��W�(�M �9�gE�G����eኆQ���~i3��X� ���:�h2+ŭM�����I��竞���Y��VOc��p��u�c�qj8ϿG�q�������feu����mDRe��dN�ݵ�s#uAU�;�%{<F��g��<b�J�s�]�+�6q]�~yy_ooxb{�WԇP�4��^��]E|�V\lm���/@�������������e��j��x.g�I ��V�CÏ֓afio;�(��f�� T�L���s�e����J63s���O)��w�gD��a"3��6�%z��ڧ��%�t�W�D=��=��n��O}��(�W��A�fwn)g��zO��ु�X[�����a__t�:��F0���ƷV�z���ZO�p���P4se2���m���d,���wm�L�_@m��K�S��Gl�=w��M)�h��uC�T]���]�;���Y��a�֔i��g��^��Ϲ�ؽKµ�X���-k[Am����fn[�z���V���(�>��&&���J����վ��t}�?bh��
�ǟ�;2�2I[��>EMBWd��_�M�#&<Yu�ͽޣٵ����-�4X�7W���4��tY^㤿���Ϟ�������̼�k#~�ȗ2���%R���$�:���gY�D��G�K���#�r�6��%�N���~/'�{m�:�ǵ{�~���"�R�m�^G�Zztu۱9w���*n�ڥ�"L2�#ʅ�;�q�u[��2Cm��Od�ӸLg[S6�cWj�-�2ϔ�M�7�{}S Q�>��3�N>~�,h9��̒$�7��d=F��{Djp��Y�9��ggC�5wU��l�t>�'FG��d^���X�ǳ�Tns�(]ٞ�{�p�Ɉ���'��.׫�4n؉����w"bz$�i���^�c�����ۢ�7;�{/[�%� �������t�����&Vg���Va�쪣$yu]G�#�1��y��������H4��S�B;���ͦ�:^��&.![���q����+t�\	~Keqr��\�e>��wF���	9z���D�C4��=I�MGH�\�Y'��׹�\��ڮ���1���h������z
����0𱻹uDŀH�*����P�n���Ñ�E.�����f�q-�IM�5��is�-i���� �o	iZ��4�:���c =	Ϳ,�8�@�"�!�5��\ɓGi#��XÂ���3ZUkN��u��+�4�˪�`v:�@��ps�λo��7��lN�Y���<�����Ei��b�1��`>p�����IntBB4���.�{��_I��甙�0���4��A8GF��:{%It��r��l���j�4����W;7�[74�oB�+�!�V��U�g�w xY����x�"�m�'qw���k�� 9.�x:I�8�I�kw%f[���M���rƓ3ssQ〫3�69��!@��4Kח +3���mv�����={q�]4�ͧ����]o5I� ��8�梧$� f]xL�ټ��5��/��1U���y׀�"26��K*��,`�L�{�24�sJ��_�Ocq�t��
}u�*�N��]���Zb)\9pf�#,�&�f��th5zZs{N�[b�D��[1N�а:�rWPу3+�p���l���p�Kɹ6u��g��-�/�:ɂ~���P]����Gt�ꛋ
�j�N̮�+�"�`;;tH_�\�ҩ�oc����}#�b� ����ec��$�9,�-Lp���ݐ�I+N[{l.9am��KrnW[��:��pj��3�'d�ZTdR�ٜ����<nR�����>2E�Y�qQ��c��%&���	����r�WU�+��i�HJL]X�nd���!v�����S5caYRT��}�;u���JYׂ�3J�]����YK���+�\�'����ZpJ�,�WU	a���	V����&�"�ǵ�u��!��[�yR� h�WoF,=�jvw-Wv��(�u�
�Zj�!�'��/��gJ�w$
�̺��4�r��i�\��h9!�6�XTK���v���FN�Sv,���],��`��^ȁ�?������B`/]��BsEJ3�`P�Dk�����.]�b�Т����Y�p��A�i�E5J�Q���ߞ
��,EY�%O-�m�u�e�I��~ES���Qi�7+�ڷQ����&�-�ƍ|��8��98z��8���,�����?r�Ȧ4��mƋ�ZԦx� ����C��l*�(U�B��8���2�M��H'�"!�����+��	�)-�"��t����6�U�sswP�\sӹ�����L����U<
��Ӊ�UAf(礌�p�ے`���7�Sp*���)o*�^3Ad%��D)�7QN���֌���L�pM��'6H�f}J�X��I���L��ʍ��k��%i�4���2�3���I4��rC�f�"�Uu�'�&��@��^ҩ�ݜ���KO�rcF�X�e
Z��L�>�Q��([=gmcaСs�HeP�s]��B�m���2�k�l�ǐ����60�p��;��mlȡ��&�ͺ(�oEύnY�?�W��1Y�p��
댎���;4a����Ak]݂��y���7#g�)���k������ݩL����J�9���P?ݔN����j�r��������z �e��6XQ �,�����՛�\�ņ�4Q�Vv+�q�}/�k����ÉxIݑ�cb:��謰U��1�$n�*�O`���`eZ˅���7�c�8�V�9�SvQ8Z'Z�B���wI|�`��BJr",�#�RZ��O�O�C6��7"�a�w���K�E5Pd@�bd%�r��\��]*��!,�i�ɟ\���^R���VN��7�]_*Ni�͜*��g{F}2}�Gl��ܳ=�y�����S\(C-I�O2v&���&�|E��I[\7W��lYq7�@�ď�R/�>���]9>^����r2β��T^̩{gp6��{��s�����ߏiN�\�l��	�9���Yd����s���f3X�ǒg'�op7P��j!Z/�x�� �]}@��]�dT74+q��͌8,V�:|��dI�1ѫ���1kxN,ܹuq�ۻN�=쨞ׯ��j�t���IX������u�����>Y�kl;��xsmu�e��\�|�<�e+U�4fX���׻%�qݱ���N�Q���6�S�&���r��Ϯ{�%U���BƬ�_^ע~L0/�.���`�{= ��|�e��Ylapɓ�,t���2��
�Q�h�M�|��[e�8����ρc�N-��#/�ЏNF��vr�X}ԟ�r�3N�����d^��-�J�	�Œ�	�{�;���(�k�y"�.���T�\'9h�����zT�n�+��*�s�
�w\,�}pLl��	S��z:��N2�P��C��ݥش��⭴8ifc��ϝ��`��f�	'��;rŮ&�_I&������u�y>�1�w��y�1�Zn���牣gh��Ʉ�:�>~�A�?[�E��ʔT����}G����5(6>�Jk��~s4�����-z
�z����]b=Į�CWt��H����K��N a�/3��+�w�=ګ�9��y��N5��S��GZ|�hwT�Qs�}Z:��z���%����4��%Vx�1�c:Ϧ�G���}۹���<�v0��6�ǯ��w��V�
�3>١���]I�h�}����#�֓�P6^�ϟ�¢��ͼ�,�)��Gю�jW�>]"���\�>CY����N�(��zU�ʡ!�cs�V���1��YE �I�#O[��@�Sa��~���?�+�ʚ��#У�y���X}'f�o+��c�F�v�ӗc�F�h��.�� �۬Hw�6��[H[0|"v��x��ٮ��UW#8�`����j|r�2�cR�%�~�y)V>���Vߩxg�z5j6�L��J�������n��p�Z����0���w����y4�W�q��u<�sSw�VZ�]u	~��ŧ�˖韯��E����e��eId����yˆ��z0�t��M�����(=:g]@���P�� Q����4�6gZ�k)4s{$b�����_v�9���e>�a8T�}OT�ӝ��6o�r
Ϙ8b8�u2�x�K�!1��o����*3�޽@����.ݮ:��ۻ�鋁T�T��o�\;4�hE�^���*3d��TC�'{�f�."wn7���D��yL�$��s�wו�\]������B�O>�c����8��͜_r�|$�aSۼy��1V�YK�9���v�;�]C�HS}k�ي5�YF::��I������#�f	i�s�l��:*�g!{k�&�@v�"�I��������\1E�)Ș@�O�b/Y�b���-��5^
���O\W}�� �)9���*d知����v�� �<nM�w�� 2���u,��q�^N�۳�S��}�Y����l������ �E�U>�8Ш�|�Ď��7�5U�����&$F���[�,w����e6NEz�|q��s�}Y�no/{i��ޭ�p�J>[^�%ߖoV�!�Ă�N3���ڏu�4a����͉s���z�S��%	�*g�q��Y�_�*�F����?X�*.�}����+l������s&Cg:��ڛ|B
�^).��i��Nm�5֦k	@�٦�n�%	�����l�9��GX����	�/q�]� �2���%�O;[;/�'v>�^4c�j���=�>˴V6e!���u�e_��{s�ƺ��8zϨD4�Q��*���9hgo��WG��Z�{.�dFv��W��˱� ������ˮ[^(1����dʟ��.�ڸ���D6�
��:���ъ�	���|(ݻW���fE�qx��ɔi�wzC�~��S���F�ϼ�q��yf�՗��}��&=a�V(�Lۡe��o���掿.��;/JY.-��D�����λWs��K�|��y����
{v�Ђ��ys��LȽO���^���.��7�W����^�\]��G�I�r�z�swg'Q�oN��wr���<�
���Wȹ�Fj���z<�"��]8�ei�Q|�c����Ҽ�g���s�&wL=�Z��Z��n��ГU�L���Xz�`S�Uc���b���������Y{o6%�zZ����E�³kwM?i�o���EF]��b��R���3^z�EO�A��n��f�����#���'�Iu����'s&��״����e�^��� E/,=����=n��C<m�[��B�[�!|�*c�:W��9����X�*`Ep��2�0��m�EV�"0���Ʒr�:b.���(ا��C�0*�,��*gsv=��f�tu�K3�e`�թ�8�H2�[��^g��w)�1d	(��u�?u�2(�L�8	U��P[@&+�Վ	G-��!�q�_��K-G�ٱU�m���E_L#�g��Ε� ����N�=J�uKfc��[Z��j���$����4K�8�ۋ!K�s�;6�4b�Be���km@@���Fb�t ϾS��癈�1.������Υ��k�T�]�.�gS�ݮF����������/|�
�q��B��VN�n�7ʟ��3��f�ݺ��k�w����^Ǐ�����s1ݽ�3���s�eeo���hzـ-6���o��]z>�r<��Wbo��^�l���!�2)��
���5���# ����W���E_�::=��5A9�q�j]����.7���ّp������,������_o�v�j��1D�<�;�����6*q�E_�;�������BV�����x�/W�g��]>r�{2��PC�vNN��#*`�ϕ]VGE���=��Rf���������Z��Y�_� �z�\�m^T���9dP�s::(�y�(��y����T�)U�Q6RF���i����`dn({%,2U%�����T����Qj��x�f�"&��B�?,��O�R�Q��w	���Ӛ�Y����yyu���{��x(cM�������װK�	�tn�|�Rؾ�V"\���o)�u����m��(�R�Shl&2��N�J�k+���<���h���q���: K����0�kD�2�\zA,��}*����3�C�Q�s�$Q��;�j�ML]�zr�u�ˇ?Q����Vh}��.��e�B���,�~����΄֡�߷@��f�缯uMo^�Rٌ݃k��O?�����W���}�x��M�9�Y�ً�x�������g��� �!5�ޤv*Ca}�~���\�2#<��s������q�?���^�]ܾ���]���J���n�H{�Uq�rTk~�$Y2	""���y���c_��^�*������}�9���������ِ¾��K�78�^��K27�f�?��ߡ�ѺϽ�ͳ����:]FƢkM�q�'r�+����ܫ�N>�ڢ ��l'��unJE|�_�r'#��u�K��?udϵ��ͱ�m"�*�{9��
�_Q�q�o.x5������%F�=����d�F\��
�я;��:����ͬ���]o �u�Ӌ[��Q��
�q�}���(.��<��s����qZF]�nv1VӷM\�&u�Ҍ�+�]^c���MQ��j����5����o��dP.�X?l�;R4p�+��v�]ȸ,�-����-j̳���_�.�N�p��Ha��9�2��Yp^�5�{[r>�d�u��X3V�d�;y��յ��u͡v� ������R�zk�de����%��c�&�y}���{$ɝ�����j�7�>�V�ٛ�s��D����϶�[���xg���s+�Z4(Vd9٫}o"�C������>������'�WŤ�B�˗\˨�;�6�:�ע��-�bE��л9c[Rr}�}�R�+�|�x{�c�oC��u�����M�ײ�~@Ƥ�N�σߕ[P<��_�������	~��
G[
�QX
����竦��׏H�.x�I�Q8�8�u�w���ڑ8���.��	Ofn���S�o�vj����B�w��~������9c���<�O�b����z?v�Z�ߤ��W��5���.��e^��i�v:7�p���h��Y�PC�o˦m���]�t��������3q��g�k�I������z����kAE/��٥nj��_f�7)�ׯ%+.N��b�ɕ��<cԧP�� �6��K�q5Zs:��7QU��,���M�oOb�]�O����.����\On�/������N���^�Xb�|�L��0�g8�Գ��
;ݻDd�#�
P�j͗���9^ЮhaVH��C�ndT��Y��NpY�tG�烚�M�vZ�+V��m�Vd��V]��}9�zwT��`^D:�+=(�:)4Ѷ���e����L`ɳ����;|��oE��n����{�7�$�d/T��]��j#{�����6�D�=�+��	͈1Q�sk/"ɳ��d��5m�)%r���U���-4t���u�z�Y��ԫQ�h�d�*�];k_���~���O�Q��٩��zVU�W������=�dVy����^͆=��'~D�oq=��7�_�J��5ME�V=�~2���=�C��[��넳�-?c�ذ�ׅw���]��.m,�sww�~*}�<g���#�?B���3F�z�͆X��ф!�Z�֨M�f�r���r�>�u����bJ=~����W�Ѹ�ǢQ�q�=�O�V�2�M��n����Uv�XF~�EL�w���;a��䳜��9�Xڊ��@B�����[r����$��o���J�Ww���GNue���W����5�C�b�׽�`�9�y�G/2���m�֨>�H�q���j��ٸƝ�1��C�I�ȸ3�;^�T@��]�BgA�UO�^�o
�..�nF]�����9��3��WY���o?d�����7�T�[-<��$N��fy}��	�ߵ�[��%��G;{��o*A�������YH��a>+��� d�IJ�.Ef�h��q�\m���Q�r���u�8"WY ~
4e��,�L2(ӏ:�Z��Η]{�����!��9+j7�m�*��^fZ�T�&t�G�U�X4���^�Dg��Տ)�G\��Uj�d�ȁ"��I�U8�ز"�f˥�ܣ!�!7M��ƣ
:f����}"DA$x[~q�v��4}	� �ya�O��~���Wøt����=�ߕC0X��xǬM��ܧ�f��e�V����/c��>���8�Ҭz�Ecs��U�ab����c�����~�Vc&���o>�;\^��=Us���$�5
}�q�h�M�V���@�vdfeh�}�l�S��0C8�R�ߧLi�Q��2�]�ޟ
ș�mSriGy��z\q��Gl�܌J��W�A���;��*O���`�����m;u��^O���e�J���K�	B�Uؠ�q�h[S�{���/	%]�y%�}���o��2v�f���R:G��}����i�|ji��g*�^����rTRr����4\���J|{~N�]{5��f=I*=���b���
g$@@�%�k�lRA�lLj���\n�)��[N��O"��=:��_L1����Z8��p�6>�_c�Bv̂d1>�2o��A�6��/�L���i=n���htC�m��������6���+H�Kߟ��7y>սw���-4d����n�G���n�4��;R��E�4\O�gn��D�|/n��!x��f�%vي8�����KNXƎ��k�y
�k�Qimi��l�42�7��IJ3�Ǫg3-�^��5mh��K�}9ў�t�	�yq�]�~�������k��e;�cnrU�bȭ�R.�INS�5N�*|W�}u�[i��{6WC�r��wR�Z/��S��_�7��כ�شPD	�ҟx���V+ik��׵$�C��@}�k-g�x�=4f�6��^e�8�>��hۮԮ��Z�h��z�t���Q�_�H��&��z� Ƿ�p������}<�����{���P?�J����*�Ṿ����Q���v�|}�ۭ�������"��#�(���[���u����v���ݝ��}���z�I�m�Pw��f[#�>"o�j5���w�ʝS[�S�.�;�<qd��ˍ�p̸��}�Y�rb�6�� ޿HG�O�/��yt{{�[љé��Uo����W����0A� ��~sHy�f���:��>���+��޳*&�����o���rY������+Z�c־,{��t>��Lg�εz]=��j�_T@&j���OFv����^ͭ�u�l�#�Y�ҝq���{?yeAl��.�V*����lA�R�a�Ξ7Ү�᫑�	�)uf>�{������{��F6hZy ��e��=��i8/���'���\A|��+����钙,��q�F�M�LB��+j�t��V.ea����0�Q�[۹��]�n⁚m��H�u~����ï!��7��n��\c��Pý����]�!�lS��L�&�X+�t���&�^��(S�6���1��0�.A���d��{sN���(�K�:\�����l�<�O�!3oY�P�l���'�5f_b�\1<��h7��t��[N���-����c��kkm�e_b眺s�I��B�w�r��������&/��]�h+�����{8W&��uϦCC)��V$I��C;�zE��7kܼ�>s�r[9� ��鹄T�3�a�Y{��bݴ�W�fdxW��:���9ݠ]1 n���Gg��;��2R�A�Vs�g�@,6��uŦ�BᙻA�ooy�S�������/�i1����I_�q��d�8�ծ�j׃�=�d�S���Vrʗ^�T(�nVG���֗��B�����X�1�(�%��*�"2`�b)5�ۦ�>�ٗ֌�E��hPqP����+x`�68�\�����$�7i<��S�+s��@և��/�%I���yp�־庈Vc�/��3-e���Vs�q<%e5e������n��'-����uS[��ޓ�~1�©�+�u�eo6�W]��� F�"S)��u����g���2�q%�m\m��N�F��6�F�Ӝ�"Jk�<��e�8��9=���J�bQ��%Z�{�)�W�-�#��J"V�ŏ���Z{lo��:E)i�1@o��X���J�� ŊL�󑑖�9F����:�
�7�d����i�W�r�����g.<
sdm�;[!w�6�m�3,a��t7{_sz2�LK+��k�I�t�U�j� �R��mǱ�8/t�r܀����U.��W��s�Ɠ�Mf����h�R��U���]���bخc�2��v�鮙��]׊�}0���w8�g2��oC-�p���Xt�f�3PF��)�.V�;��v�ET������[i@��G�v~軈�o�)y�S����1�� b���9E�,��u�]�B��;EC�yka��r�NX��깱kn������{Ǻ����~���uZ6x`~&$�Պ��<��ϣX<s�ͥ������b۝R�2�'�i�#`˿!�� I�5U�"�p�\y��>��k2fu��T�T�9��'��$��I���3\�1ˆ�Vc��w��f�E�x��
�ח��7��֬�v��ɳ}�lMS��NJ�����ԫG���	f,�[�0-�rة�[jm���(ԯ��)p:K��9m����Nڨ�Y��}4i���z"T���#��DZ{ے�efm�%��1�;��K�[��>���mM�eL�|���ŋ;�EYW�6��p�w�β�w�穼��]��{�p�N��*tx�*&jz�޺y���9�w��ʹbmY�o6����O��ǣ}0A�8{W[ޫ��n�|�]��dOzJ۞���T{�}����$^���LW'���\�Sо�����F� LC7��P}�y12�o�D�F=�ͷ��v�����f,/{�|�b�<�u�=��<�|tg2Y�FO��S��d���e��6kpC��4�IH��.����<����=;j�zÝu܁#����2�V[*�G.�d�/�0+�KN��ۡ��:F��#t�JgZ����o��*+5��Q�[x:��!"���ˋ���U��KK��I��V���݋LoyzB��8YR��v����;�Mv{~s����g��U��-;��8�T�½ֳG��)~3�Y�ɱ2��7(؝8�͑������<2 h4X��8`ɀ]&�.��ꦝ�D�l]U�;K��_y-+;�ܛ^�"�Ɲ���T���v��mnp����N��W���5q�o�B�����|�&���Om*��ꊎgK��JU�峺��#�*�̾l�)��:!y��!��{���';0�x��,	�y�_K�gΩ���Ba�ʗ�p	���\��u����k`
��d��+0}v�yy{���6߲�R�ֽ��ݾ�	/}H^Vc��� ��@�����<X�����zo�9t���,�{��E���m��jû{J:�j� �&�k|�\"*�o[8�˝���v�w/7����ڐ�`F��Ȃ$ā5w��f^��\�g�E�9�u��U�f�zǵڸ�9gׂ��FĘ��@�؎�J�7��+���Jjc{z�
a��llI샩Y��lG��k.�r����͵P*��'Nh8?&�n]a˻����ڵN�9����w
]�c�NV�\�ő���zU{}��`-(�NjA�,?9�-.T2��[t��e�uY�R�d}��,K�Df��ў˝�H��M-���]Q�.`D�u��8mLV�D*�Q���A!��A�˂�"m@�[���'��͗Y*�D�[�q�Fw<�Q������>ʝ@7
7$�R�_��������������{��;@��PL����ɞ�rlq��yƖ$df��+wu6l�_I�ή
��-�l�������*T�i�vO�S?1���\�oB�OeL�l��ݵ�ۯ�Bw�W��Uz^�#��������̊���s<�c�M���F�Ob��n1�Wog�Bx�ϴq���Lm��΅�}Z�k���`L�7�-�&gm?V��o餖vT�[ӿjF�����9c�_�#"p����J�E����>���u���*�p뭫�~��:��sT+����H�q���Ϗ�B{>��s������]��,���}�tǂ �0bv�Y�^�T�wU[��ו���[�b�U���d��a�~wWʼ�	MCt�nM�=<��;^g�?NXw�-��w�r5�D���V�E�Z!�%~�;�̅S$q2��,���8�s�^ӽ�/�۴f��o�;5�X#�k^��	i�L57����n�f	�+
O��.s��X��0#�= �Bۮ]^r^cH=���:0n*`��4�EÖC?����.�v�%159-WP����_����c�l,ĳef�Hx����ښ��^җ��QB��{���0;��ȃM�㴈�T ǩ���.�ejjF:��踨ò=���>�{~aϥ�̣���uh.�Z3�&d/j��H����뜭�;w��9=�%遹��k����;>�r�]��
�o=��R���K��gU���]9�ޓ��P�]o��S7�c�>*mK}���yQ��I�F��ٸޖ�J�:���͗�W����{��r�pw#<�*/�s�Ƕw�J��Ϲx]D\^O]x��z�E�I���>����.��G�) ����+��%u���I	gu�(ϡF�x��ʔ���1�'��v{���\o��:�
��w �������X�M2_�����}OôΚ�4e��P����~j�O�3/*���n��"��3=5����3Hb��Gz���u�(�߹�&I�1�~Wr��(tk.��o87���m^%�R�/�=>*���5�=�ZgTx�_��q�q��jHwu�u�5]^,a��F����Q���n�4%}�b�:4���O���>OE�%��&*��N�Q�WZUǖu��6�� ���'G5Y߂�t��Zk��&S�ث8���c���e�O�ǽC'F
�6�_"��q��zpS;J����.���@b�	8]^�G^��� 1���e[�.S���������x�ݴ
�P�]$i�͏/Nw/����7 [�;�����`��;�J�]ي�#�<�~~�����_��/������>~�dK�����>���	�+��-��N&�ç��>�CԥT �o>�zC�r~u�5SE�������>E���s[Y����/�foՓ��}�+e_ACZ1|Jt��}^���y���}�ؕ�.�Щ�% �"ial����ڭ�L̒���?Ѹ�=!^��FM�	�}s���_o���7=���9�˅%6*Oe錎|���ӗ,�l�`��mi�ړB���O�3o�	��{����<��i~���9Sbi���J�.����j����$�ތ�݂��Ţ��X3>`I�=��73nC���l������@���&���;3ͫPck%͵õ�g����)Y�7���콕�fu��r�N7ג��M�Mw�Nu��B�DZ	�%u�)�N�z'15]^�7�^��vB��C+��O�!�OF��u\�Q]c�υ��u�]����l���ɖE��.y<��rĠ�Ij;e�I^��])�#Of�'��"����\%]���p�v���A�VeEt�[�)�wq�#���x�d�,Id^�v��6o���D��N!�ݮV�Q��݀dH��^��5v���ud���Y�K��d_{��m��7��b���*Z�y�\���WB���}�����f��??M_�!�V;s�V7m��9�#��"Q�S��w%d"�������+b*���N.�W��T�=������|�ݕa�g�����ԝ�a8v�����ˊ�f��'����ks�V(ǾA���S��.�8Kӹy�������C�.���5���$UD�N�O!P-�a��� �].N��w���Y7�����ʄ7���g9K�X�y�i�ĕ�<�>>�dI�)p�DXSuj��߶��W��Tׯo>Y�L��7���f�-�࢞t��W�k���܆��Q+���EY��Vp���u���{��n�¨�L_����L�kމ;�5����A���;�{U�8y9pf���ި�~ó���F_>�t����^�U�j;TE�pIR:�1�C�ٳ��}���(厅�9't�4�q��t0�����nn��#�ך߯m�9�F�����&�$���	)7���	�R;�S�f�Q��g*)u��A�-�E15˲�/��S�m�'�>GI��WM�q�-Wy	Z�x����u]̈���a2:�@i�h ��"
�["J�^��b�Ù �(6�2Bv�%*	UDҴ��J�_�qc�2刍�]���k3>�b\rY�HJK%��)�t)���'�B%6�� �*���0L�u�$5f6��V0����;
ӣ�/�_B)9���7������}v����r�Um�V�_��+��:��s5������=b������*��=��3T�=RN�Y|KK�&�t��qw��>�3����*�4S��m=A�V�^�77�^�7q5�s-�2��ݾ5���j���:ff$	�(5r�"��3�l��.qE��잺�s�Y��<�J��YU�g\T1�pU@�D�yp��^Ҷ�}�;8��������^g���|�I�O/&�^��m����5³�2������㝱1��.�~�Q�F�	��0�;.Z���.���pm�\^�`L���w�u6�f����\c�j��뛢9�y�m$�k.������ؕ��������<��^����2�1y�Cz4�4Z�!UR>�Z�y��1%P�B�b®�������wT��S��х&�����l�-���Oy(��37�9k79�|�j��!۴�ʳ�hd��Yg+P����t��R/���O�R�~����V/�=���#�*I��ݫl㒤�Ϡ��_oV���.��R���lk����	��pɖ����L]��a㢟g��݋�C8��%��(���=u�0��3G��Ȋ'�_H�y��>Rw�{�=���n�����t��d���yR܇�s���,����;��T� ���GǺ7�u��Ҿ�Q�N���:;n��[ZW9W��p�D�uI���F�i8��0�Ȉ'�w�uuu�S�����e��=Z�֢ǥ�����0������Y�F��T��5�b��p&]Q�q��4����/.&X��&��7���5Gb�o%�z0�s�O�$���o"��ք�z����C.mq��N��������I��Һ�j���ٕ�,�R,{}�-ٽ�<�����.4���\0S( Q��QJ��s��D�V��@�$��RZ�;福�ϻE����;��i�ʝ��N��Z����T�����ي�1CN�>2���K�Kw�j�5���d= ��t��y������9y�/���TC�e��W)��Ͼ��+� ǣW��j�o��+mC~���;��f{��s�׫�yzwJ��oQpq��Y���U�OQ�\�Qb���\p��o�\�]�8YU1�˩5\f�^;)�p�U��/��{�N��J��ҨΝ�P,�i�]O5T��?A]N8�˷�&�]gf��TM+�#4{�(8u�^I�v�In�`ܠ2M���+M׬ǈ��n����k��M\��u�|a�|�U�SJq1��Bp��L�B��r۹�ĥ��U�cV[SP�S���rܻ��\�F��c[U�Y�9%*���Jꪲ����/��LU=�G��t'�B/�0�8�˜+��$��Nv淾�	��Vy���v:��Ƹ���������h��.��v�X8�W�#v���%�_�����UdEh-��/��"cV�B�YBU[E����y_,�����Q�}���-t��T{X�J�w^��S��YAZo>����)���$�v�wo�k5$,�e�H�{�G�U�Ԅ�gjK��,��K�n��m�M���E�e��ۿZ�[��������t�=�^�we�E�[�">�;�(�\�4��dqg5{�x �(�+�]�/�^��Vi��kY��5��;�w�>s0߲�kb����j���.3{iJ�(�t�<�)��ԯ�ƽ�>�{��\o�^ K'`*啐Ff��h�]u}���Ux�lo�4k�|�M'����8�K��a��|��g;�G�x*���6�Q7���u����\����ǡ*}�2q;٬1�{R�Z�<�U�F�d���69�yA�.���JSx��aq�%��bz`\Fݲ������7�^#�Js�����O�?�ow3n1�LN��9��7��:��Qvj���Lu�z���g����U~ʾy�eD|��ec�I�7:|o�j�GMp"���n��|��d����bU����\?v-��r){Y�#������t��
��&W�P�E��{S�AY���EUG�ՠ���k�O;r}���\�����)�7w���s�fo�a���鲗%~����&o�+W�`}@��������&�������Ve��"��&����Y[���!�������6�c�u�G,�d�p�L�_)�o^q�]����8Vn�q��+��s� �=�պ������FK���ϼfg}����eo����u~77~�Ro����Y�������UO�*���v�y��&�#���^"/"3{"yU�98��zv�]��U��_����s>��u>_3ﯴ��k�g-r��(ynu1h��+<<�1�{֡��Fl����݊�P���֌"x\^���ع(�.��9h����#@��^f�h.f���ه(lV�:��1��5��ttZ|Fe1�������������Lr��?O4VJ
Lg�G�b}���w+~�SNu�������W�ҏk�qB{9ZF��F�Xw9�N�C$�y�N&�S#k��V_�J�;���f'<MRj���w����~1��Q۲�fv����Y �f���0B���Tw��^�6��2�
j]�٥C|��Ѻ�����6���2�j���c%��y�q����@�Z�� b�B�Z�OMT�C��!��ţ'�������P`�jܑGy�Q��w�yu�<D��#۲�u�)_c7Ef��V�}��,��J{{��ȶH=��jɅ_��@�Wi󛡐�X���u��Z{/SR���{�����Q=֦��N�;��50��뷝���up�	V*{���/U��Kd�D��UZ@�V/d��޾E��;Ux���i=V����w�9X���?�v� 6��ufP�{�9dh�[�����W��z�
������歄R���|����n7��9T4��έ־�t��#7NWM� �.yZ �qu�m��A·Vn6W;�ޏ�R�tڝ��u�jRV���R<�v���p�V-�yh�R`�OZL>J	���?�I��rr[�m�L���<i�-u����t��`�,c���#$�
�y`˧i��nJ�s�d��G��1��������m��P�b�JJ��*j�k-mq��rwZJ��+�:1\��Y �:.EJ3:_Y������Q��5����À��5���L�����'yⳏ;q�2����}c�켠��"`��,diZ��^��wG�;m�Ԓ.��Z.��8������kv�
+PN:6�-%I�|�P��I6��aMru0��u`�<d�j	��9*n�� ?��"B���);����[*x�*z�Og֜������D�Ac(P@#�[��;{k�V��ۃ�&v��9|�b���+�Yak1.yF�9�^^�7��MM�E�-�]�WKB��_Ax��])f͵�e�N�����W�(�˙�%�LZVP�e(�;AYv!���n����4
���%[Su6#]na�Aĭ>�#Aɭ������V;1A"�yrLTimq�'U��r��]�m�e7@k_�tsyu*�B\d{b�8H�g����ƭ����E �,�k�u��{��^��|'��uk�T
��e�������:mx1F�md%^���$�F��!"ZܒI$/rY��q�A�jd1"�.$w_)���0蟣$?EA��.d��IM�|	ڣ���,f�Y�����&i�aWcú�9�&�b�m^scŦ�!bXf��mM�pso\�i�f�`���x���-��̨-��J��&��3mu�i�H�*�@�v�&Q#�n+q��8��SSe�U�UV�m��0�e�݌k,�ᰘ9��2�c�X�w��jŞ�l�����͆�!�����+�ڥ���p�j�l�3f�kW��[&�>����][��1E�j2)Wvj�aqi	�z���AR�܈**��+d����B�-1aR5']F^
�H��Q�ۙ� {V���u9�9k�L��NH�L���ŏ����Y��QPV&͹4Z������qوJb�#N�4���"�M <O�;�� ^k�I�JL�Ú=�vT[7$��9^,S��;�"PW�y�
�q�b�K�c� �^;����R���I��L��U��Y!%V��ͥ�T����w�{���S��L>�͙d�^�[�d��s�`���� I%Q��q_��7(����㌴�.60S�����^���uX[G��ڄx')�T�����6�b�HQ��6�=�謏���[2�L[p�<+�S(KH"�H��(䮵Wd|*o3$�2��X��(X�An[)�%�*ʫl�xJX�n�W�Mm>��U<uz����d�Y�T�:U_���%�(��;>�K�����U�/��
������>�NT!^�1�,κ{��2,CG�Ǎ�\������Y�[L��Bj됲���?۵l-xa��x�>Z�#yٙ���@��\�*x��^�����z�}�����f,MW�W�a��Wo�ox�*�W+�\Ἴ͞��`�~ �69���i��o�F�ix8O�N���!P�B�ߏ��a��3��{}�}nb�K�$ۢI�ڥ7�_q�ĳY��=�5B��	��?�H��hL�`���,�h�a��j��ߡ��*�Ǡ
�_[��?EUt`������#�D� 9zBT":��-ף��}��庽��vTj"�͸eb-@�U��b|o�o¥�;���k���O)qk�>��F�'�C�d��Ss�c����-�T,x]q��f�|��^�D��+#��5Ң���X� ��O"{��T��5%�����h��(�"��[���ZGeԑj~�Ĵ>Q�z�h�V���r�O�����������2���yk� ?}�'Zѡ�<U��S���=�?�"L���/�ܔl���ӭ�=y�l�5����3s�/@76��-xV
��ZtF'~E�D(���A���|�;��탩�X��`�q�����3��AA�ᵅ�6�ظqŤu���{��Y9�C��BCT��V�Zs�N�sdX����;���~�8�����*%EA�6�:��t�G�f��i�3�l�病����Rm.Ȥ6"�mb�z�A�9���mM�_\U�||7AS��c�=�cA�/�Ά����E��jy��~����ת��a��N�zbt�!�N��{+��;Y��*���>�� �"�HW� ���B�xR�޼�O�vF^���k��=#�3������}Zs��I�ǹ:�^��2�|#�;����>��>����I^�|M�dR&u-�h��$47�H�J���1���g
���5���iK�ۚ}~�O�����65���y��� *_c�Y��1�9k�]�#�j,�l�/KA�n�M�K���STBN��i�rB�ܝRbﺑ�z~�~����M�����+D
�5���F�Ѕ�z:r���8���˛���ķMj��*���C��t{��G���tv;�H�]�"��Ӻ����#�]�j����Q�=fn�UfK�p�8Pw�ym�,y���}䯨Gz��CgR�I���qf<S��o �Y�fv,cmҤ0�
:i�]���^Z���v��v��{Ӷ�1wC~�t=P����E[GFnnAw$v��ЏU���N�',ҡ�r�Che7�]ݕ��V'xe&v�e������൛lm��f�\ ����\[Q]�N��N�m-"���w�h$���^���Q�Q����Ɩ��xT��;�1[�
��>�#��f��?GEq��VY����>����F䲇���Lz3;��5���9Z�<�	^D�~>��0�yn6*�uf��D�����˅}��S����pD���l�@� jq}�҃�W=Й�����{7{m�j�q���gyT.��J7�p���&EH#�xt��@�G� ��x�Dx�N�P�߮�H��~,)�Y����v'c��,V����$R_�����?n9�����(|��Ǥ"��L����聽"F7��휿��U��߲q����I��3Ty�DPש�Aba���s�~��)�S鱫��<��s�7�]����/�z��9����5rb��sU6_T��U"���9���$�G��s�7��/\3#U����ћ�>��e����^�'N� G��qT��Ҙ�W��|R���w(�������7#Y�.'�A*v�7c��Q)JS??_���Io�U��}�
�
P�u��e^�f6$=y�۩�H�9,��=Ly݉��h��=_k������'6E�ǝ��0�Vj;��u��L:������;�v�S![ �c�v�mXH]�fZ�_ݧ��[ۚ�H/�>Ԅ����3uևY#_Ì���3ʝ��Q�[i�tgJ������:E톘�]H^�iV�1uS�=b�O���X4 �A�����.eЊ(��&�}���tj�M]V^v3U�r��f��&s'į\K)U��.mb���@<[ ��k� N酌8�'����(�\��8����:~��Y54&V���y��ͱ�O�r�&h6_{��ϻ"~'�z����9�����N�sE;��m�a�����N5�b�>�m�H���Ύ����L�@�_ZV�ҫj)��K���{���!;��xb��~�Q�\N�seo����N�@�z^l���O#�h��[>�⒗0��73���uy�,����zU�F���m����nk+���>��j�'W�Œ1�{�#�����z��T4�y5̺��&��>`�� 4Hk/7}�����V�rs�y*��j�uT���qSR��)���t6!��Vi�e�Fo�˽o��}��뵺�!"a�Wa���	��+�|ť��z�l��L�������K`&9O,o�g���,���*O��ɉ �y! p����Vg��$W���^&����p���g�����ZI�ۉ�i��6}j��Q9�R��Gs���q�j����N�;#-�j�zo�e�(���7�+�h.�%�x�B;^)�Q�yp�Rwm�5&Q"��|N��:�^n�wN���*�֚����Gw��=��:���K)P�PD����%�F��k%������jL�:J��׭��1���&�ߊ���p1��J��*M���Bh�ܛ �C�&��v�����T�TMR�C-ِ �|�J�q��<���#0�\�f%��������'[�'�yx���m�%ڒ�B�
U��X������_�1WJ�K��<E?��Qö���J�뎯}1غS��g�`^\��o��>��a��~<�z��;W��ޒ.��3�fدk��t��o����ߕ�h6\�ʋ�x ,����Rq��|7���m���R�U�g��Gnqh9��	�]�*���g�f�=yn>�IS<�{ z����Fs�U��P{.���нbЯDL��fKD���W�{��2���4�4��@W�g�|N�s��Х52�ĸ>��|����ΝK�^>Z�T���h�S�J=�02=h1��a�@5§���<dgzLu��I'�O[�~0�W��i�#�Ǵ
9�Ϣ6z�����7)Y~�d".6uޞ+;�|c�nv�o��b\����2��W�*_v�ɑj:<�D��u�ş�����_eE�����~S fi8S^���z}�e9��I�wvb4A
�ɍs�}+-��yyF�r��o���xl�<�;���f�⁛�=���|R��U
��Ad&B�B����?�j��b	��O�Q�g����F���������­�Yu�T`oڽnf܉3)7՝�r
�e�E�z�TL���,�>�ev��󀮺�Du�C�T�O�K��`ϝ��C���rM��fh�����_t��.�Ǐ7]^�]���U۪�x�E�"޻)lL[ۛ1�a��+���\z-Oy�e���ݹMS%:��LiVlqs|��K8�԰3�2q�P��Α���^�U�1���Mu�l�n���a7�����K�/x{dr-(�Yǯ=�}ؗ)³s�s$���C�r#X��c��;�����gf
5�'�K�d�li��D��Z4�v�O���T[���3���ν��qs�p� g4Ս��A��&6��-!�~2��zA��iJ�y1�E�w6q��N3��:+A�ߴp�\�3s� iaZ3�Aη�}�_Jφ��
��;�O_&��]���@z���^���^�NN!�5J>�.�L����c�\������u����2��w��垽� -YMf���c��w��/ �_�z.2]|	��DٞE��=C�c�m��?k'���X
� pI-�$����;>�|*���	��T@��ۇo����7&$9âoG�ڍ���������o����=��HU��i��Eo��OF%���������+"~y���C5U����JP��>����xR��S�`�d�<����Zx�e �������\�zc��}�n��8��B���z����4�}�)��(!\�^�_R�eTF�V�*W�Yv��>��lwDL��#2>7���m��eb��,`�<�eh�h�J%P�d�/	��/@م�!�\n91eDmkǍ��Ү7�7�'\�)\��W� 2P�\z�-w�
�	��9w�[�5#	���25��x8.-c�)������Y�x<|nЖU�Q�.�!|�g6�T]�˼�%��=_F���k;n�'���W	Ŗ^��U6�v	�L52�+F�D߁�׺����<8�T��&}��W��.��'�<\SO�z6�ɀ��)ҏ@ˏI����$*�Y
wy�|����"�׵C5��9�����Y.��_��ְ}8с��*Z��J{�ר��^L�O�w-�(Ⱦ����q.�ݓ�nPX������Q�(`��`ST��(�ܛ��!���uF�Ow�tm�>�>m���Q�C&Ц�AJ�RE2����������eB���]�?'�����ۍkkHcs�ڢ�yI���C��B��={3zf��v>����uwwA����b|@�5���.���~�#�E.��
?�-+����'_Fz��x�i'�=���s���&c dC�e5�9�WbB5�c���[����)���yf��hG����l_I�O=��02G��w�@�M�ºa��6�>6)�絞��պ�P.�q�����X�;�&*�z).W�v�*
�M{ĉ	�qR�օHUN�~�};�>ox+�Ou�8�i��m�����5�Di\�}�U
������ݵi$g�C�P������{��D�9�x~���9�pX�0�k��Ɋnw��,}�tv�����p��+-)H����Cȝ�d�c�,����/�[T؆���A�V��`<쥺����q���n8;X'<�Т�L������v��Jnz���-5�-�z���GX�(�s�?�gn�"���->��z��v,ր}勲��6� �G8�g'������G�OaFA꫾�Ǎh���ʇ�7��w���]�/"���u�]��c����>��f%���C����x���y$Ă\ ��'ЕF�PQ�۱�H4�m�rr�Ӈ�E����NJ�&�1��sU��� *|�f�����Y��4��Ӝ�y�Ͷ�����`zf����N����X�z_)�Ōh����G��z��n�D�nG��@JS[}�w����V�6'�[y�hW��LD�z��+ywq�{3�#��C�����:������<��Fro#�[HvN���~�߹���ÇʾYB�	��_�3���s�賮>|�>��yi�#t<{���|65�l����.	�4�<�0�z��̽�UU���9q��g���翇�n9�Qs\Yd�����'��c؍��&+{��s�ބ���ng�%�����g���o�nnw�C�������9�EkX��	�N{�w���(�.t�kO�C�e��{�w�jq�n^m��ﱥT���"��c�B�����]G��#�}=�<kM�u8Wޜ~hEd�}�(`�.sg-��)�?��N�h�9+�pO6Jd\�X���hص ��&M�a��td~�;h��T����R���)Wc-�;X�S����g=�^��QJ���Rą��73Y��Bw��D�>�|�a��kd{ ��(أuQ��&�ǿp�L��"�lm̈X���#���+Bh�(�f3#���B���s�c��c'eů�U�ás�"���_V���:t�4Jl"��f3|�\��(Q
H��vY���K��_ñ@�C���9��n}�y����?�LT�Q~���}#.7�^���8�ͼ����B�E�&V����8ڵ��Y_f�z�i�����)z��>�`�\���j�Ҡ+��؏�v�����}}�>.9U�u�C�m}f��+8d�����s�莘�ܝ=��x�"!�9���9�f��_�%b+_��Z�JC���Tzs���Q��⢣D�5�������o�ə���j}b}��\�)Rb��3nj"|�z2*���^z����{}]���{���޷�W�8��~��g��c�J���}hɾ)���K��m��y�Ə���~�	��T����I�}O��q�������gM﷊�i:C]��ϕ���h�����.%EC�w�K��,��O3wDt`t��p�q���kҨ­]�8�e���"��w���|���e���t���W���Y�ۢ�����L��2�U��R�ӕ�8�*�U������E�(K�&ȻQ��>��7꼻sFp���ox�{��ק�Zi���χ	�:ǃV���e����s8=; X�6�����]�����<Lv=��EŊ}z]AYӋ�9WEZ�b]L�H[��Kz�+qѷg;k��IֹN�͎-f�D��o<j����>�r���Z{�g��[-7;�~t3V�[��I��k��JN�HY�/��WU�b�ߟ��*��ە3d�8��e���W�.�/B1/
����6G����lz烣�&���+ƭа����d�޸�z���,]�|��z�,��<��s��W����z<��=o^{�{3"̱��v;���s��]��cK<�7�}7�Ɩ�/1�����v*����m�2<����>�\�3����fb2L�u<��A��s�	���q¹W���^;���q�y���?!�9����-'�+Þe(p:t�{E�k0��L^6}Q��Dϻ�1oѼ�6�ĉ�߂��s��G_�4�c����b'�:TYA���,cеpY���\6d�6;��e�U�cti���w��Ư^ \a�"i��������ǉ�V�g�]!�ft/��}@�ϫ����ZCa��וbܙ��1b�)�Gᓎ��s�e����(8"M��CڥDg������7\m�@<Ûȷ��,�cr=�٘����f��L�bYT��0�=����JgN��Lh
ž�;�����(�ƶ$�=+�]r|㧰��Wټ5Fqh�j��§Ύt�>9ɝ�	؊���k�X̜'�ZN���o�7��7�+Q�Y�M���m�A4	f����4m�,��E��Y�lj�������x����M�ѓ�+�j^N�M�4[y�l�Wq��y�)���/"B�K��P;�%Et�N�}n�<K� _,������'y:����s�뭮�JspMi��]�2��h�����sʥh<��v��qiwɇ�0����N�v�!�7S��ۡ��t�[�ƛ;���z-�Z��:��d��Ŷ��*�=�Rm�|r-̩q3�,�]퓂Bc=F�R�^v��H���L�tw:�3�i$+�Ӭ������=���|67eS�r/c�Q��XJ�<-����J	�]/�t]ݽ�dcl`�`\��g�U�_V�ձ�7��N�ٌ�w̷n�S��7A�@㮬���+U��b�wGLFc��L��k���E�nK�&_Gf����uΝɱ���F�J�:��/�4yl�U���}4��a���.�K��&n���O�Ⱥ��7�6�-ܔ�U�1n�oD�;�5pmr{.jk��aس�������k݁�C���,#�q�T�q�[)E��D�ʹ���ӳ�SbU�Mʖ�Ĭk�����k ;]Kfsw#ۨ�7�n.��	�J�*�|��ۛO�Ѕb�\�z���Ƚu�3Y���/��ѤfH��ؒ����39�Ut�����U��凹��k�=^�U���(����]��]3}u����P�k3��t!oLF����7r��Ś �@�z;c�"�p#ybS&��H��J�$I$��F��$��%�����vu�y�!��+��"����U�XOM)��T��zh�J$�-풆�k̊���3.R$N/�\d�[��#���(�,u1(i�����M�5��Idg5�{��\+�v8�Hj�j뒃'eq��-!V��ٶm:�K&Y���f����Vb�R����+�g)��|����g�(�K�<�<a4���ٚ�Ȑ�'�����U�%���fMh�mm����:\��)�>[�َ�'j�`�z���N��"'~�r'Ԟ�L���)氞���`�<��a«�I�ڇc��6�]�R�4T��T^~��@�E����*�V��=$�y�W)oa�l�K�z��Ʈ��Y5t��{��F���r�0lg��gu��Wy��;��ߦl�$�]B��T��ߩ��Թ������#�ۤț79�Ϥ�K럷;˹��	��|�vE:�q�2S�^���OSt\�~K�)��S�dh11��輽S�����q=���vz���$�o�{���]�H�'��}O�D�f�ږ hz9�D���?.�#�WZ'ƀB�O��KۦP��o��򉋛o˓Z�hR6޴�*>Q���q��h��
�9;����o!.!�~.bk�(��) �<X�BRl����S��&r��R����:�=�w�ݱ��/��~2&����c�|�U��*�������
`{f�P��Jr\{��F����xj3$̙����܎~&��/�,���O�5p��y^�u
�q����� c;�>u�u���t�p|j3�Χ>�u� 5�C�z �&x��;�8���okݞC)��o
~�E��2
�/�_�;�l��^xQ��y̯d^�� �� ���ӆw��+�3�E�W��,TȬ���^Xs�f���20��:�v�јp~��s��Հ�U�.��!_�=@�(dFE�9�р,�w��{�%Ⱥ�>�����M7N!�șT��W��e��@�_U��q�[��O=�z�d���n����z�7������u�	]fv�4�ʟ�S�=cq��F���
��hQ���
k��*�&�X����y%���E����`�V�q|>����,&��tP�'��s��5�4�*�Z�+����j����ic�v��d�O���@wY�	�[��"�m{Nˈ����	���{Ϫ�^���/��Ѐ(����9S��J�7�P�1\Q���nU�~���xY���9�n�&hz_M/n�>�\e�Ő��8-��k��1&g�us����@z�6{�[t�b�z�'�1Ѱ/�6�����i12%M��g�������9#��-�������y��F����NH�M��S��&Z�N��,j���TE���F^����}��sw��6�c=��P�|��z>>���L����.㝪�Y5װ�9�Z��~d���I�:$�T�u�ͬuǇ�4�A��u�^����ra���bc��+Y ��m�U+��J�\v���[[��߷���y�Ў�qQ��P��3�7���IS��ٷu�j�^ɞa��b�-����]�f0+�>���+
���M܅�D�F'1ݤE�5���/�']M|��u3�������%=̾�q
��o���r'o'�[;;����weX�����ֺ�|x��*7W���Z��M�*VU͖����f�:��T�wrdyRH�h_�u2�dV�3�k�&W���Ej��ӻ���	�V����㪫#��2گ�\�H㚊v��˿Hy�b�n۹MQ���]ƉJ�`c�嚼���eЧIe8���n�c]%
	�5�����jTt����0a����c�Lr	TV��0��b(Ѕb�������M1��6�o��7~$�~�KE���M�n'�!���R��5r=d+�g�/��N�Uw���!��9lYC��������v�A3�y��yG�Ls|E2"�:⧰ƨ��楷����|-�. ��e`iǠt{�����X��=>�� ������J 2nL�uW�؞�N�1�~]�f��n2�|"g<��ɔ<ռK�&�x2�ȷx|�ш��>�y�|= ?eyN|*RE ���{����DAn�LBI���5]��N�(Vl�N����.����W+�@>���'ɶzO�w�W_$�v=��RQ5�R��)X7���2��na��]:.�����C`_�yT�2��������>7�_�<.�>�>3MxST�CC':b��*��J9�a�=��	��I�s}��|bwW��������)�0���]�"��3��*�ʘ������>~m��n^m��"&kvK�a
��Mr�HUm��4ؽ�r�K^,���pu���|@�M�Ȩ~0H�JL�X�Ʋ��K[w�0=*I��W�&���]���K�!�3�N����Va%��L��`������fF�N]�I��r<wr�����B����ݖm#�鱖\}q��۟9M��/d��2"z���5�ŋ����3��g�����b����b����/��ӷ�����t�����NIP��aY���L��oV<��neU��]�t�0^s4�Ӭ��;"d%S�}��U�J����T���5��/��͟|8a`��`�@s����&l��̽��Gs��_/���6߳lE�"�~�j{\�wls��6O/p̃S��5��d�z;ơ�D���������ϱ��7>��t�t��h�����{$^wg�Oܒ}�xkޜVD����y�+��Nu�D�#l=L�����ǁ�H]�W�X,�r�g;w�����Yn=ޚ�m�v�S����*
f���yώ��G�y�`�_o�S�����z�W�s�=�Ӎϭ���$y(���oq�����}��H���:~�wz=�xu�m<{ؽ���Ī�����/F���䣭MD ���VO��>�#�t%���B����3��ȟ�x���$�@] x�"��q���~��h��&F��h��t�(C����5��7>�-�w�(}h�����A��O��x�!sh\zy���l}�*Lz��Y�Fo�MF�崃��҉?xVk�;��T��b~_��۞ή�s8�X=C�F��xIu��]t)NO�w�1VY���f��E5 <��]�M����;��G��"��wN�~�ɴ���j���	��>�A�%`�ԃ�q�1�㝣�A�zu�{�#2W��߱~ֶ��F^2k����Z�f~�nc�"V��~�ő4
ʾEF�۫|�����f�kv��峺����9��mPU����ѭ�G�-�Cu����\Kh���R���H����5��w!J��F���;m��[�!�� �YF��G|��fS��D�[������*�.�z��gk]=����Z�骝�e�޹/쨗8��<0��wn#l����&=���ͪ�|=8�y��ݓgR�a꙰�4������"2o�N�C�̬����QQ�`��oq&��i����ʼ��{J�:���п�
�Ņ�3s�����e�5�U��ҽw��ݫ��9�e|<ˑ�sq����η�[󂾅Vl6�RR���D�D�dqPj�lw��o�b�}[�1�>�����ra3��R��z:�P�(ܤ��K�~(.����c?Kwԯ�/��i�z�9}�]h��uC�#r�����}�����\�ϯ1v�\��{}����ʧ�:'v���Fz��K��#%�>Y��t�	��9�J:Ko�^��{�����=!��R�H�_E���³g�oޤ�,�ub2����r��'�|����m[��Ð�
>ݺ�]E�+�O+�)3>����"ҩ�1�x� =Oyu�]}�5.�[������g6��9~A�@�i9tהD)�������p��x�~$�1��&ݟ�n�G���oTȄs�|C����OE��Ls�w I�1�aZ ��Y\4�p�Mf�24��<��:nse���k6�<���ǀ��D���):QgN�b�6��W�E��bw�sW�p>��{�/P��{�ޢu�1�	vE2	@��u|m 3��C����}��Q�[�7���=Xv��:�Ud�����B"z��=��ѫ�s��E@��<*{W��鴀���g��J�Cg���V���[��g�͐{	��s-v9m�n*��������~����7�����9>�Y����^�5�){�8�I��6�I�t/�ҍ������7s6�3K�s yuI�%�(-��B��ƕ6��7�����#K���U����ּ�Mu3lM�21���wD?OS����f*��ɦ'�zL�`�ɮ�Yz�ӫ4����w�D��|�u��{�����C�y�NJd��B�u2N �>*{�6��F(c����y"��;�}(\P��}��0��:����n�6�T�}�,Tⱙ'{�|�|h<�+��@љ�����zI6��8��Y�}���f�<�o�%��L�E�//)�F��t�ֈ#��V�W�+����b����Q.⣾�t��n:�Gr���媌��u��ޢ~��L����� ���d�!��k��wV��5�(�<�l_��UY��1�>qV&&W���a�TZ��Dl�B�Q��	dW��܌��5�	�9z&�������aU��7���R��cy�����N�3�8l���S�|Z�a��:�T�˝�O&�[�v�`D;��I���F� �c,�[,��^\��r�Fnꏷ����{F2,~᛬Mf)th[Y��׮Vs�]6�)-�+Q�Fr�p[���Y�&B,��j9�QɎ����n2�j�UV|݊��"QU9�&$zG��%���Z�
��-��3F��;8�n)���y�^���`�6�l�����d"a
�l%��D�C�3P|� �X��ϥ`��	�D���چ�Z��<0J��X�l���A��#f}bu���o���%yfN���XԞ��sz�|)/`;½�F���q��A�&�P�ZUY;3&:�_��F��#_;�~�Z���;���z�w���u��~���>���f!ּ�#���{Ic���o��w�*����1�-��NJ��Lz"������7�^�\{?���_¯�e�b��_��/s��7��1�U��`㟹�{���v��>�L=��D���W�{u/�����)Q����d-��*�~��k���[�Ɔ��Q��Ǎ�*�|62=u+�:F��D�h�.�z��S "�ؽW�_��m���y/��W���*�G�ˣ����sT����1F���3b=Y�:�ޣzT�\���B����vl?=!���Q�
0�nr������o���/��7���9��L����G�~Vn�aҠ�"�Ts�M�YT�`Ұ,,��݉�X�x�vbL���t�]��Q��9����bQ�������F�?*P1�� �~�Jt���y�aC�7�˄�5	qxQs�(�7�^�.����n��H����$���Y��{p�������O��	�(�Iw�O��9x�
]ҧ`Eܹ'NAG�QQ��(�]�]Vˠa�]��a*�zo!�)~.��n9���WVowN�y�)#�v5NGo�����h��̺D�h�O4mz��l<�Q�ޯ�@����"'G������Sk�+�C�F["C]�G��b�q~��_gf�o��'�V�n����n���^>�L�D	�ь�����s;���Խ.�|�r�	>�{�^�-:���`���۽=8��à�qS�r���dK'W�#�pt��]+V��	���P�����x|d�@M�t����_J�!��>����R`v���EY��ɞu4�����kT�Ѕ��^#�<��!�~>��;��an���$<��z��"f��آs����N����� ]Vz({�M7׽���j�$�3
����77�3�)��r�^�Q�����b�_�؂��@5a�+~�x���	ܢ▌�J#hv&�d�X����q���è��X̺�X�����.��<7j�� �Ϗ����FW��L>�̍P��]b�s��f6���=�k�(�fo�	3<�ޥ�Ѥ\:̊u�U���a���6��05

���0��&���H<`���ٽܬ.DT03��c�;�H�ߐ��@�j�r��̓��;m��ډ>'Ș��S����yC�v�k���kB�:zq7)t�z��h|@^�Ŋ�`V����#m���;n���..�u�' �)B���Y���x�T��lJ��#M�n�q�7�+{&�9���5�Ġ�E�:kwf,OdՔ��j�>c�-������#��זo�L�1�b������ �7	�FS�R|��Α�fy��]7*��~��ƙ3�n�@�U�E֓�gߢ4~�'��k,E�	|���s��3v��Q�D���Dh�9',먝c��dS^u,��ș)�)�`-�WA�0霳WI��~ޚ�~�Wl��ٮ�o=��>^�}��.���wS��қxG�k�s>��� � ��F��\ob���YC�f`�������� m�*�J�H����
/�{���|�U�b�>ň�4���ߘ���
�������(�.�_p���I�w�M�-��&f���q �U�sӱ7�Av�vO�$�}kn���lpn��a���R�"ͣ���e��@��L�A��L�fR��߾��@Z���F����+�l�c�J���fo�]�~v�^��6��{&f�x}�l��&�����?4��B������9w_�-�Dw��F�3WQ�:6��/f����izе{Z���-�wT������ɦa&|�`�=��N)p��u�ь��z����e��^ɟ(i�1���K�z�ݠ ��Kw��6z\yFe+�L7�:e�.��"�+R�*�����f�9� �C��c�M:t2���.�c}���c�NP�9��7��0��w�@q�}������1���}2�nYwi[������ 11��"��X�L��*kz��Wy����=H�A�9&:q<�/��l���'֧�3T#����~�@w%�o>;<�S�n��] @�E,R@@���4H�]�!+-�����2<���}�K�p�˕ئ|��Q'�G�]�Xx���~](۹"�h�vmKRlݢ��RU�TUf<��$��y��Q�jKnG�fP�}���F�E��?�e١��E��9�M�Vk}ds�};`��SE�����%l���a]���F��Q�Luu����EA���>�f`̢�P�1�R�{�w��F�B�|)Kͫݡ�!Ϟ����_�u=���ki��=�ʮ����Ҹ��G� D׮�:[��2����ܯ���{�J?��z�b��Wnj��`�*R��-ʒ����$6���D��1���g<V�I�KuUol1&}�N���ؼ��d-��S�����I����DW9�Ju��yS��Mtzf�[�����������{��u/~��ʧ���^�:�\Ó�B
��(��p�P�&QB)��Wz\o�d�щ`!L�v�&Y�x���G)N9��x��`/d�t����6����-������(��������w�ȅ�
D��/�WC
612.��!�$PC:��R��P�@"�*Q��(
c�� "��"�ޮ[K^���B�*��Z�=�t��_����������7�ο�'��_��hx��*�~�OQU	TE9x� ���!��9}~;P��P���_��(�*�?�יÑp��?c#���wO��ݽ��EAPA(""� �*̫�8�?pQVEq�[���׵������C���7p����D��^�}?-�y꛹=u��2��>�~V� ��|`n�vz�{k�* ��QUo��lQAh�Rr&DEUp����R�
�OB��w甔ib�(0QUgc���DAU�3N�]��߽:�������6��k`��" ���ۡ��ӷs�!�����B�>~Gn}26���������m՚�����0�hn!�9�|�e���oM樨"����3��F�QAz��);�>���d�MgnF�� �f�A@��̟\���x���D����U
�@AE*
�*T"T��)TUUR�R��R��
�U*�R*��R���$v�2�UT�   �                     
            ��      �Wu4�+x���i[���&��MźRͪ۞�{m&�����Y�7�ܥ�m���Pir�٦���3�kk[6p {�]���ۡ�n���e9��R�@Ov�<��Z�'J��$mw� �U�
h\κ��
��5�Ԟ�!G��/l����^V��yx ���y�9z��h�:i�(�m��G����P:롪��`�x         7���cLnp�x�N���@בЮ� �yn�y4)v�+Z<x tR��r���vЪ��Pz:�<����E/3�4�r�km�R�� ����U��u���J�ӳ-��  
)Zۻ:o�l��c��Y�7��K� ���E����-�/m��nQx7v�^;w��(����9{2Ȳ7 4w�uU���{���n�����mD�y���ӝ��^<7^�����@ �         ��0�V������;�w���v�u�ۭ���g�K�x�zޭ�f�� 7:�z���5͉�V{�w�,6���9U�=�x��z���x �͵�e��ކj1��.mX�4m��k4�nֶYe��=׭���]o :�e�Eɨ���j�wvT6[Y�7T�UfN6R�,�n �{֪��/m���{�����k��֖���^Qm� 4�U��         ��k\[���)�����kZ{���N���m�l�=�(�֪�����6�=ۼ�D���m�w[fQi���^�^� 7{e,��n텥��,��(�
 V��z��Y�ۼ������8 ��u�m����3������,U�nٕ�Ms�w���)x ݪ��\�u�Mv��w��1�K�\[iM��:N�i�@(	-�p         Mͳݻ/.�S5�=�-��[�f�=1�o=����w� ��l����+o]q������v�<m{���l��˶ʱg� ��m[m����Ų�=�Q@ �f�n�7u�X���{���� n�Yf�^��<k�tڼ���Ŧ8���b�w�w3�s-�< uW��m��.�fZM��kjUm7��uK�:�f�)x'�R� 0��D�*   �b�   =�� �� h�A��@��m	� ���$��hF�4���@`S�% ɫ"��mh���P�҉�,���_��I,��$S�8�bIff\ŉbX�1<K1$�3?�%��Y����I,�ǘ�,Kf-����)�5o�Mme�L-��f�{�X������b���+D"~���WUм��)Nxo�WK����e*p�C�ܭP�"��� �/��}:��!@��QmM������J�%j��3���%�waSN�}`8�-��<�����̮��\�"f�Z���i�Qi�@_B=1��c豸����F��ѥ���T>�]�c�G�E]�HD�V.�z��W�7��;N˒��0�/e�����r���.��F���i��8��-squ��\�N��˹��Yl뼧Zi�b
�����n��zi����~�aǷ���1�\-Yś����M�ib�1�ǼxSVr�v�h��ٷ�L��-ʠ�B��[l�a5B�0�a
j��W.!��Fq����,U����
�o2�[�r�w.��4v.�.��E_�RV y^���%%u��rxv�0����1@U��6�Lօ����ݼE�x��j�Ԟ	Q�,VV����<�iݧ�MF8�!)�B���˵�OD�B�±�dn=̧�ŧ�ݑ�܆	!{X��w��r5��uf�l�cj(k=u��`�@wWO.C���ܹzrW�@4�/Z�����v0����A��8����˹w�LT!�l���_�e�Q k��)%虱;ݲ�L�����̦��
�yv�fe)�%�Y�H��g%,�i��n8��h�D�kϤ:\�ͣl�i�H��(ضЕ*
�I3:Ve���_�jҪ�6����L���� 7F��Ԭ���F��`a�#�l�T�\���;�%�Z�6X���
�rr�F���;�(ƝX��P۸K#M��՚��(G���32Gf=D۩�d�ISlQ"Jy�� �WZ��P]��Q�������H�g7R���(�\׸���&�-�� �L25��z1�r3���U��N�B�m9{.�˩4o,�T��iYr�yPe ]u�6$�&$ve�(�,��d�r
������������R�9�4�[7-dbb,5�*t��M�4��F���M��0P�\J���%�0�T����@�-�zd;�@m�2��P&$ͬ����ޝ���[sB�+ŕ|tI��u�M)@���pB"����S���v�Ʋ�ݪ�:�j��]��S6�[zr�IY��[ 7.���D,�m;��m�1hq�n0�xj�0#�Zf�A�������ɘ�yYy��ݧ�n��'[�M?[zV�5��_�6����[�ͤ�li�-�6�ݹe4cɨc�𽘨M��R.��OBr�fP�q�kq,wlX�N�i��Am5�=B���-յWX���ԛ����0f�v��Y���[u�յ�%��tZô��:.�����Ӱ�(ʉ��;�ǂ£�C�72i8A0�zĆ��3kn�Q�Քd`���(���w�J���:���,k�jm,��z�.��ټ�MGsc��P
�gj�{����b#�-G(���^�MD�
Jlax��^�ma��i�{Bҽ���;��EemUţL��M���hT�r���S�v$��B�3{K[טS�p
ؑw5^-L����4�mЦt�����
5�Ǜ�*�n�Br�.Z�͊�ǣ.�ލ���CmP��b�:+o\����k�o2c����7krj/:9��4Q����d�޺Bʆ��V��j�X��2�NJ��ZwC0�^n(�%:�
<�*��Iy�F���e�\�D*��6Yޝ����YDHP�0ncX���ɡ���-W���ֽWv�ͧ��)F�ǜ�o1�V����工�`�0���O7kYzi���;�).᚞
{��m<�:7Y���Kҍ)3�Y�w� �&�7��ec %sv�ԯv�o7D`�;,�Ͷ͍���Rj7Q(�NHjWA�a*!{n�D;�v@4bّ�L^�[c@��Z'bA�����e鐻n�Ȕ��M{��Գ�[UM�б��N��p��J�ӄ�+\YB"���ͫٹ�g2�#����:p���֛��1�f-�.+Fs {m�(7p-K4��N�FV�mÍDM�.�Ś#�`H�y��TS,O�n)j��b[������[Yp�9�n��f���	���GTY����%D
T�.̰�;�c��teB%7{Gufj�w�or����voŶ�hnn*Zre��2Ӡ�:\������{F��j�]����khmҰ�V-�jh�-�ƒ̺�4V^�w&�=�+$��LI��7X�X��ϥ%{#̷X��wR��U��`�9
�;F�;�b��]V\J�<Xޫ�mET��i�2�f��oAEfѕ�7.iz�\�� �Ǎd�Tˈ p��f V�
���wca���ɖ�R�8�z�ʔ�<�Mއ���.��,f�6��jE�0�ݱ����B��")�M"��u����Cl�.R��ة9B5L n��3Mܡ.�h"�9�P<ɐ�p[�bn*j�����qVIU43\�[I�XE�5{Md�Ac�n��bQ=M[ѕ֜e���[�$[E+s�槰f��Z��v�8Ijx(�$dq��V��r�lp���n;C&�hA{��TA˕v5���Jl����WEiհ�*\�Q�4	8�$Bm�LXԫ!lָc�J���n=jZ�֕i�[�h8�.��&��56���v+2����āB=
Gjd�Ц�ͺ��n�MwwX�7��e[ڿ�L�ѣ[0D2��۪;w4"a�x[v�I�NT:6��v������9��e��LRf�+���M�5B-$Л�!�X��3��v�Q��N��9��v<{��z%�u�;�l�Y��4�wY�LF�Ɇ��@��9n9����R�ێfT�[9��AJͨ$djn9��+Ս꼳�.��i�i�d�ݐ��P�[�W�0���j�m)�W�0"1٪ݩzR��F��n���N� �X�ߗ-g,��n��[`�Y1ɧ�V�����X��95kR�=َ�:*�O�u���/���T��.�����������N鿊�1��h�s�L)���j�>P�u���z2�E�Dա�����חz�%Ӧ,*l������ Ej���&�k�"ȫޒ�Zi�N����vK�^3��J՚ʐ̥m�6��t#V��	�6�l	OZ|�$�em��9^��y�u����y�͙��v[���C݃d[K[�x����U�,j���s͸����K��`����ͭ/�
mK�dt��-��懱=A���Ǌ�l�HaVu<�F��:�"�
˥���ǅ\Ca�n����k�!���m�6��t
��m��i�[�YcZ�A��|�т͸T	�)fE
�\�i�U�M��".�	�\WhDͿ�i��CS�@e$�j���Ո���5��A�zV�jq]�v�����h^H2fq��/.Ȭ�L�lV��C�n�k{	9��,��9�j�����3*�x��@l�P∱��pn1(Qe�)��j�n�n����B�|�\�A��+���Q�x4�c�����e�x�B!�{c35��8hH�	j
*�;e��3/k��oj��vh=�̷h����a�وn���.�nV�4�ӧ4U���U�N�M��5�Vn��0�Z�h�Y1���H�ͤů�����FIn��	�`�K0c;K	�H��K�ʫݎT�R�N�+V=#C�T����&R�+U��%h�M�y�v5���t�L	 ����Tw\ǐ��,���/Kǂ�E,9÷��*����ܤѭTA��O��J���g3,C�C0^9J�nò�$ސՒr�IT�94RS�.�fK��3�X�*�A8�Y�!��D�yomHI��c���`-�^�"
����:��6���x�#�f��26�fVM�����W�j����`�[�%��U�R�A�5��Q�r�^��5�������n�`b^m�x�,&����h��w��Ix�1�"nDIxd5fq�I�%�n�ۂ����h��JU3H�J��р�ۡ�'r�ݔ�y��*A��j�v!W2(]��Y%r�Uyl�Ǖ[{����/�7,dB�cm%(R҃�݄tm�����n�T�G%L�ԑc����Bv�-U5��[dI�V�Q%iR0�Q�0S ��ɔ�������bIW��@�Q�N�L�N�nf���4�hӖmYnKۙ:�;2�R�����h��E4��b�j�̶�w��٫+q=��s*޻ݴY���؉`v�َd:u�����Y�����p:"b7�4I�{�r���*�A�[�iXy�f�c"1�w.�1A�v���I��e ��*��l���&�(f9DU�Kih372�ͽ��ۼMBj�JF�HꜺK�n[��c5�L��M���G;W�3Uw�WTqc�ͲSg0=����V�+ս˲�V;����ׅ��v��c�u�5���Ф(���h0�e����9�0i:dW�&�N4s�[]9�.�%��*�J��n��Axi�[j��Vum�.�Ao9�x�`����V��KV������5�VE�R:�qA���V�ܳX���)fV���ʪa���2��CQB�-[B��$��L�y��:��	��FK��[��&����o]ҡ��wibb��9*M,�ճF�b[�)���6��IT�1M�aMd�WY�\�O����Cj�[�o&�y0���y
�rp��tf�5�]� �gu�{�#x�+ۤ6M˷�3V�u����"X�ΎS�K�i�{[(��SB�*B���v�*z��zs.���JC�c�x�6�n����7t�V,QR��/�i��[6ᱵ�����U�yCH�����IQ��uysJҌ��b�&�SoI`�ڳ�����Z-k7��g�kc�̐�2��
�۔4Jq}��n���3q�XZ�(3q���h3u���-��s2��#�4%�V�޷�%�@#�^lx�ڥdr��������vM�n:�f�͗�kS`�1l��y���z�F�*�r�y��T4֊ݍXQQ��n2�
VMp^���t�K&:��2��ӡ�V�ʖ����f�5�5k��jܷ(4���'wr�+z̕)�����R��a F�K�Nj׆��ǆ�7wQ]nѮa��vF)��	�E��R�YA�mE���^�Qmf��q�/v�tb"X(��Y%J�b�c�n�ٕ�����(�TV,-�)��4��Ul�;���X�Ac�&�՚�;�ݷ�������gD��TV��R+s+7V��2j�j^��B��{Nlq�ze�Lb�bQ��oiե4`�����;O�Fh-}O3,6�ʥ+8����m���hڈ�ה��ZNsYv��V�^�:�(U�([3�����q����P�B,To31�)ʼқrc�q&���ԡ��W�B����\�Y�͉�qU,���6X�uS3�5y��34Y��^�t(���w]j��[�ҽ����V���u��8Y{�n9KK���)"���ͽWu7��4lF]͵76�@����*]�捗��H$y�x- �jtsN��Ѕޝ!��GF���n�K2�n}�y�T�4��ci#Kb��y�W���u�	�H�ˆ�]�6��srRKaY<8|m��ψ*�ଷ��:�/P#����1�ʭ�E�Q@�Qi����"�Z4]ܔ���J�������d:��4ܤ�n���j	R�������T�[�5m��&Jx��K�5ɳ.J�9�=�IR�ڂ����Q�iwV��4�EJ:l���u�f�Z�_/���b*
ʖ���š�6���Hk$�4oUB��l���Z�$�-ŉ��ح�l�x�2�$VU�!�&�p�ڽ��"V���s,��AkYx��Smn�5��&Z�qZ�ı2�M���u�UW&��Պ�׹P��GZg8Z+kVR�T��%,��U���n�#l�#f��5�٬*n�T���6�������G^Arh�α��±b?;V�aBY��i�H�{��ۺ���V�+��O&�b�N�9����ӧ�Ƶ����6����bK��v�:+��}�r��[k���H�ηWW1��k�?�u��l&���L�4H ҨGZ�%USB�v^᭣�:�7b�I�Frty��_ҹj�43u�9�e1z���d��sIH�����3��y�;��^-<�A�<���
�R�J�}��	�+i�[*�sxQ�-+��^3qI��+��g�fH�U��CrSۊ�8��6�+D �*��Љu%���m���)��%���׆�֯*a���*�P���0���e4-�E�Y;��yqQ�Hh��9F^(���4S.l���!mՌ�ZK�ݧ�BI{R���#YY��	����²8_�Ft%������/�8�C3T�0y��C�r߮�S�/�n�ƊT�L��]k��\خѭ�(�z,�V!J�|w�؞>���-h�w��[�n'F���Z0�6��л�Q1��qb�	)x���t��(�I��G���ӭ}ᐣ���22.����<4(��ӛt/���Z�)�bXcI@��G�ỂȺ)��%�K ���2o*邜w�1f��5TF['�f����I���՜D�j�1������U&�U���8�44��X-'��h`�B: �!9���(�]��l�����yD�/nT���Ǆ�i֪��
*v�2��̼���YQ~,�KL�/s^SQ� ��z<��ɼ�4.<xɌkj����gM�y0P�z����eEx�pֺK+t`�ըu�wTظ��2;�i�i�;�ʋT��-r�"��js�d��� ��!�6X׊�OV�32m�ݔ6�Ҏ��-���[E��Y�'&^�3wP���/��+KO��j�6���*һ0 ��U%V�T Flà� hj]���ջlQU(�����Q������j��������v�����+�9jU҅P\K�TUΊX��m����Yg��-g��%W)�*U�7k����hխY��� .�ki�G  �]�VU��j�U�U����:��8J]
l��n�K���1�#O��(����}�o#�ݹl�7:�{i�Ӭ�v���}���}�G1��#y�x'd���xϘ��n1��/�ڸ��ȷ���r��ΣB.�Y���C@�X[n�v��xײ<���;n�g���؜G�CŖ�]���^����{)�@)�N�'�8G�S�m�z��ǎ�nt�]�N���I��݇;�.���1�'nN-��]>Nm�uu��������=��p�l>� E$�f��4J�㩨���j�Y��D�ä�Z��;�K�ر	�twd맇�b�q�=��x8p�'��.��v��Y9��N�KC����S���[�`�v5nynی����x��8�yY�v��ݮú9�\�coF��Om���mu�7�Wt;ɖ-m��n����v��N�F@�M1�M%�H�(m4OM�Dr�����"n�ٛ$P)��؏W��p���%��\�+	׶|�Ðy��q�m�v�����'!v�<��{OOJv�(�.*��l�p���ۮTm½�����r<-��6w)n�^[\ksm�yu��j�h�u�<��,Y6���9cy�p�ԗr���\�4�������δs�*���r�#6���׮�����sϸl��[Y2m0�G�:����u�:����V��a}��d��h�|��|��X���� �g��YN��:�0;����>�7.E�2�c����ջ86���啋�;y۰,����b�f��']K��7�r\�kk�Tv�D�(�3k�Z�bݝ��Q�oK6s�W���t�:x87��1� ���˄]h��ΑSs��(3u�h^ܣm��\s�Ǟ0����^Ҧ#���p�L�S�n9�{Y���=;Wnh�ݷ���'�%>x9pF�E��F�#�*�sV��6�v�u�;�^up-�Ei�S�>-fY͋�g�X0Y�FKjF�Q���vds��v7n�TF�e��&����3�?���n=&.6�^
3��a���m�pL��s�yK1�޹�wY����man�/}֕�//t��b�(�S�+�s�'o\� s�NďB��D7m����МrO}�o����hm�Hvb�t��;L�sV�4O:�;l�t#�c��%4���vɑ��b���\���9Ě.T�;`����Ԟ&�{N�O&�Z�E�Q��u�˨�m�1w��Yw��@�Ӻ��D[��$�*�������Yݜ�ku�K�^��nLlnzp[��i�\xLt���:A�^Kl�-ê�2Y4���I�&٪r:K};u�/�	sش���Cy�t��y=&�4۪;��m�Z���x�\�ٓ�s�n�ݸy�Ei"C�-�nsg�	հ(��um�6}=�ϴ
��Ov{\1��k:σOsj�;Wm�]	nm�[�v���xƺާ����y:ȅ������ú��ڽ�5i���1��.�͜<��ۇ�vok+�j����#��l�l�n�^��-���$�U�}�5���D�m�I�s�-��ɒJ�sڦ�v��v��	��^qm�N<"�4�p���q�yy.�����#�dݮ;K]��Ѓgts��7F#�'g�ń�j���u���d�p<n5mg�ۘɮv�nz��n���q���>�o/6�����M���h�\�eV��V����6�1c���W�^��N{-�k$���n��>�����qɵ˹�Lm�tu�g�Ч:�	��v=5��[u+�crr�n6�3�NXs�Tc���.��vٲ�e�J��<�f��'����s���-'H���E� 8Q���k�����d���Y���	Yd'��TgN��[gZ������75�c�{��ݶs�z{ESqѮ���li�� ^κ�1�}�U�j���zpN��x�¥G��X9�(ۧ�w�-�Y�z9���Kc�+��x��-X5�v������]KB��tj\\$�H9�h�=6x7mK�7o�݆�[���ܾ��d��-9;�`9�^��0�T�7K�v��}�i�m��=Uq�ӂ��n]-\Ɍ�ecu��O2{&�6��\�'��)�{�s���<9�����m^:���^]�k6�q�v�@<���\�m=C�u\�uۇ{�<nҤ��n4gk����xV�:f�0:lV���B�N��r�rE�v:�!���s��;�϶���w7\-Ʒ w���]%�1"�Fv��k8׮$���<�<�*�'<�J���Hs�n���vN�a�ő��x�*4Z��i۶��x��H݌��s�\{vv�і��L�������f��wI��;��gv!�7n�),�nٰ�\nw`��bye��7Z����1��}z�6�ޣ�B7D��kQ���$z��":Ƅ�ܘ�{O�;;q���cH���<X.�P�b���3���pkQ�K��ֈ�M���pheK��u�`�dݶ�0�WX����SSN��m��9�D#9w�H\�׍w=��ݺ]����L�>~��
� [��Ɂ6����Zx�:��lx�X�wo;���]��6޳��5�=ez��G¹-���]�W<q�lxNI읭����I�ۭ���0>�F���kg\4mƬ�:�pm9�ɢ;p�v��M��N��blfQٓ�Wi�[�� ,�\�۫0�q(�;0O�n��;c�n.iq�uvN�[x�s��-��`[g;�}v|������Ӽ��]���`A���wv��n�<��7�v7ؾ�sͲḍ<�nw�\zJo<]�2�IA���ݵېS'V�ƛ�rm����e�8nƱ,/Y{�Vz���3�ګv{L����kY���Ts�^7fLV{�,��;�2&�u6#@��Y.ηWBv.ܐX��A���&��sN��F�ڏd�&�;ݱqn�uڳ[s���ta�&IMv�7"��I>#����t�܇d;z�a��6��m��;�>��\)��[T9x�.ԏn�|h���G���{v�D��&&��8���a�{X��%��봓{=�zW��q۵	)�3��<9�;x��;[k������Z�@VNwg���T��S��yp��r{^o7�� ��u�Ã�������k�e;)�[u���.���h y#>�3�6��d�ۮy
NȠ.ܖ���ܫs��9�f�����^9�NmE���r��n�δleK=t��YM��̍��t��TՉ4F�J��֛�M�Ƶi�P=�n�h{h�nr��J�[ۡ�%�V�;h�'�u������/Vӈn��l�ʜ�s�ݭͷ5�Le%����ؖ:0)�f�������&,R�ȁ�e�kjv:S�v�8�ywcm���CvL��������ew���˜����^�4�s���ƞ���;n`:�A��jKg�vЛWg�;vM�"X�]�Asϭ['z��)̀hms�ۏ�����y�!͇��q�3���K��۟!gx�7:��-<������Te��x��\���s�۷��k�x.#r���4�r�&;U����;{^���u�6��2֑/mƺ�U�@ ��G�箴��rr���KZ�9��^�q㎬\畎3s�x�$�ڱɮ]�|�j	�\�N݃��n��m��qG��;6����b=�8�d�wT1��n;b۳��n ��ʼ<$q[�����^k�s��`^V�vz��ܲc���.(?O�N��ͺGf�j�gOk�����X6�}�f�<^Ӥ�f��m���Β{rٸF��D�r3�2��sֺ�ۏ��'���ݏ&���;��uV�cm��s�j�ڸ�SUt�!�#�mc�
�lN��q��['����MΡg�\����ݳ��Ǒ8��Vƶ7=�u�㛫��������M[��ۃccn#�w,[v#��k�7���6ܙ�����wkz�y���c�e�%X���t�Z����Az䓶�����+���oi�S�Y�3[a2\�x糤�����n�����=�n�$�m�9ܜm�M¨ �{h�&ŋ��n���wp�۶N�.{T�N��%�l�UΜ��͓n�z�W�n��6��r�^v�R).�5�n�n��w��ҟ��<u^���n���z㭐b�t���:�i���ӮJ5�z��{>�����9�[���=�[�[�xmb
y���k�Fk�$��hz�^�M�����駷[1�v���Xom��3�Ƕ�%:q��'/h�6��W[9,<��'m�f������k�u/����cf�9�ؑ�ma�y�4;Z�ï���؝{Nl����=���C�[:z��k�*z�Aqv��mζ}��`s�y�0?J��y�׭���&zy눷(�Ʌ��N'%s<�6�L��z�=���+�un�w�=羏`n��o3VS���9:t#Ѷ�g&ZqoV�+v<!�WS۷s��]�Gi�30l�E�q�Ӌ*3��ex�*�m�T��]���"��'nNi��m�sz9�:����C��ٳ=	v�[��[�`�kU;\N"9ݷ;� ���샱�b��z5i����?}۝Y��ܴ�L�C��z�Yd1�q���];&����`�6��( ݞ/c�ݼ�t��љ.�s�s��ֹ�ut�i-����q=h}�!�ۭ�uĹ2og��.^`g��S�����^2�}����qN�u�<\�^P�qu�'�Wg^Ӥn�műp)lkŲ�Y^w>ْ`6)�n�;=����.���/%d��.t�V�������c�wo�7"����gs�s��Sm�s���n,��Z7��lt[�:s�y�G����$r�ٶ��9qɷ��x�m��^��]q;��{Z{m����ǮMҤn��\�.y޳������u[�z���a�;��Z�Ѻ��z�o3��N^8�b�h��T�N<���.�,n��nջ�z�������:m����c����K1,Kf/�*I$�1f\K1$�3,��K5�n�Ch�k��2U*�!K��j�*�VtT���YZ�s=�sۚ���d��yӎ����[:��[P��D	c����n�2�V]Q�ۭ�&#�m���n��6�v�6@+z�2
��0�	�iU�1��1O���	����W6Ӱ6�0�k1;n��Wo<���P�l�.��+�6��2��y秷Ne�<a�v�9��ۭ�P�V��7]9������Npx��Xp�w<��[K��yJ�xD�ѝ��7c�����mn�^����LsK�i�R��ܚ�Ag�s8c�c�
��d���{{e���Œ�Ųv��6HGh��<���S�;�n9�*d��s�9�ݖ;`#�{o%]*v�	�XXۇ�&��Ӑ�˓+�d������&z���マ����&&g��M�a怸�]&}[l�ػ,a�!�Y|WkLFS�8�*A���=�˝n��>��[��4�s��.�ۃQ�AxE�{sI�ѕ�瓷h�qv�hW�=�;���x���:�
rt �6-8�;�q���n7l�N68�=X���Bv�qmڻ��|b�v9���<�p�n�s�ƶ1-��Oh�����&� ��8���h��7�Q�c����K�vvD̶��Y�m�&�8�J�Q:n7�޸#�lr"�;Lw���c�Z6��%��%���	V�l{mĝ�t������6��	>�od9w
�����r"��G\/!���g�������ת�Vgw^�6���c���u�x��%�ޯ8��N9kq�c�kth��;x�j:z4f�{&�c'b�������$�r�tq�m����x<ɩq�We:�v�n��Y���3۷�ۋ����rq�l��㊷ �n���:3�̻����ؼ��׆�nL���m��6m>un��w3�f{b���	� �n��n �/�xkk$�nqׄ0i��6-�nݤ	M�깊m�6���s�5ȕ6Q���y�a�sqɶ۳���A��]LA��fb�����,ĳi%�6��I-�������
�r�bu�T3u���n��;2�my'���U��'�|��=��v�vѮ�8�Q�yn����>,=����o���9��MA8��^Nn��9��ۧ9�x�>l�`���廰��2�Ʒ=M��.z
��p���g��J�6n{b�-���t�W����n�ܛ����El �X��+x��@p�vў�m��9�uk=)��ŘV�N��dB"i�<c��`3�����v�`�9q�Sx��6�P��/�s[g���5?�_99��Вc1����et$�Z���M�k�v�9F{L;ƞ�J�� �6�{}�����qD�)'��^����e���-�d5:�+ق�mԞ�T���
#/#�)3��x���yMs�y[��jl�r���������+���vf��+�y���#��x���6`u,�+�
�Լ����9�Ǽ�B�*��_�J״t4CB�f&�_��S�4���G�6�e�����<�-��2NL�"�Ҟi�O ��q�{u)�.�y���!u_�0�"�B2$�W�lhA6��7�e���!�������T��!sy�a0�i�Њ��?{9m7 S�z���3�B�G�&k�嗡�����������R���; �u[Z
ꋯ"�l ���U~��91K�=e���|��fڳS�,�^F�#k)���� �$������H�
��tR�eg6�p��x1�i��T3+�	oH� ��vH�������t�oE����T:�;���f:�lb�U��;��x86y�:���%Q���%�^��9o ����&�����,��fV�_C��ϬU<������ؠ1c�8�&Ґ�S����Qʡv��fx�Fׂ+އF�4G�həC2������uM�[5v;36r�S8��9!�"�Epy��/n��x�җ��h�U�N�r�Q%�ڙ�s.��ݮ��T,�Kω�E:/7eƣ�LY��҂f������E�3p5B�����gY1�r��u��/���y?sE��NCg��MB�����-G֞mi�I�0vU
�D��S�a�<��'4v�y�SY��Q[�b�Z���;I7��;P���j�ӫ�N�����J�GsddU�mF�����=�=�����=f��R�^�i0� �
2Z�����/�`=�B�;��p<+q�A"��9�*��;<�`8���Z��1{r���z��r�K#�4�)��v�Nvt�Q��V1�i�Ｆ���b�n��XY#z�TR���:h�%����fV����V����5�嘯k�Gַmj���i!I^VtU������!�o0u�I<��iSX��v�*�T^: h)	08Iȝ���A�_m�d����}��e�ӬHJ�/����2V]v�X<�����VA��"}!��o}/{H�Q�-D�b3A�ԋ#l�����v���R�>"h�����g��������p����ע>*^b��#��l�i-�g�ʮ�E�~����w^��g�vɱu�9=���m��ciWM���h�Hy�X<F5қ�7kB�ޜǔ��Q���Rf��Fu�uf=��j��:aF�s��/q]�L�:�<r4_0FaN?w;;�RT�#�}g�[9�8�q�ջ^��h$��	�;ћ���
G�V��0>׾��M$	�K����ܺ�pz/<�n�H�C��,d���
�&c�j���<��bS"�{J������)8�n�
�/G�=C�)z��W��]v��3��A�cws������EdJw�zwh��v]�j�3l(6iF�5���U���I����y��А��=rM�F3�&e���.���iH�Ǉ
��vRɛ�2.Y��-����2.���lX���1$)Hj��>�t�/6F��ذ[QX��l"��О�t`q�S�u��%G���5.D2�mW
�~�^'v�`���u�NN���u��v��f3���:��4��X���Gj1�2X)0B��������j��,l��e.$���X�J���,;"��R��6�Ӎ�!K�jv���le{Ϊ��(�0HcFH}�q�u��SH݄����	б�D�5;s�T���:��Oa���+/vs��R{���-�s���ۼ��sj�&A e�p��s��U�f|��]ZV���J����>ս�ߑ�8n���Ma:ʳtWgc�~n�*�����aq0ܑ�g+#�S���-�-,�ɬ�+�w��x��j`H��3�y���VB2��>���y��G��/(Px@J!I!���^����B��Ek��C>@�Ӣ�:����5'�	5k�y�Dq��n ,�,���K\D�Z�=�ï������xݧ]\�K���[���Ы�����ٺ/`��{9L��N�3��{�9��G��ް�C�I�J��������Ͷݳ��μ�jգ{]nvッ�G9�ݎ��q���f����}gQ��E���[�Ϭ�o�kmk!9]����qD�02T�thPC���"!����4�Z�㶎X���vŢi�qs���[�mvѮ�f����\��u�n��B��M��8��\��-�*M��W��mb�qk��z
9���!�틣%t>B�\��x4=8zɬv���y���ڛ<�<m�\.���v�\���e�Tl��n�a���G������ץ7�@�;�]a�D�������K ����fj��J����}f��a��	Y� �6p$�U�a�����H+���L�c�V��gX�9�#4�.'Wl�G��5�&�ۓ)ʚ���{X&XUs��B���8��-ʌ�u���N{Y���c���'3s.����.7�)n��<�_M�Ns
�����6�l��Q�d�����8���J����)]'l�śG.�VF_:L�v;B�q\���SljQ�NKL�"hEm��[�d���^Z��d�>씯�{�c+FZ��u��w_�o��}�]�e�gz�u��t�6�J[�|��ډ���]m&[k)T266Kƺ9��p<�}��qq�bB!���`N+�x	��c٥�[>��z��0��p�4;Gdبpb]��n������hΎS�~';qA���Z����J�"%�W�o;Hx��;]�*���^V�GX�
�ɷ��U�v,����;bb��G�8���6��YÆ:�!�{�(7/M�R���+p^CUf�׬m��r(n>��,ˡ�����X�@�;�D�"�2gQ�C�Vt�U�ť���0B����b*�_s�fu՚ݢН|�d�@�9�.)�i��r�U�,�2$W����ւ�zP�fH�
0Te�UE�Y�zMU-x�I�g&5uUfY�\�2)�Pi�Q:��/Wi���k��9nY�梓ov���'@�8���-8�����wX8���ȲV!��w��4�U���v�rڙ\�s/qZ�gB�[yMv�3&�N�D�.�G#zd��b�4�L�w�F1�J{z�<(F�bn:]�8vϜ�����9!��	�ˁ9
ǻ�]�nB����R�S��g��o��ۚ��0���ވ�g<��
n������X.��aT���c���&���}��sհmB��}����BS�ݮͼ�Y̧x�|j��e�o��ig�=t=��/	��b�$��x ���7
H���^C����N���Ws��ZR�W����R'�[��λ*��_S��}H�cv�"5�2����;�c�-�k�=�i!w���,�g޼xծ0�эd�{=�-��)���ZX�P�uto��W���8�A��o�U�}�wc��v1i��1E��S|m\V�_�C�	m��R�[K�rݤ�.бn�jp�XQ�Dш�P��n<�TẨv��� �$����%�(���o����q��y�r�����Drv
|Z�]H�Cށ�r��4b��
 ���$��-$V����.�:�b���*��v���v�)K��	�#.Iys��'e���-��T�@��n�}ǒWحڭ�{g\%�í�Z���L�l�%ֶ�na��"�Tf�qеn����U��j��׊m[�N�7&M��rI��Bˍ����Ťf6�T�w����q٘B@�5����h$8���������c2�<YM����f	�s�/'��!Nٕb*��������c�Q"L��(����p�˲��/m_p�/KzW��ĵ�wwUf��F,�L5�LQ��m�����/��<n]e��Į�62�yA�q��J3���W
rVR�ۭ�oBƞ�R�5��.��)ς;�l�u�7��S�!�X�s�\#��Ϯ��jz|�|�vP@�,���
Ob����Z�n�G֞-;�	���i��˅m��{(���R�����zg�&�f[}�T�]h��d̻�=���]�b�%��vs�q�ٺ;��V��#��n�8$�)�:��&�S�����9�'a�8�Bb�����yu�X���"w3U��sx,���+o<�o�[�R(�Ć'�Vd	o����g+�W�"ko���Ul.�OrZ�����l+�ʮԻ�j�݋;�����л7���4�F�1��0���F�X�
���_�Sxt�x�+n��f�m��T�����aa~e�}Xfx�v���'e_z�z@c�SF���L\�U-Q���*�c����Y��Nz���H[adt�a�)g]ș��r�[�S�ρG6�W3���O�*�BJN%XZf�Pz�{�󾊣�`./llOD�#Թj�ݾ�w�ܢ�(�e�Գ4�O���{E��D�hR��=.8�MO)��(p ��{^Wغ�$u��'hf�y�e���S|�;�S�k��3s�l��g��szZ��A!/�ܻ=�g�f�]looY��M	��7]3d����>{3/gj�v��,�îV��də�&���O�_MN�ʗn��Ƭ�B3h�ݚ;�';�N����[���oG7n�k�6�Յ�ϫ�Q�:�=��Y��繝��ց8��qy5��oS���67n��N˂�����I�\��Y��Ӎ��ܵ�l��˭�gO���������>~��4mofѹ�x�8N�r��l�ps�;<¯]���-+�p7-�8���;��_:��������yc�2d�t&Dr��IUVݻ��
��֧�f�{�M��n���T�c$����C�������]5{�c��l�wۃ.�S&�k	0��V²��M�E�6���g�'�����j#g>���?6��cAO��	)'!j@�=�§o&nzo�7��7�_����;	�>g(th�7�mM�=W½Qw!.�����jb�X���ih�&8�Q�w�{�2���ȬO4�������ͥ����hL��g�Y~̠�r:�k��n���64/ov�Q�p+YC�m����R�R6��Sz�jQl�f��wo���2�\��[�t�����g��Ǥ��q�����a/I	�zw<�[=���-�v�zZp\7�i�JG��4q⠻z��r�Y0�
�Vd�������ͣ���)�N�
r�D�i��K��q�Œ�:�<P|��R��H�RO���BjDc�)$���+�Q��I��a����ڿegi٦�Gq	I��e�3��s���˝v��!��Ԩ���dα\�P�HT,U����r�e�X;o��
�ɚ{�{���)p#f2�m�ޮ���Djꋃ�����8⥤�n���٧��+1Gg&�r��t�ŗ"�������Dj���޹+o=��K�;��,iڽ��|��F3�H�H�~�Ҽ�J7b�5Y�N��2�Ӏ����k�pP�y�2j�D�'�S
�s�b�s�}{�sF+>��Y9��D�	�j����}�n_�~���ʛ�ԨEVc: nJN�J�M�D�)k���'t�^V��v�_��M�gpZ���[�h�d8ëS���sʁ��S�#tpa��݋l2OX�\/=�Cgv�7���\�h�y��lH��ha����F��(�U���6�F�
�nou��=w�ݺ+%�j��#�`L� �I"�-�M/{�l9ՙ�lh2�Χ�rȸ�Q��۬V�"�ZfQKiVR���P�W���Sc��&��SH�8���{)���Vx���v�oj8@����T�����{P�,�Ŏ[�}%��u��k�t �[㶯��p����N�ݴ���ԥ=[��	��47Nn*�����Gu����A��R9�[�u���U�๳�w�7��N�r�ʻ,����$�c�̅L��a�]��틘�a�R�>:�'%fub�	�#2fʷ|5�<��ޱ�RÑte��Ν�\KgJ�ZC�.`�}���ꖫ}F��_uw��.B���K��"(h��/�5���	�ن��ub���}�0
'vގ�s�� "j���fP����Z9���}}wR�4���򤰥��s3xX��Bn�<�'{v	M"z<�����g��Z��=w���#���w;躻S�1��8���9y�^,�=o�B*ӻi�b�Y�Ŵs�Z�� U�-c���C�LOOi����Wi���n���^�f���m���t�����:�wA��̢�Q�J���oF����}5\;��B�`�ָ�ڄ^���uvhX	�'v=��q���e+�@�/����5�-�@�nY#�:]����r���{5N�.J=Y[{B��CD7ղgoLS�n���`��x6\�E)%ɚ-���\|����{7��8���°ev�m��
��X�pk՘�q V�9l�d��ᷬmv��q;����2�7�Dq_Ex��WU�M�X��KY�U���.��ܫͲ�� I�J����m�RY��R�6��p����lU�����"�;tS�$�y�����:A$��}�Xx� 3ֺF� t��y��>" x������J����~s��F��,���+���V�T����"r���6:�:C��<]�0�o�~U�V��Y�G�{�?�{��$0E�d��
"���[ߜ�����(�7/�t����d|�(�<І����u�!ML9!�y��l�@� ag���|��A0���o�H�Gq�%���|�ÿ����g�$@���:`\�Y�QY��B��ydo�_ƄhC���i�+lCΐ�ٖ�ښm[9ԭ'��n3�3)Pb<\�,�]����Gnc��Kͻh�!1GGlh--Q�I,�.=4��̚Xt��������H��+�x\E�>]�+т(y?�P��1���o��}<˓GL�@�]�'��F�<�!)�����4�].x������i=m���b�Ku�������6��?|����0�]�h~}�HWyG���C!�b2�X�C֣��y����P{��}s4�?!0*<^ϲXG�x�vC���Q]�;�y�.�['���K����N��:t�xOU��#�>Uoƹ�i���#�A�B��_]:�����z�T�����\oP_���=E�����a@����ޛj� n(�g�?�0�fQ����Q�8k�<��~��7�y��<Z�λ��x��ظ>�]�NZ��i���h�ju����d�_۴lp����i`sr�y�>�mSK3;D�X񶝝�;I���y�|�Me^��~u2�LX͆�N��5�\1��#�|���]y�"�����Ԇ�Q�~ͭ���6�(壅��(���j��`�ī�ϴ�L�PDQ�/˖x*�>�D�0�o�G_h�|��ΰH�˴ �pw�����WV6�^��Wv#dy�������vy���OϽ��"+|��F��@	/4��&�YN{+u�w�sHY�5�={t��%�$���8�����7���a��k�@QA��j���^��|F`\��y��,��g4�<߽�0��0�_���y�7� ||\���i2byS{R�,��"yDh/q�<dfw9�Z!بӲ����Rx�p\x�����
��;� E��y��(z�-�낳v|@��ӿjcOb�i
ɟJ���"��!��+<��u��:x�(bһ�\N�w����Z�������0 Y�G$7����
>�P@"/�O΢@pјlFG��@�c�S�����_r�P��<�g�ga��Y��Q��07��* Ť�{�zY��YGO�M	�sҝ�ȣ�dB8����1�	Mɀa�\Jأ������n��!�Ŝ��]p}�u�x;nH@f���r�p}x�!��'�����+�#H��x�. <��+$T�]Y�<������PV����cГ���T��K7��_��?�-�_�x�A{_���QQ|C4_f@ǰET��j��/�E�A�a9�>k�eu �w*���ϏN�؈��@eJ�.��΃#N�x���44���7�k��o���]�+��U�;�U�eee�W}C9/�8,E.d�Q����o;0�]v�yՔ��'��N����z��|����N� 9$�(����r��l�n�v�΢|�/i�K�x�u�Z�<viX�]d�\�����b8��ґO���m�r�rN�v�[12�K��N5��B�����I�p��]n��p�2XK!mb�6w�/ ��Z:%q��}�.�t���8v��<��;��>�r� sf�I�6�ήܯN��:�e��H�8��c7�r4=�W'�\�@!���G;l����m��0m���`��+f��ι�l�p��p~��"��}ߘx6���|GԹ<��G�{�t���H�B�!jzEG��x�ծ�o���dw}ƹ�~�zz���,�����;w��"�WW��Q��6����o�ϫ�"�!%fHs�O(�FBK<'�ۧk��������ޥc���Ϣ��}��B����4��G��Ї�� :�k��*A(��c���f4��C���qC�x+.�+.�ו���W4�w���jbl��c- K,�\��gZ��J�qѲ��Η�|��xyyG��]N
#/��*�W��^��+���Lwo���ޔV�]Zp�G<�MG�h���W�w��4��e.A<��%��N&�@�䌧%�ȼ\�
���'��G`wW��� �>] /�(�<��c�����`'��LE�����+�D�~#�,�|����\^Lw/t�=��Ћ>�� i��>��<�(�Gϻ��I:H��K�j�-����үc�{W]�ʉ�#�s�L�w�U�E���+���ߏ�K��@e����r��ϥ����f�;5�	���@x��߾tj獞� ^U࠺���3Ny�D�g���{�ڪ��xzU��4[J�rج�T�Z����p����yv�I\�xt)8���k��d��C�t�ψd8�S%�O�{�C�a'�Є#��|C��e�j��B>��F � #̺�QU�u�9Y-��y�D���`"�,���x�%��N~�qW�����߃��Z���
.G@#����;�H��/1�}Wߝso���w�y>	E�\Y�u�e�s{�`��U#4�1�8�b]:�۸�j�dq2�T�Nj�6�-���o�s7_D:)�su9����25�5�Y��!	k�D"��q^]����G�"�pB��ق��R�������a'����tь:p�Im���;������h{�g�Gl���JdBR
P5#�<���\B<$
���Ur�`�?/d�O���F��}��*4{8�${so������6�1�51��W�r�Y�ײ�0�:��E�TEI�}(|~'������Y��y��^��!"R5�+�G�><]Pٲ�,Y���g��aΎ��|�}�(B<t锾!
 2ȇ�AX�u�!Ǥ
<(���]��S����G���#�}���e�B��;G�W_�}��1�c��t������ThD�n����!��CФ�<���ߕF�8�G݇w����������6���~�|�H�!��/
#)V.<��ԣ���b�ٍy���QCЍlW$����|�5�ɲxk�1�-���<-������X�q՝���ݜqkDM���@gڰ��Y�!�<���ջ���0���G��_�=hQ�Sߕ ϗ�8({F	(ty=��\T�i��v�e[�,�<��!Y��ý��.x�:g�W�����?V>�u�Z6�`YdN;��:xȇ��1 Rm]��(�������d�|�(��qn�rc���X�><�q�w:��	�"��~U>� ��b�;γ��|E��X�p؁F�E����<`"�
f"��ǰE�VV|+�xc��g�fx��Z#��}����J�[�������"ň�f�
�I�����!W��J�tC����{Q��q�r�#x��s�u��#5�Tk���j�p۫.��B>z��h,��!�yG�DY���V�N!y�x>�g����2`�7�n�RVh�
G\��Ju��������*�v㗰z>�ُ��th1�5G�}�x�Mr��J�� :v�ӹy�Cʞ;ߕ���,�P�4��v�(��x5���NAd��w�Z��{��DYz�g����8@����9���c��j�p���N��	���B5��tF���ä&���@���u*,�5��H�B	���~�R��C����h"�R1-8㎪;����ۮ��cP��h]��D��Щ�Vh�B�i��~��!�{u�Py�V��F	�}��~�}��`�0Ǻ�Ү> 2���\T�p��o�Q�>��A����DB{�C�D�>U(�_��z�(�x>��I3:��b5�,�����G���zH!x���W #H^ߺ�?wu����"g_;y޺�������C�"������D�H� �^�>#OӺ��o�c����� ��!y�70����^3@��Tm�2TK^�6�}�z-����J� >��]pa�� }�]W�M|��}�^�yn���{��Ū�%�X�i��C�;��QG��@z��l��#�{���4~=<-�Cͯ����^d0������䎸,��0H��ڥY��~�a<��<aG�ۿT�"%̋�#]����"*�:Gj�Us����sP�?^�UQ�gβo�8h�H��c��˩v��3IKO�'�ig;W��ۤ��+��M��
1��i6�\�.���kpf���%^���,6fM��T�v�:Y�-J�Q�]��P��#���� Y��cXh�"!���%pf(/�OH���OH�B0����4I�!�h�[f�����Ȕo�T	�i�Gݿ@��u,<�j|���Q����`wW�@yl�t�����=h���SŽ��@~��SC�Tq�F8F���M۱�7\=cq�8�sq��3��	�玨^5v���l��BJw���*G����Z���4�{��E\�x�k��t�g��\V�4�A�G�>�0�!��k�o1�9��!��i#�<Ӈ-pU�l�Ǧ��W�y���G��B�����BE"���GMD�Y�4�d|G~N�R�(cϓ'��xv�E�Yj�c�i�ט�]��ɏ����������G�P�D��C�u�U��#G���ojMz(xs����4�@!�!)��o�N���kN�hI�����C���:l��iG�.*,��Ľ�x�pu�\���̽(��z(��U���{�>r����j���C��x=�f+ߟ�\�z��|�D�h�ZF�Q�$�"έ�	�?'�g}�d�f���2b�#����f�dC/�|���� G�y��!�Gb����*�r�8y}B�4� p�{�������-���'��4E�:ϋ�~ٶ���۱� �!��Mb�θ�<�(�d`�Z��ʉ�z���t2��V4;�Z��Q�̙�!���\�|~��!�:���+��:h�D�HD$��~�_f<�da(��)p��<?���V�z��r�6�P`��W)�/c�Y��	o��-�Va{cA[��0��>�1 ���4��D��w�a[�xI]�mm���Y2mZʹ��&.���!q�Ŏ�(M�d�ۇ��]��z���l�Ӡ�y��ϖ�;�up]��e����ٝ����^1ӍE��=vm�^w��qG[�����>w���۲��C�on8�ڇ����&�]��nݷu��L���τ��O=]�ʨdů ���ӧ٘-�)�<Zeܝ\��v�g��.t�]�)ucZ&z�`Fgt�p��p��n�َ�Y-uҋ�n]�@��mu`�Z���ڳv�E��!�E�DC����腞Y�@���o�~v:Gڹ�[�V�*!g��rȮ�9y�,�V_Ƽ��<�p{���T��#��?!�K���b��0�C��V���#��'LD5qQGRH�>6adv�il�3���g�G����ë�X+����I�#�ܺ5����p����ψ6��R��<���(T�}�!"A�W��@����g��yj�4�����E���TH�Um�YY%7���\Zx��a�:|h�}��T6h�!e�@a�XB��ʾ i�fȰ��{�bszb�ӿ.{T��t���� {�yi#���X6�P�������H�r�0�*>$.�A�ۏ �O4�h�8�W�)���r�u~�$��]���wel�~�ú1�WU\2�|�a���f���<GM�0�����xF�����8�,H��NQ��z�˫tB<�Ta���Scqa'��/�����Q�"L�x4�A<����� A�b��H�,�i|�pQ߳��w샬�z��0� Ȇ�D^+<{x��u�v0�2�Q��lՃů��ƕy��e��gɨ�����TO�ڵ`����!m��5��ˮ8�	X�sl�؝��R���fZ���:6IS�*�!)�_<��������N#�k���iC��@�+S��l�yX��@i��Ȇ�����/�cH}����s�d���m&��h��� (�4Q�Ϫ�������bpQ毘�^=$��D��D�Ɂ��i�C�(�#
0���W�-ڡG�GY.�]"Hh�XF���Z�(;P�!Ԓ�q��$�j����*��5���fd;�v��r�츔z1*��u�������g�D#͞�� j����P�CІQ�,�ƣ�ĥ�@�}�Z�hQ5Ƿw�c�C��>M�p_�?�@7d��c��1z|�'����9�m:���/�m�4��D(�=9���k�Ha"ɤ0�Eς��@������gD�k&<�#�w�E���\4@�L��i:���2��pi�a�4O!��}�4�{e&�\%�	d�!�C\t����MW�%�݈�"8h���[�� ���F��v�ӧ����\
w# Q�V�#��,��pۯ� M� 3���d����������W���C0���U6@��kc���|��P���Ki�����~^�x0�#��U�,:D��Oqr���z(h��T���|��~��j���;�aY�B5�F6�yV0�ڍ˴�a��.��tv������",���z�>�>��#	Lj��A"�<�D�L`�$����.���m��
�"ެT!n2尬���ض�5���W�J?�r_U��nJ��I�>��@�VI'M�����i���<��� <��d�����2!F�/�`�3�Y}H��ܡ����<A>��1p3�ܔ˩�CE&L6��8ydC���7hN��~����&��aV�Le:x-����7��5�<��vKQB40E�`�����t��H�<����|�#�|m��جwzD'�/k�. �/�|B�AJ[e|m.5�[ꇊ���\­1K�|�4�Y����2-��̻��|@���(��Aג�����2�3�)u�u�t�	ĺV���?=޵E�3r�]K;�	y��"�}��3����/mp17�b�ͯK�߮�ұtyO�#D7<ED����G�a��8G�_#�Bl�ٺ�:���)�r"8H�{��Cp��#��>���#�����ψ�k��v�(�x�|�e ��`�.a�6oԢ;�tk�|�iϣ  ������9һ�O�~�ɼ���@��<�Y��(�#�h�˻jB�`�T����!�i�yGևH���ݷB�;�g谋��٬o�,���?}���m��yg0�b��Q�!� U}�:�$Y���#��}ht�++��Y1�GO��x;����s�^�jݵ6�J�+y����sͷ�X���8���ظ��Z,�qJ����r�m�C�<�76|��<�BȲ<p����\E"f�&�|)}�E�E��^�#��+�Ɉ��@|;�+r_��y�}j�O�<���G�<l�y���4��l֢t��\�������3����d��-{ŷ�k�z$}�H��um� I���^iD{'�&���}�3�!��W���c���� m*!� ϭY1}�d�vP֞gO1�P��g
���!g[�}��p<��|�b�kی����#%rKi�4�E�oun���>�<�b����\j�;���>y���75�Qdk�#X7������G�f^�>��t��Z���:G�7�4���	�3��A�=[z�G��V8GU��	oqw�t|{y_��n����OM�x��}+�4�r��	�Wk�����s�q���#���b��LT0a�= m ��]������JŜu��v���%�0�5�]�V����7����\C�n=8��^]��ƞM�q������R��b�|(ilz�sPY���p�������	>Bΐ+��h�	�dnJ�#;�1d6ko�	���i��Q�<߂�Q�yߐ6��|���UyW�y�>����]�V���%2�u�#�<a��ǹ�m�y���@3T?(��T�ԣ��oϢ��iЀ�NܤWts�="�u���O=k;>u.�oiь,�YhD�HW#����j���Z<~hB;�����j�%�]�dY����,������,�[]hY��Y���-z���g�}]��'�K�,�\�-q�/Ɔ��t�<��%��˃��uFF����^hwlM��G�I�����Nʵ�%63���x>]�� ��\��j�QD?(���3��@}�h�a��R�<���w��N�i*�����~�M�|E�_��E ��dx&d �Y1�$�/�ö���t��&��y��Xb4z$!�|�J$v��?
���_�!�2Hg������pڧ�Gԑ���|���>:@�F�8x�<��Q���i_��Ϣ���In7��2'$�!�dx5�d#�~�a�����a��
�C͟�-�!�}�(��5������F �ӂi��
5�]>��~*��y���E����~(��Gǘ�6Wudi��#�!=ό;�i� ���׭�%ǝ��ʹh�mf���Հ��!�G��\�����w�D������G��B�+���J��:x�3[����}����?k��ia�0�9������t����Wޗ�6a�ye�1ԅt�3�C[kA.	6����+�����+���ۙ	�F�sb	���6�c��#��ԊM�Y�snڤ�ŗ�H��TA�x����x8��R�ث.���������3M�0\�X�f�&X���ܬ�đw�w�����D3�+�`bHɤ��>�\2b�߭�c��v�r��OcyWN��!���[��*���R��>� ]�S9\�8ގvw�6;����K呀�/���_��V��ghn�|:쮴K}{7.^����}�qcm��V�f�g6J����Z�\xoX���C��Y7��ޕ}�A����o>R=޴wv���Ȧ4̦�U��8���oQ�ηY����	;(tkF��5�uX3�N��^7O� �Q��T���(���^�ogX!Un�g����tupRt!������+�w+�W,�z^�w�Y����v�D�3�!O4�[���a��r���v����f8��5k���
�̓�&�;�;�]X4��ӻ�]�oj�F��+ba�U�Ì���Tְ:>٧&�Wڤ�J�Y���r�vwÐ��[����Q��gȌ66�� ��X�',�0[�y��'��n9e,n��:ɽ���s!��[9�|[��Yf�F#��,��kIG�����Y$���a4a{�!߯*�"��!����@�>=Y�b��ܿ��@tH}pu���n����ӕ��(vVc-U��o {���՗��1�e�+l q�]��A�g�$�\ 'Fs�E͎���%V����V���x:C�P�:9^���|c�YÝ���傌5+��<�U[��^�T;��W5e�1�f�xv��s�� �6�2F�9�C�
�/ZY�u���vˁ��
��)�,�s��낥%�x��������a�t9�+w�6�8�w��v�M�����������۞t���L�;n�חqltb�`�yǴ���4��Q�۷<a���@=�ra��ݳ^�mv6��ٷm�~�v���nÏ?&Z��(krn�Wv���V�����F��7nx�H���n��Q��4���sJnxOَ���u 3h�q�*��yC����V�&�����n�js��g�s۱��=&�i%��3���"�*v�mn���Oc�I��p�5e3�ݭvadi�;;�cq��n��Tqe�tm�<��v6Axv8�y�	=�4�[���M;n�ݽ�������hX��nض�.�r�έ>,m˟Z�,��V���i�mq�z����<d�\�'+����5��r;F;�|ux�v�zm�}����u6A%s�JkknhЉi�qO3�8b��������x�����:5`���z�6w���[��X���b��k�tX�u�U���v�ǈ�L��'Nc�QY�ʭ���T�������p��y�3�m�=�������bP5�B'�K�n���ۀ�������T�>���v�c.L8�	�!�յ���lJo�������s系�M0��9�m�ͱ���qs�h�f8+�Mk��7n�u76z��cv�i%,g�3\[�����M�ojqn��U��:�w9���7ok�f㞤�vk�|v�d�ם�&�ۮ�����\�m]*���ݝ���f��:8˳���r�u`�5�7�5��Ǯ�
�����']�b8�O���e�k����^�%��`L���Eۋ�k9۲盵[�oQ�g���\w�;n�몮�ڃ�g���sۛ����9��<����	��=%�gx�ݏ ��nr���=p��P.��.��z�k2�2��m�Nkv�����I�7m������nYUk�};BM"t��p������u(�I�G����Kv[�㴶���s��#�뷌�s� gt��fn#p�n3ǐ��j�V��ػX\+:s��$���y\��X�=g��B{m�4�L<`�o6m�n�kE�ngf�m��on�;Z���L�����ܱ��W����Hg�O-<-������Y�*���do:�V4�Q��O|iv�E����0�C�� �3M�~��?Lfݧ�m��u�#�>8B<�"<r����t;�+�,�@3���Q�>܃�p|.�2���8��WO(�����(�F�hp�"5�Vqѯ` �M�dq���	���3<j� ������2�D�x(����]�<�W�� �@�G���3�>io��~�u^�77�B���[�{i��4��y4�:��	n���}�(X�"��DP�1����Ĉ�����=.�U��
,�&�>��ا��<�����r-�!�A���}��e��	��J�� gU�@a�j�_��~�(��B�Y^�q��B4zF�Es?e�"��ߣw��G��ϵ�Y�1ad޺d��Y��񖹤H�=_g�r��\D�w�����P���4���C�!��!�(^kO-�j�:�x~���*��!�%�ߩ���.�|��C���Т��7�`#�u.C�v��xC];���}2��E�=�r��K��F#����a�3r~��Dt2G��� ���E�,zOf�@h�H�AHG����o�|ޏMqpd}��,Q�(�RV�wh���Y�a��c�i��L==cpꋶBђ�����y�B�(�K����Y�:C8F�����y�O��t���k$B�B���h�G����TV�zy�8��(<���$t�'�Y�4y�4f��?5)�|~_5���쐴B�����!��E��$�C9'Nw�Eb1!���[�S_,��*�շ�1B�0YD�FlW;V��E�ҥJ�
��^2PLj���c���ݎ��8�Y��xv��j]W��S�鋗~��B.��<�-5"���+�0�z�ȇ��b�=tO��t:x+rx�#��v�7�o��6Iz�<�{x��j�t���1��m���_�k͕��F�㌩!����d��H��Y2eg֫���a�~�,���\�gղ�N�]LDP���P��#aC4hLɺ�V>$�������(���w����}�@|p��B���#�4�NZÆ�	�_QAd�& M�drIB�Iy��G�M��+����۹��$Cό5�Ӳ��a�~�,����
���t�����Mj�R���_|�B=���E�D��d_<e�|�� t^��B�u��|@e�<�}�ꌱ!	C"p��aGƁx!�G��ﾻ4�#���u]A��F��o�)��/k:���E�!���ȇ������ʀ���谁�/GDQ�33�a')i
�o���3R"�hY�g�D޿�3�`[�*���r[��1���'��^���p㑍�����Q�u1�nӏRv�߷w氲(�B�"���N�A8F�C��S<�/�'���Q ��t�<���������f����o@c�p�0�|�x~��P��"�U1��OL��!�F����[YKM���^k�O,�ȅ�)���v<�>����S�h��4�E��F��D�����Qdw�n!ms�ْ�T���
^@�y�;�����|6��?S��K]�ȸ#O�.�|��p$��q�A�����4��G�h��}���5�P!� Ra������qc� "	-q�s2�=���vi�鱥��˭�Y�0�]@◳0f�޼�V4�^�SK9%+����a�&r�$�w�w;�Km�E��l�h��z 8=������G�w�ǵ GK CIQ �<�C5��<��}N������\��.�b�RH�	u�~}x���,��߷㣠A�d���di���V}t ���;�\��_<�,"g��KON�$u��+���:y�W�$#��)��o�\��$t�<o �.�!8G��q�����MI9\J5
�P�9*1@�D��E�}�C=~O'4h��E�"E�h�[��Mo�F���vW��s�>�!�A5��gxy�ݪ�HgA���4G��I~��	������3PDQ�,���A��ж���R�NI�]��Gj�S�\l�5�݇���,,j� E�c��%�[�ߛ���0��Q�?Zu�,�{��\�<�Dw�.�t@����;!}����xx�g�:FҙLa����;�{{��E&z��p���c���D|E%�/�Cqt�H�h�H�!Ww�{��q6drIzp��A��"�ϫ���w�߈Gk����J�9�\�H����s{(x����r(��	��G��g�U��E!F�����fJ=h<�>��(B,g��!�wW,�DQ竽����FQ�@c�8y���p�Y�ĝ�$Q;�}(i����ȇH:-�QK�쿾W���cV����[�n��<~�����j��=#H��udY���=���	yd�FD�5�ՠ[k�#���,Q��uR\�Ց�P�c��ب�᫫|��j�����kK=!x2���B��ϳ��֋1�(C�D1�f#_�����"ò[^�`�z�s�h}5�Y�Tͪ�|�g�a�������*N뷧c]|;̝ӻ�_tO4R�F����7M�0q{��h��ɥ<y!7�08u����=����N���s��r�f<'k$��Z�!+r��K���Β��F�k��D6V(Eo>Ug��B�X���V�>Av��#fw��^����d��F�!+|����MqZe 0Q'���5���<����E�dӄ^x�~ύ߾��N���h8��\�j��V;;�5E�W%����Q��P��v1=z�!�4��>#�1��D2A�}!g�]oθ;��ȣ��HU�I诳�^�=H�x¢$�P����)�L�w��|��8D?8����͟+��v���#v���d�����ƍ���q&-�b�uGش��l�"�X������+���EhK'q��4�g�#o��x${E�{�
�}c�Q�0�8�6@��2%}_JG��}=#�qy�g�n���^w��hU;"6�qn�o �(B��Bw�ʆ�r���7��2}ɧ_���$Y�3��߳E㺆���!#��%'��F��{�X� p������K�=�{�u b�����d���{�,�e�2��y�����4��YG�����==�I���
I�$pV1k�;����ʺƾ�_}��J#�ʝt6Fy"(�m!���G����,� "�x��qa`�=_{�L؇V�DR84D��#��-�΋��YW�s���A|�E�wߠZ�'�vNux��R8R�f�mu��{��T1G�i7��@Jۻ�k���PG�����X"�#�}���������B�~`h8t�(���	�_j�L����>�@�����$�8y�5{o���_/K˿AH���3�]Ce!��Ti��F�`���l78ݛ��*�4H�*�������`쥡���$����*�c�δ<�F80���=�ˠ\�|�\cj��;��JPimՉ��]�C����]�ͧat�����1{�N�Yݍ뎲�r�cl�秣^Sͫ4�2:�a�aͦ��p��3���˧wK�I��.��c�Ì�>�(;k�be�6�.�ݝ��]��+���kI����n�3RPi۫=�7<���m��f�� 8������)�ܜ�?�[����'k�R�튝ڋ+���v:��&�{�Ƹ�M� �R�8'VbA�O8K�|���F��(�)�I"R���F�!�#��!()Hn�G���k�G�L�P>6zG��a�h��2kU`�֛_��� ����8��#���A�dn��,#
��[��'����N2Y`����	:~"��4��*a� �:U��{�P��>ྀ;��Z�����F�H�>����O+�2P~�h�#�,�}�O��<�>"Y�:呇�D<�!�B<���𨟏��p�W6�g�~����a�G÷v-	A�l�\�
��D��yU�"{4��/��P��(�\�\��	�7J�>��΀����4Q��,����#��&z���{�+�:y"}"*��)1�q��G�opP��t����ߐ���ɫN�z�Q�5���v���3V�����}�[<��{�u���z�DQ��=�4�q}N�>��O]�=B��\]B�#��ު��0�;f +��|�}7p�9�x=[��3˧�����k�ʴ!��V��
�����K5��?;L��U�&�>a6@�#�e$�����&���B����@��~ϬP�gς�O>&.d(JYH2/'�(a&��ip�&IV!��va�;����:y���?�Y��|xEx�t?���.z��
L[i�al�&�ǄL�=��z�E�kY�u�[3`0g��������T2H���I����<&ϼ���b��m;n2�8E�P�ݵyV�]nٮ}[>t�a�Af�AD�9����0��t,�oC�Ee�h��Q�Ih�HJ\��ޔ,�t�,�Dzq�F���y�y�0���-5�o�8H0 � I�1�@r|����K���p�wȾ�E��ƾ����To��<Tvc��)ᝮ��u^�������ɕ(�*����m��OZ�$�����5:$���t���w���֫�_(c�g˹E�����e��B�~��	<�%�?Q�� t��^���m����m#6�0����>߭��w$��Ad���.�1�M��J�>'��U�l�CǔQ�����F@��>����1�,{"��h���u q,�{���ӧ���".�=&� ���KS�C��q�l�Y�	T�����I�� pƚ�4�!����Hp�G펌��'��,��#�o*��ALX@
"�C�@�`� `(Hg�D0�ҍ��#ٞ�׷M�ǴFX�hb�c���f�*�g�4�A4���x;�b�&���P6ą�$��M�>�@��G����dY����}��[\'�"����/}�y��ޑ^��P���@�.v��|��Y<�VXa�Dh�߳�+�N��$ҳ�&��y_^�|�����7N�(�%#)IdRH2�;�<��⺭�K�Z����v ���.���wP��m�$s�Hf5e�+U�.���|GA�F�}*��L4�$]hIIi$�{�<隹	4y���ʥ��4x����l8���۵�F�#��&X=Kz�!>ϳ����:x>�l���������8~��kP�Z�*!"�!�1�����h��لa��;r��E���#�<>ހ 'Gk��,�[�{��\�h�Qdߠ��d���$�~�4,���Αx��H���}��T^��J<l���미�����x��ǘ��4@�t-?'")Q@㎃!%�	'�e��'�ܖA:@�oq�0�"�aF�p+�#����f��s�"H����cdߗ����!�F���
�Q���<������l���'Q�NRQW<�p.'lզ�`�,�鰊2w�eP[�NX3/N��O�?.��:^M~���Ԉ�{x��<�mY�O���:�t�~(���E���hq���⵩j)
�k&�Ƹ�Br��b���ޕ<e��"�G-����O���:Z5d�}�`G����Z�}(a$�Ϗ_>,��=�V."*��I���P�>%��	<8���r�D����?\��o�$�f����"c�4M�OF7��_�tL�q�c���7����
 �A��� �&z�t0�kܧ��!��c$"�<�c�~v�Wy錄;��sH�ΐ�Y$�\}y����}��\��:��Y;���7��4H�0��!�lM.b�x���G�6���Y�Q$� n�0���g�A7-퐭s&a����z�V֝f�룑�C�����#�x?�:G���G�����B#����B�$Mt�� #{�C�1�	���H��	?+b�.��yS\�^t�<�ϱ�K¬M�,��ҬP�Ȕ�/HN.[D�Ow�c�  �#�̘cF�"c���Z���,�Е9i��O��4���"���7�2� ,֘�pߌ�ۍ4�ѳ��=�_Ɨ)���	��X�#E
�X<3����o�U�Ι`�1BAX�*��}�� ���?B5�~�����D'�ZD�^#Վ���"��-�K��'74�hy�U�B�T���·I#J6�E�"wfV����]$���J����; ~1�7���<)�b�B
�Dsݟ^���`�����]/�B(�IHQ��̔+�i�(�x��}XRI�G$m�@X8Q%�'��n�	�Go0&��sQ�H0� U ���s�����K�����Й'��/�a��{Z?3*]���1H�d #�m�F��F_�5(\a~���rg �Amlwe�b����@{mqbΫ�].�UCp�#}��gf�u�N��k�7�m/�R=��x
<�[����#㶡%�A'��n^�ݔdN���%��c\h�&��@C�P����uX)���mÄ>.��(YԆ�gra�������ؙ�tԺ��R6��Z���0���<��>_�fܤ���q<j�p�f�!��|�8B<��Vř�� C�b鯷�:7~���4[AI	0�#�8k��9-��D�����hz��i��$<���\Y	0"���8�M* Οh��k���6. ��	J��˵�l�HՒǼ�W�S>�!ŐE	:�+���܋��?���y�<ɂ0�ŉ�Sh��P �Vkت����B**�i��Ҕ�c�w�N���+\&�NC�<d\\����C{�Q���<�1�}��M<����dz$h� H����PM�5��M�y����������@�kg� � G���>i����wLb0�'�����8b.���^���eV��b(o��$@�h�X�,`�&/�4��/�`3cW ��a�A"��5[��n~�V<ɪ�p��0��������ӓﾋ��IQĸn�uX=!���~@QDQ1Qe�K��0���E{�2��Q���������D�i0D��I&$���[�	<6�<���Rv��b>�������@=�TY��*ЄCU���s؁ǰC�,�8@������o�#M�<4���;@y��l�G�;_̑ |]�M�#�Bp�M����ad��6F��
R��9i�]}�6{����	�|4�#�e_ڮɤ0���H'�bD��wG�g���\>��5���1�V.W�#�ΐ0K����(���B<��>/�u��y��W%���B�0L!���=�W}Vn��k~�P|]�^awR���>�*f�-��
-N�C��lpk��t��Ia5o3�o{pf�P)��G�7�q;�ZE;N!dns��܏g��펬�iz�n���J	��Q�l���&��A�q����v�\lf�[<�k��1��F�3Q�v$�nw��f���;�V�H�s�t=Gr�눱��,���.��%먄���ro5��ኖ���V�K����+m݌��g�Ro\�m�κ$���v1v�i��َs�+t�:�L㳡n/v;�&�'Um֚÷;q�ۛ�;6=r�I�y�9N�\ڷ\̗j�YaK��nm�*}��G�+:�Z���'���I���V �cQ��t>��W� d�}�8;���(�ψ�}�O�^������:'����o>#��(��"� P#����5`�#DB � ���Y�!(jǩ�'AF\�8pp�?}���� {D�hP�w�MK��0`�!���e:�j,Iг9��(��� ��|����8|� *^� I�����M��8C?F	��DC��gƅ�뜝>"�N��.?W�b�i�b,�`� �{��g���)���nL� �PG�M�"��5rx��}ߝ$�(���w���������7��:F1���A�:*{"�p�8z/����cfP�=@o�H��؉
���ر����6p��:��q���@̈6\�������I�(�	�/O�A�C��@;�����Ii�\��
�^ Q�Cp9��x�H�~'�� �* Y�q�)溳����V@v���0D��n�QS� t��U� M�,�	��f�$�\��b�pdϖ���GXKn��cVzu�hi�A����/��c�N	��T��Q����ʌҼހgٓ^�mD�%�dx�#J=6~"��w=j��V��H�ߤ�(��TEbῷ΅��$�㇄T� �5�DU���"}�Ȉ���m��~�n^E{f�#�[6ޔ`;n�v�xnX��y��VR���nk���Uy�ˋs���j��F�D��^�W,�8�<�A-AEs�Ҳ:x}b���A�B����)h�>0��_ά�!���CY��æ��\6[G��OP�׽�b�#H�<l� ���@A���Wkh��V�H�ܶ�n����	���G��!\F��n���P���\ry�����D��#�������VՆ!��ӿ+�n��W7��Ě��Qu�%Ag����-j���4Uur�>v�����$5϶��?���z�Y�\�d{"�r�аl�x�!�"�c)q�X����"%�ԉ$�7�u�#�Z�����\�H�j��<O4�a���>��J,$w��[��mR�n�Zݴ�n3��Z@�P�H�|h���� �F��"ݰ�$�Wh��WڬY%%ݲ�����ǣ*V|���G��E������8¸��*@#K�T�Tzh�׷�C����OP���ifH҆��k�)$iH$f 䎅�F`զ͒yf��O�1u��d� CD�?��H��/W�0�}+��A�UG�w]�n!��F�h��if>3�w�*�H��f�ǶʲD��4���񁃾�υ�T><:�.!!�V�d�bBFT��p�9�Ht��pQ�}_P�P�~1��zW�a(�D(���9Hy}��;�����U�@�y�Iĕ�E|��*�K�b�?�U�E�4Vk�D�iI��X5��H�����2��J��7��l/�g�a2�E���r�x;wݭ�2[BuqV��uRi�O0�X���L��.F"���}���o�u�olZ��u��W	>ϻ�Ր�v����<!v�{�f�u��we�i�D`1��N� q��|���*Ǫ�Îa��t)����!�ت�5�哈",�l�w�CNRGJ#1�_����s{߳��!7j(�r�̽�_�m.��"H�ю���=��7��(6���v3�H�&�ެ�"0����kt�oP�t�g����ȣ��n{�r�id
,�I1�x~TY!���گ��#xƏ8'̂E٬� 8p����χ業�48���n�mpl��3deH=_,��W�<�w���@D��}}|�u�>��������Mo}�o~�9{��#�t�7�I+�ǻ�XV�g�e��K:�8� �c�Fæb�b{]��h<o"���kEt������Y˭`8L��ܧ7�)P|�seJ�C:�YG:�芬���K�yC���T��n���	L�촊*M�sm����7�dۚN"(�9��˫
�����0iR�	t���˥���7J�즐Σi��h�-�7��O�ݝ��]k)L���r��*^6s�F�noh�ڋ�A��"M�Y�x>�|�V"�}u�:��-kҞ���������B�R���p�����aF�R�qh�";rV"S*[�m�]]x��]��1�����P����*��K[�K�v3�����Pm>E��<����ө10襫=��޺�S2pFB�|�L�!Rh�r����Ν��Js!�V�iB��ţf�
���/*f4���Z.���|��P�K]��1|�`�w�����Y����ّ�ԯ��w����d�s�� ف�犲P�ܲ�^�P�u�3�`{��Wڣחu�^8�'s�u�n�1�j	��n�F������Ju�[74K������������ DoN�RT8�^A]����Ĵُdi�9g�-]�������]�r�aKN�œ��ޓv.�*��-V�i�yӓPm���m6u%t�\��**8�35=;Q'��u���bي����z'H��;�E�z������`�-e؝ŜD�ؖ7���+Λ��C;@��.�h�F_j��������l�ۧ�goV�d���T�ʹh�����F�`�����;��C�|DH�'i��$j�X��ӣTr�<�#���VISa%��M-߷b�۷��z�o����`�JŪ��Z���f��n/��%V�t��T�h(��(Xw�ҌK77��!�J�>a	N)$u�0�7.JC�������DڍS2�֫D �_���P	c���u1W���d]%���#��
�y��>v;̺|o>Y��k�4��;���í�ywlt�-�:;���%䇡-m<]�nq�-]�9�Q��F��zt��C���r�e��Q�	"k��7ψ��Q"�>����S�S**�e�o�i��1a��TO0�ڄR�!��苶aM��)H�wt�jc�zt�������{�ݫ|-�ܗG9�pmׯo�٦�AC� �O۞�d�YW�El�U��v�4y�dr�1�s�zǺ�+#��l��m5	�I!�:�Bx��D;�m�S�6�g�'�lC���ʧ���Ձ���e�S���[�=_v�h��[�v�o�wt���I$��]P:-��XF�ּ�6�UrT��I��
�zX���:��T\E�jY�9m6�G�p�����7�N��A���+���{KPv�2�x��6D��V�71R�י�WH*<�$��r�uL�6�fs��'j�9�.Y�/�����8��ٵ��,(1�ޝ��+.V���e�y�&������eo�e� $H -�^:t��w�TN�<�gqBɵF�Z��=׽B��|�[��M"�"�n��[}3Qp<{H�̙�NM�1�����<����gD�i@N6w�26��|��z��dMuaV�ό��B�5�u(�0�)�bH�������q��"�����|�k�#`U[ճ�}�}H3
��5;5hL����Q��f!�����W��[��U^�xm_�Cf$�@Sp��g�5[�l���q��x�b���(3V�
q��@�\"�Y����tȂ�/M�,��U���J�d��������pm!�M[�
�W��w�Ԍzt���i�,�k7�+T�(R�Ko"���x��w�,��f�Z��� ��V��� J�إW���%D�t�T}�Aw��	T�P��2�os��e�\�7!-�7���4_8�i';���U��yT`���ɧ����q�� ��<����(3y4��W���G����p�x�1�/޼-x�L�l�c��;�=WpR@0ۊ��
�U���l^_u��%���s^V|��A�F"{���tzh���!E�e!+�헝�v�D!i��y��]}ly�eŒǽx�t�&&�v���]�kr>�Ks��]�2��N�>wY��a�����ͬw��P�r7W��嗮j��v�����}��,�t�d8�J8ݶ�^j��.&�z�en�n��r�����2d,�m��F�S�|n��o8���M���ou��齹q� �S��U�ݎIU�O%�O3n|U���'�OQ�8��]����H���kn}�������[�z{&�mpjz��'m���C����J��]x�:]�ێ���܎�M�ݟ]m�	�u2sm�Fy:�G/l�[���3�>L=�Ç�#�ٻu����VVkïU�X�r���CO�\�,�$t���Xuo���.�׭��+�(Eя{X�����������ҭ�M��W��q�2���ږG,�c,�RKy���2��7`�<^1��;����{����iy!MR��'7E�]�����ݫ�e�/
�H�+~��2����F�^h�\fgE�� �W�@[�����"�F��ЈF��=v���>ƺ��]���y5Y�������0�]�cۗ}^�W{>Ǫzc���o-"�q�$�n�o�X�+ Y���E<<�H�Rz\ׄ�3u�X�����2�H��N����y���ٯ�/���(x�Xy�F��0���L(مIn�/x�ܬ����(C|�wc���Λ�qhJ�W�bDH/_MFS=��z�w��_��PP Lha���fG���l�R-���F�gnn3��z�Aî۵�ٻ)<y�5h�1�s��3uA�A\-i h��~}�L��Z�ʕ7{9W��I�fc�.�ż��g�ϬH�޹�¶*�m#�%`'�@��U	k�����o6���ov���z�m4QPrV��xY B3S��i�h�y������u�zZ"E~Sf�1ƕ�Ґ�)l��	��[�KTd1mtz\�5Y|mv���`�H�畕4�Q����4�S�0I�kCO!f�D�Ѡ�e��4��l��*����j�o�z�-�0�������k/����� Yd�	����u�e��$�\����4o4��:@��/�rW/ʒ��zޗy�{�D3͢��v�UKHA�f���t7�HO!���ڿ [�I�#��NA�aQD�9��/�
�{�Q���P",�*#*�2^�갱a�� +��*_�ܼ��Y7��MƐ�ߣ��%���������o�Uld�d���fa�*M�֩�b��fAP�	�P�1)���T)�����\�k=�wE4DX�R&���;Gʏ�s�3�����e�3�F�k�9�}(N!��o��q�h��֎y�l�W:�1pgqs���5ɳu�����vS���L�uJ�]MO�}��%�^�VnKv�f�"�~�k�z]èqT*uF\�"K���8��a}S|[�;�'&�����E�� �P`�ےXÅ�7L���!w���CH���=�Q��(�� ��T˫�xf 
�� �(���{Xgޗ}Q1��\�D^����m'�1��#:W@	Fd�$e8{�L�}y��o�b���4)n�/s����{y���
�����w��v\5{�`�P_v�,m�<)5�8wRA��A1v����3�z��d3n�븠'D*�7:���yG�	Hal.��/����b����Z�ma�Q"�솷���;B�ٜ����L��|֓bj���mrZs#]�\�Ǐ��9�V,��Di�A>�E��9f�/J�͈����cY��!JZ��Y[����*��!%>SB��x�֤yF���!��t���a���V�,BZ��hy�s�5j�}7��I^rYgз�?��Q���aY���VNH���Bʺ�
Yp�Fy>Y�ރ�p����ieR�]��a�ݎ��n���%��7@�\��x�A�t�.Id��=�� ӌC��}�J��J�򞊺�V��.�f��X�/�2A�oC͡�������
Pn{^f7���K��@u�f���Z7�=։�N�U�������&�w>�S�U5[�owb�K�
���eFeY��U7	�����Ȋ]���펂6�)\�l$�e�xM�G}}d�.���)�KC�3<%O{�/�)a�m e�l$i�b)b�Er���;y]�"���L���O����g��/�";�e>8�kxz���0H����r�Jr0gI�D�.$`�D�_M��`���=�]n�3��懶���kFVF��s>M�w�j����Qi�Q�#ܖr���Ef���!5mb�ȹ^�c �ů!V��P�]��|xmc�6�w*�S���{�O����@��t־h��eJ"XKn�m���C���9�2#N�
�v�E�Ⱥ����\�
P�Bj�W������E��P��^�uxC�!A�;�!��O�t��mΑ5d���%���m��k�ڄ��n7>s����0<pG8��)]�����	F`%#�y�F'Lt�E#o6�g[u�#�9���5����l���lBgڪf:V�맣�MF�,30p�TF�}�4,�N.3��h���(�L��I�]D��A8{U�B�[4_9xj�+D�����	6}!֨+w%TZ\�ԫ�9�����Og�;�hU?ni��N�{Uëj����͖�[�b*"�
q�ۆ@��9w�3��+��ܷ�j��Y��.��S��eNH����p��T��B!q��,��P������W��vEވ��G�N�Q��\=^0O1�}re{K�{�ڬ��tn�l��rc��>W�����h��W�,�*I���y�B=�}��������'����mFI���p��jm5r���j��~}����R��❅�t/'��x.��1B�*�YW��9~l��) |Bx;cj��b�W����E���mK��Ub�������zB�5j�Se�u�uI.sW}ُ�=[d��@혀��ƹeG�2�K-���f�:��Np�ih�N�����2H����3#�1qrh����w`KKj͙�]�-���\�mhBi˭����{O�Eg`�'�q׀۫��j��;�Ә�Wl5ґ���i箋�i^��g�Qm���N2V�ػXv� ��Waw��}���r�8�;-��k��Н��vNN�s���櫲���;�%�<�:G����m�x��'3����κ��o�;���T���q�]\*��O\������kv{l���3nܱ�sx�#�|��g[0�ݹ���ku�1�[���w��"�>�g��il�\la	��(�!ه���fC{ҏY��g�-�v2����rf�N�ں�uE���7x%�p@ۋ4����F��^�u��Ԡv����'�x<oPlu���ܹ�
��7�� Ub|���v���\���x��gI9��Upd
��^���ݱ��D�h��+-���zjka\�P[�=��u��0Fa�h��8����.ͪsJ9��0�oiY��Ϭ*���������J���N�!��M?4ـ�`�GN�!h\���y��}D����Щ]n<�_�,J��﷦�P���qt�*y�{��\r��;���ɏ�{�8�SF[�����M��4�-�$)�"�a52
���qr�AM������wb�ŧ���޳1v��6Ә��#/X�p)��7ڽ�A�	����MC���yw���k���r���d�.l�.L���Q�Xz|��X�LEMݻsɯ4ZF�8��%�窧U�o�JE2cA]}�N����٢���WV-�!�T,���Mw�򁶹S�n��t��T���]���w$�)-�rۧ�3�a�6�TW�C�nEp����q�2bީ��ֱQ��Ņ�
� XN����m]=��^1�[�B
����CHk$�fsw`�Gӯ��oz�L�X��9Y0��}U0���*[�k�f��<HD`����}�jة��d���y]�,��<W�1���e�!I8���u)ag��z�� �z�x��Pb�c$gU��xmPe�j��b:���s�}�����j���������iy���-5��oҐ��-�Ea)���EU^�k�V�;�n�؍MD�Qf�����4��l{x�7����h!ѕn�j�w!�K��'���J���<�=����Ie�I]A,����@wLI�屢�!�3#m�����N<6��{�7�Џ!�q�J��\���I��kُ��y��B��F����
���B��X%�L�	p�.۰!>mլ�ٻqc�Q�+quZ^f)&Dq�$�<G{�Vy]��ů'��kL"w2��}�����q�,��/w:�5�I�xyiW�EB�u�^b)T����^���4@�b��0�"A8hY��4Y��v	���T^ՎC't���=6^Q�~�4bbiX0�`CW�`�2E$� �=����׾ͺA<�U;x�+@����7dFFㅷM�"���z��Z���ڳ��z��7MꨊCj��aj"�5u�s|���q�a�1��ܭ�� �Ve���N�MK"���M�z�MN��:aU9���^�1���<��"�t�Pz�s{l��n��+�Og|�lm�l���kU��VEOhq�]Q8�X�u��5�t1�(�!$�����5%��QcD�k7q��]ls�����q;#69�f�ۦ(H���~�Ӆ��.r"Cn'W����G�!u�F#}~�STx$�Ҭ9���ƞ^�|�B��a��ځf�n	��C"�K+Ʈש;��c�f��OI��Z���pRI�����3�-x_n��.:5�o`YG�n�l�xF^�Wg�4�V�� ���&��^{���{&��h(�o�#1 ����&pj\$���z�$Թ���xt;S�(qlɝ�P+y��.v"�r���0�d�
PF�点�����e%�X��bW�-���8P<5�(�ѣ�S���Q��;�MO�E���<�C��W�CѴo]�=q�{���/ݺ>�o��xO�����RR&T��U��3������i�m�z��]f���̕Y"�m�n�v��E����@, ڇ��.Ƥ<=	P�M�܎�y�)�(�������żb���(	@Vu��#��Li&؈A !C���j���3C�G�7��o�'�-�G�^��fb�[�ߍN�l;%SFJ|z�guj/���vԶl[cf�H��B�>�Y��a�V6���}��q>!	>�����k��-w�.>J�xUJ���y^9<��w.�筊��0]%V�IWWdϋ՞��_%���e�ӫar�S���NE�8#jj&)�D�6��.�tI	��6;gϋY�v�ڱ4O8��a�b���(��&9�����W���..ҷ!��z]@Q�.��:�dʬ�d^�[�@?k�ѵQ�ԏ3�`��M�e�����U���4o��m]���7je�x����&�	LB�Gj���Uj���ZK�x#���e�{����C�xӡ�k���qy�U����LUs9QU��`���(qN�q����4�.P�2U����j�j�@>�W��� ��˨׆f(HͷZ..�`�`c��Z����8�r5X���y��5i��"���C0�	s!8�����雷$)��*B�p�z
֫F��yh��}[t��=��}��^2�^�����ݳP�z&��`�ǳ�m�Y\��"x�A�d:�{1�z�o�P���ZӍ.]�~P>E�%l��J�3JUq����T���L�RuO�d�X��3�"���������TlEi��Po���A/W�G@q�%����^0.�}�k�*���׺��e�x��f��יJGX�*�
W��^t�+��yCN�ڹ�����]N�>��WYL���Η%�T�L7Efr���ln2�'սu�z�r^:P��=WB�ַ�0�ք����{hRF�bu�<�N`��,����X����7����I�T��78���sV�;(��z�Ւ��0�*��{���'W�ٗrHʘ ��avWu�ĺ��݌с���7��skvT:.�rk�N����&�aɛL����;��W�^A`��"z*4��;8�(+h��8�ͮ����iǷ5t�Zo:���L�uw�7)�k��eqգmf,�mQ��@�C����4�hޏo�t ]�9-�潑K8,K��ڲ���Z�qjL��f%���/��ӭ-�s�Gz�j೧�qf�n�>2��Z��ls����-Cl�)�CEh�p7]��G&e.���o9
C0|9��2��,�Yu{���cE��:�n��Z����D{�����śr�]	�3]�]NX�Va$��NR�]x��u{}�&\�r�c���e\��>����{�Sn\��Kdݍ����k����N�g9��f3Ag
�1�;�O���EZ���j$�gv�j��v��Az3�`���B�\�Y��V7m�u|���/z�.�	֝�%��ٝ�'gd�
�w���¶�Σ�y���j�X���)��:v���rtӽ;�ɺ�mJ%��LN4��U�h�]4�$�B�+0\T�l��9<s�������-̮h2��<M�5ً�7�9热*���g�:
�;�;.�ݬ��Z��J�oB����u�A�`�v���k4�l݋˲bdR.�m�M�po-ۋ� V�vcIz;i����hq�l�K��]Hݱ��`'���(F���nЬ�˽��G�z���V6Z7����u�1=�>Bw)v�l,l��>�Nw7�ہ�u�s����'�\n�/4��7]�����0T�G[��m��ɶ*��|\񷇴�rx�ݸ7\����.8�i_\@g$�������]�k��ܖ.�ۭ�Rg�^��>�kBk�4���� ���Чg��r\��aB�jKWj�[��oa�g�����O'���J���� fQ4Ny���u�Իv���t���{r��=v�wf��.������x�Tz8Ǡ^��,��hO.m�ci7j]��z�ǳ�q�7gv���<�	�s%�ۀ����zŧ�{w�<d��Z��yp'q�7e�	��1x�qjfם���[�l�L�����N��e��îܘ�\k��dg<uoE�2�mݚ�N^T�^�U�-�۳�7��F���W2���0�=�n���s�21<�nw.wN�1���hA�r�w's��m�Ot��oG\/�-g�kv&�C�n���V\��I�NR����ūIZ��X��!�{�-�N5���M&'�hcj���8�-�M"�t�r�V�e��6.y��^����oE�p`qb�p��S��]���A���9N��q�v��5��q�R�%6.���<�d�ؕ[���[����<�����7f<�z;0g�z���g9-(d1��\m�\��;es����=k^ǲ`�����yp�;EKf���a�Jg����۲v�"sk� b�K�n���s��W��1mB��;k��Нr�9��N�8�DKs�hm]�kl-��ZS�Urv���8.{շ1�d���9���%�@t�z���ۍ�b�rU�ӗR�f�;V�;N�-��v�Bp��a񹍞eY��6o.�W��G�Ѷ5nF�\;pA�<h���5v1��!-&��+N9v�n^(���,=�nvK��u[�"�/I��e�G%���j�M�6'�{�oI��:�/;l��^6���x]E��ԁ �I�pnf7#��;����Y�;���p1��nĝ+�]��<#Y�W@�i�X�n��ѶЮͺzWl�==hT�j�m�SSS��@�h�G\M����^����A>�2j��(h�y�/]�r��m�ٷ�Es����|��vx�!��O93�� 3݁����|��F�ʝ���K�a�)�&_}q��M�v�}�t�X��HV R�y�R�b�9.���%�[�l�X�Ni���j�CH����rDZn	��r�H^����Cs�+"� #����	�Z/aI��V�H{�����X��R��`a����@>���V�6��r�C�a�
D(P5�@��b�K���3H��!�
������Uo�����ªu�@x��z*4����UM���^=43�Gii�����"d�@ڂB�1��\`	�]�����('2��a.��:k���F^A#��H���2�j�t)��uO�k�u�N�	��k����)KGhduK��H%+(�m���uh���kn��X�F�8��s��1�ݒh{e�qO7DfRz��������Ҍe�ʗ�^���:��O��/��S,UĂ�9V*�Y�^�\5N1�	�[��ʺ�_v�v��!�r�7�'���Pr�KV��B���$��+������z1Y��3�����v�rek��YM�j��V�]YZ�m��!
�cD[ ��y.i�E�*�[ُ�e�� 7J�߸'t�%'ª2��S�
��u�Cݡ��\e/TSru��q�h�e����qQJ*�;e~�4j�����Os�k�޷�Ir�-.ݚ�&-b#K<�]�I��M��z��W,�ׅ���]�Y�k�q�����^f ������I�tq-"���m^�}��Ԉ��Gx��h��yu~�*�!ͺX�Va���C�nb��LP�ذl�on,�֩U�e.	+o�;�_�I8�p5
r.߂H�H��cU;<�c�kVUD�b��x�� ��U", ����fk�����1E��ׇyU�Ul�8i��{�w���L�k���룚v�;NF��t���ۦF�76�p��.�C����H�X+*����]k�V+�QC�a�P��Q29�\i���[�Lf
�_%t��>{�ѻ�+l��Б��V�G)Be���0���r�"��|���R�i9w��B���{{������x+�OU�
���OV���O|�� F`���>���U��q��jz7��m�3�Ϻ��=B͹Il,��ٵ�ꄙ=[��w_p����i�D�ߍ	h2�<���`����S�`�����iw� p]Ӿ9L-@�Ů����ϳص�������L]���;[ �F�HH�����9����Ż����ɩڇ|�>9;��EJ�%=���H��-��qن�ajk��@�C<����fL-�5�yش6��6?V�6���Q�~Ҁ�0��4�~7�k#�����f�o�׭ٗ���U~��1��dBWX��H��kf��3T�o$R�"N��n3� %C�1c�:F\�:6������-`�x�պ_uZ�nȆ��r�Ev�5 �sA��8�t�Mƛ�0��]�0�t��'���Z�}V��3���|�{Pd]�'+�&��������Sخ7�w^�`\[���Ŏ·��Y���a݅Q�v�U�[U����<���IQ���^َF(C
�v��OJ[����ʢ�7q�N�����󙽍�Gg�T<���7�0���]f5�*�ub�f�p�FQ�{�cp�b�NEy��+n��v��8��u��P��?Z���:�ժ��N��gt�	�.�����;F)׮���<\�&���[]\����-��7s��䩡�xo��תߕ��]��r��I���MY����*م�]�ʢv�B��7,1yyi욎���x���뻹IK�ؖ!�[K��a���X��މӺ�QPT���(���A$n8،%v^2�#��⳪��2|��#i	!M5!�1�bU9�=�M��'+����q9=����;B읟m�=���p�4e�F�r<8@�TǶ�TW,7~:�S�Ր�����lv��tw2e�m�1�vY�omŋ���DWb!����IyJ��pV̤R>�664��X�1T��]�kE�2�ޯEAn1!AC	����j�����`����7�V&p���#&[YX��XڟFd��
�^��o`�J��3gj�Ct���ԙC�w�l�ӨQ�}4<o�G�&v��`k��<g�L!���l���쩎�Pg�80��Ѩ�����8"n���DJ͂�4|*�(��+�8!=qGDL��7Z��@��=���k�/�Kn���m�6w�^46f����a�ׇIe�P��IH���E����H�񧏢�{Y#�=��B���Ung���,��vE���}l����y|���m�@w���]_:�������0�7�KFƢ-���������v�n��Lj4���4&�5�Jx����K� �d��H�`���:�\�h��2ѥ�W�OI~MY�P.ޕ� �H�(�3����gte�ط�ִ*c�[@Մ��aؾ��F��M޽�׽e9��r�E�v�KG��n6�pD��B�� �V�x�3�[�j�q���y�NK� �ׇ��&N^ֵaS�+�cF�������n�b)�u�����v5m�ۚ9�y�6K`y���m<t���f��[�7Y���ӻ:�#��.����)��ճ[��,g�ڽ�m�U�A:�mWf(R{��헢ꇐ:Ӽ���V.j�74�먅����m�85{U�48uQ/����g�ӈ�!�v�q<�(�:�n�0�ݝ�����
�����p���w�N۩D��z�WI=k����")��=�j�&��v��e���#�n�9� I�zG������D�#N8�]��ٜ���ղ���F�WTz1])0)���V.��f�ђ/Crm�?�Y¼�^��||+ x��q,����D�=�[=��!" �e�s�Pi�hÍc�CF�ٵ�5w��1�N禚�Ȩ�e�͓� v�E=����@OZ���v�r۽%����5$L��!��"��%9�ڿA��zU�l�9�h[��	�}��d7���WJK�=X��+��6y����,5��Qz�e���XU��ɢ%v�c�" ��\���L�ʤ�:�ͯ=�V���4�I�e��Zf�=qtDL�`Q�0fz��zj/D.��7-;�5�D-��}�z�y�՞�v8��]���y�7lR2nSeuf��H�Z�y8m��ղ��k�;C�^�vx���
��<�t�ݦ=�j�;HB���*Q��۩����=�v�j�ҏ%`�rR����hzҵ+;�����5CP�Pq�?#ӡ�ApFL�$�$k �),�ھk.6��+%(`F�#B9��4�wu+����:����R����ە�u�]�)�N��Д�\�=��e�k/n�t6�!�I�]�fwoMr�Dh!��i��/p�eN�SP���T�;ݭ9�@ڞ��:���	��!��N8a��������
���u��1���J
gvfv�k�X9�!ޗB�K`S���"�j�bK�Gt�i�2f&P�¤���\��tZQA�EtW{:5l���<F����.׼��!U�G3<<��w�a�QwK�"�+׶K������ԍ���q�
�*!״$)^]yy��b�[�fdL�sa-�I���`h���fD!�n�T̣�dH���`�̸b}5i���=�㾅Z��No�%>R�e��Ib,��ic�]�;��qs��u-d�y[O���[����-�l$��"=}ڒ�5�~Y���(�>��9)\�;	W��6B��u܏��O�~#�gc�*��XhS��՛J����{���@cjGaև�f���fV��ٓ�+�\'42.��'�ԇ�Ξ�����&ŕN�3X!�BQ�O���XZ�z�pӸxH���]�п����S�0�.C.�!y�s��<�;��"���烇�>�D6�7�/'K���]��۸��v�C���=�[�!�=�v���hv�m��:@v�yƦ�����a�ū��#V*.���n�Ȱ�Z�\�N�M�I�J���jH/vzQ
\���v�f�3f�UZ�)Ԙ���\`�@s�b�a$}xhC�\�K#q�~jL�	���/̺9F1��;L)"1!"@��^.�!�VE=����")`ǺP���ଜ�� �����؜���K[TU��G�+�n���S)0��NՑR������Z�����5�9�ݩ�)+�[�q���7C���z`%�;�=2>��)E�u߮�����;��j��!��bL2���٨�;�DYa�%W�Y��ז���U��������n �%$5YˉI��5
���Y�k�,F���2��B�WU�\5zk��=bA!@�M[3��n� J��F:2wcD����(1K���z��̉��%��1�[�6~�N�O+(��]�zm���e���X4Z(���|�C��j� �M&�Ŷ��tl�Ge�ﭢ�:$H��݂n:���!-�ywjf�>�{�F��a۴rZ����&��'�.[j=8�)ڳ��vu��'^+��u�wM��T�ë*u��W�CK��������Ρ����pn�ie���Mo)j�s��<�����V�؋3�׃��e��Å"��i%��z���*��rllX��������g�.
ߩUoL��)��:�!��������p6ײ�n�f�^C�Ŷ��F�>�m�8�ܡ{Am��Z2$`��6�n^����vj��GY�']mX�c�����aD�弜�^Z��(�
Q�.�4���ы�ϩ�|k�x�%c��QK{^���Tn8һ�(���<ӓ��ӵ�Lv�[w�Wd�V�4�	t�����m=[q�Dٱv�Ux�Lw(L��4q�<�x��uO&I���ʱf�,�W�Ro�g���7 $��4 $'æ%U��u��~엾�Oe1FU�N�S��NK����^�u�B�%�����ć-�$�P�*9N{���BqR *�,�3����
�ۜ����;�_R�L`��jfW�յ^��Ĉ���Ϻ���j�<%:up+���h�Ñ�9�-Őa�ݤ+���`��r(�A��*Hs.]P�]�E�����(|�q�eޅYԧH�}^mhU��Z��>4'j���A(P;���ׅe)G/�X�+�2�dB�	�wb�2�H�-1VT��
�0�}�`�B���3@����Ņ�>�l�4ޭ;ү��]��Ox-�#Z����Ĝ���/ ���nt��q���=��=�>��Ln��Mňkvחm���yδm��:8��+�zw9t������7����+sj��>�	��u�5��͖'sx��/Z�R�;�Y+�Pq�"Fݸ�fl��e�X�gs�e�'l�{!۳[v;h�C����%���l��8n�vżs� ���"f���^�}�X�	;gZ�";.6�9�$s��u�-�`�}�۵f�-L��$���]�5$�;:���v ��&����n�߸v�',�>/mKq�ѿo�hX36ic�"�<���&���9j�z���'#�q��v��#�Ö��w��twQt����$�j�V�����6 t�B�a���)Gc����_b�K/Uv7|_OVC�]�:,�O�2U��Qz
��`��
MHhVg�n��3x6N[�Q�'�E�ٴ�� ��5R�H##a�շX�6utʻ�����wb�9�dFҿ5�d��a? �.2DRfj�����L�2{
}�4p+p�>���("��E����5f*�T!lȑ;uͮ�}�nT��F��ޭhf�Υz@==x.5K�֘�|ߖT
+��ԐP���2y��Z2���]
�Ch�Ω/��t�Q�Zs@���H����P��#<��^�Z������*G"s��t��H-�G�,s�����[7�Wg��<toQU�c�[s�S��T�n9EF��K����T�s�,u����e�fH����pt���uב[J���'A�}.*���hʬ��y蹳ٖ-��±A>8ɰI	ˮ㊕h�^�Z�8Ľ�4T�}^_K�vv�W#!����K������������X�ث�
�P*���zE����`��1�{�;q���F�c؉�N��-Li��J�����n��W�X���o�kNjU��-���_���"�B�2 �B)m�n�������f�N��1:ni�ġ�kx���`���-UP��t����ĠN |�n���K���k��XA�6M������P-X7f�y.�^s1�v�����׋em�����e�bP7vq����˾���|ɬL�u=TA�ff��I�����߄�ϱ+�V��]˨���r�C��8}Z�A��=S[4.s���Ҝ�!亯46���M�o@���q��1��E֡3]S��,*��<����3��뗔�qU0e޺�� [q��qw�8�*�[��:��5�$ �q��N�Śsn�N�6���4��$&do"���\XIF7��zs4Q��Ucy�	��!�l�`��pN���2��T��z��%Oc�����X�)�.\G�%��V�&�W x�ʘw��
�ػ��Q�m�j����d�#���9\��YDah�ԅG$h�H*`V\[�/a-�B�0��Ǒ\�4�Y�h�=6��{��$}���pBX�w3����Sk$޷j �fu���дu_��kw:ԊCQ�d�PA�޹��-1*��:�V�^���U?f�9��������uEl��nW;��#�ڝ�7Y$;
�bed���!��K��"��N������X�㭄�MK�=Ę�1�PР�5�s��5�`�9ǋ�nʈ�JѤ�9O���G��!QS=k>mIbJ��ˬ���ǊYս��mnV��$"#���tʌ�컫/F��K�T�T��~뽋1��j�J���a�X�$�>����N�,N/;��+�*�].IЁՕf��.��@�ˮ�#��m��moo��vw3��b���[:;N$*�C\��=��Xobe����;�{��mCw}/�Z� ���;�kUG�zA1��BŐC����W�R�@����w��܏����0朆�2dU�1	StY�9�XI7�ϻe��sg(b�1m\n�y\���T��Q�MF*0�DA�0=�2�&jx'z4m��pʉ�n�s�h�sw�XY}���k1�͇r���n�ȗL�������r��a��i��ц��i�y��7\�*>�<��Zu7_\G.�:��vkfʹK��/w��$C�\
�7ȫ8��޷��TZ��mhU0ݮ��%��S��YZ�whwY0��l�8��ޱmϏY���y�z���p5��ܾP��=shڗZa���Q�vq]EϊY/�˛ƥ9�Ra�%�v�n�m^�x���^�X5�{�i�roN�Q�{��%_G|(Ĉ�鮽�g�aP�D���5.�w���HU!~�Ω��m��)�&d��UB�J�v�R�}�nsu�K=����u���-K�� *r�t�L׶�e,a�U��w�"�±�yRPG���l�!�j�vF�qgW�T}6����Rx��O���ԝ��_�ro�`�{t} �]M���2��/G���������3Yg}	1a@�L'��3��(�1�c��F�5w$9��\��hh�a@ܑ"q7!�~��r������4m�Z��Ȋ�]+�Z�d,�1�E填�E^���A��W�p_,X�b��,�_F�N��8�L!��h�B�ڵ+|M��~ɛ�}�Q���GA�1���� `�=��m̨.�`�1X�S����}x�w
I@��6�' E��Ȍ�U�]�S!�#���Xv�7\�G��9��D[���nѕ��C�!o0{K��]\�������2�ɻ��
�ڔ5��r	$���A �Y4.涹���v(���J�(AF0y;�5���0��>�������go��W��\t[�f0��N��E�^���s`��
�ؖ��mB)a ���b�R�IL���.[w�����m��}ݓ��������M�i�ԗ�w��\%���������D���;�nMZ��n(�����*�H�g���~��u��%߂2���Eb��{�=ja�x2TJڮ�+�")���C��;`�Oa�kx���lVMl���Ғ�����"��Ҫ�:˩�c�L>�j)���U���Vf����1�̛'�gs��\"�76h�Y;��x�$Q����JE�_cUpB*�_
�v�J~��\1\����F9��J��w����.�^�S�,cެ�匔�ӽ�8tX~��:L��Xp^!Բ�����Kt<�V�y�v����O�oy-V�N�?-�x�];j�:t-���T:@]�+�,��^�г��.�����i6���J��!��w�ϴط6�6��?CD̙�{��m��ՓG6����S����K:��c1SF`��mA�U{��.Bu+T�2P�Yd�ΚO/�՞�|F���5�}��w1��l�{.�M	U�4򚱼[�cV�EI��U�Gd�4�'��)�ta:*?�f;�`�up^e�{��Aڹ�qf��Ͳ�wpt�X{T�#$w+
�<�E[P5oz�{;��F��][U�4m��w1@��H�� ��@j-+m�g��s��^�݈�Nm3�����ͧ��c��y���Η8X�^��n-�g��_!\L�nN�;��#s-�<����7P��T�n�o[�mǃ;�c ���j��z5��p����`�8��Ѹ�:� Sc �����.a�t�l�N�\g�l�k��=�]�ܝg��uq��>Ռ��b#[/[=�d��b�ո�z�q�Y�wFȷ9㛝l<��ی!u��9��V7
mѠ��6�Y�*՗TSw9ٽ�^+����UVc���Ǫ�f��۠�k����c�q�n(��w2$3Y[��B)a|~��S�A��_qڦ�	���ת����\���{�]P�+���<�_x���+z��um���̗4˝P�='�9�띪��}�لm���F܄�"2�L�����/��xo[�~��U�x���������l�3�q�o3:nO6��HbP�v � �Miڶ{�˄@��aL)JE���Y�������w�}�nx�e��~y�.�wd\oo"ś�1@�����Y��޽a�%X�&w/'�px��⦬�w�����J��6y%�%�E��=�8�������iݲJ�.�E\�`$]�A)D��2l��[��#xsǥ�R^�*��q�]�y�;�U
ZD�r�x)�A�8��g�.1�D���m*fݮM�g�Y��j�g��鴣1��"KR�
.%/F�{^��}���n��{�BAu�O ���o�4�&�>1���
���hW�{jN�_eGNw�qL��Q$`1RC�oH�Q'5S��ڄ�>�3R�O0Y��[��ΚI��J��.�!��8�FY|����=8	����.�M�M��p�*Yb�r�억�ǤhiU֝�B�d+H/6|��4�n
�ϟG��	��i�w�M������G<��N��^��ڒ�t��M��(���p%z�����͗lbeɪͩ��z��+
�3vƫ&���Am�77��JOW�YE6�Q���;��u��?[�w�Y��(�]�>+�V���X�7�n���>�6�	�5;|�����;�/C��z��w&�h��2pa�����r��[g�O=fIo���ɥ|xΞU�)�UGɓ�ދ�Ř������=�M�i��^���yp���ɧ��瞌�<^������6�ӹ���<,c�k�k�-���6�$���w�7k��z����D]v�p �S*�2���X�.�<�h4�8���)�i��k����^vR����V��N9Ą�F᪾&z�n���ʃ�^�]̚b���~�X:"��	˼1҆�9C{��M�:���̚�k[K%n��)�P�LM%Q÷~Qbc34T��M�U��VQ�+[���ן@���%�����o���y��Bۧ@@�d䲓�VU$i_��(�eeJޠF���9m֧:'y�!X�6&E{��[�j;�X巜"�T�H"4�U^��N=��];��*��H*5%Hv�����B����)�'�ชeL)Q-F��;���aX��zVd��c6��H���GɌY!�3-����o����$F`)3,Ĥ#i���+>;x}=�rQ[h^��I���R6Y��7�����q|ԹAz�S�X֯K>C�Ð^�rdD�4��ohmr��]�������M�6؝�ٛBu��CF���j\O\ɢ)�v�� �ڠ9���&d#��%:���r��
���a���6z��;Ϡ��b�?Cxt*�uВ�K���Wb���x;u�� ��Xs�$Y$/{�]u�������
���n��D탒�5YٽLH]�ЊU}�x7;8��.Dxѹ]�u���R���Ws4C+m�È7N3!
4TE�xn�2�I��k�xl����e��6w�5�UL^�Y*����u���i���T22{/�}���XM�oaͭ���o�����	I	�!�Rfw��*¾zJ�]nOs����L��^��d��g[x�w�@aD�G>�*��Q�\���B3�j���Ŋ�S���i�جO5���ӓ������a,��S����׋p�?U_����VW��0|A�@r6�;��h��J��y��z%l��r��%"3�6&�nY���I�����IUf��w��!���Z2Bn��e u���~�x^����\�P�3����^��3�\<Z�uqLi8,h��g��������7�����!�^����v��U�%��p��[�h�!�_�J���A�~�G޲�u�"�.��ҷ�R�E�[�2��6�G[H�_Y�]�O?k���L�$��x�f�[�����I�D�3��3 �	�"��]�%Y�T㷻��o)+=�^�)��l�m��+B����Z�'0('Lu��t]�{�a_E��*�@��Q�zd[J͟(l��esjȯĢ���)��Y������eb�t}��/&��L��E��Udæ%^+%��XǏ�7C,�j@{=RǊ�9�\�n�iw$h��wW�'2�C	�w�}u5Ex�kpװZ�1
����w
>��N�0ҡH������2�*b���E�9�p2,P�c8��u�}���P��=�л�M�xڷ��n�q��4���fg}���9v۩�m]h;���30�-ceZe�b�MMmF�mn���C��'is�^lp��]��c�v��u$�{h�3��ܯ��CuF���܉a�cn�s�ї]��8�/cۍ�	�>��bnx�=ieV���r�<�gn�V��9�����*2lⱷ��oE�\�t<n�&���n���6w'k;m\6۳�ɲ��m����q�b�!VYp-��{�뵶l�m�nx��֜[p��$NͶ�>;an�Z8�(bv��D�[��i�ݮ��%R�}����z�vv��o��33��$^݊�Y�\�I`���p~P2� ��m�S�c�x��H�Qv"T[Y@���a�7d�:}�����m��������bP��:L�A4ob��ʙ�̳��0;1�9��k������a�gr����2`"RR#-�+��n�z�ywv&}N�]�nuGZZv4��\�kfA���՜��b�e�Ǹw��F�0�k���RD�$�z����pl�{��=ӽ�yml36ǅ�������+"s(mQr�:U��(��J���u�������z]�k�d��ox�[�D�l�0\�31�fu��������ZT�	c�1�<�|���n�
Yڍ&��X��
���,F��Ջؐ�h�\bS29@�����n����z�m<Y3�w)ԝx�p������Q�z��k#y��"i���~1Sv���,�0�w�Sa�r���B\Dv
�a)��$p�xQkV����g�L��%@������<��\�.�ܧ1��liq �Rx����l^��Y����lJs���}��˶���M��mL�N;z�w�Y�,�
I��_:����m@h����N�J�}cwr�������lP�Y$���a��ٮSc͔7h@��}��ylPQ�bS��#��3���E�w���<%ܰ����%S�j�N��_s�K�07�����
�����=u;�]�H�":n��*�ц0�!G)����ފ�E��خ�np`GdKK�:ŀ�s99��٭�ba7��{vA8���R|
�>𭷽�뭼8�^$��b��qf
�����^w��]W����Vv�\OyyD�J6�=8e)�S�}E�իT`.�R苾ʜ��>�g�j��ݽ��:;ċۮ���m�C��l�;B���ok�]F[�մv+�mjIj�L��vD!J�Jym�W�uv�V3ǳ��R��T�i�P�M,����6�Wm��we<��g��o���U��]v�[�V=�J2X���8�\d��q�5NUb�!#�)�:�g�;
wZn�v�+:FE#Su�n7<}��Ώɽ0���^�+N���WC0t`�V���т)�s��
kv���L��������ϑ9�+���B;�&Dp��W*w!ܮd֍`Ɨ�/�βS45+�{ku0����NF����W/.��{k�S?�����\�
�R���)�wY��YN�ͼ�'�y�t�"xlx���]�I�]�q:׹�L�$�>���:�xq�G���y.v�k�ζ^[�b���t'���
 �1�ӵrga�s��G�QŲ���|C�'\!U�
P�q�8-LX�3��w\*�½1����:[��������h�������ZH�Q���E�M��������l)�������{@d��f��I�뀶R�����eyu`�y��g�f���
Edkw���SC-����9��`��,,����ٴ�u�Z��e��o�Ƴ��P���ۭ0xOf�"%�0o��nކ�Z��N>׳���v�_.ᗳ��{P�(�:*f���*�i�|�d��;~Տ9U��Ok(���E.@��8�L��r�����S�v@�ӰF]���2��E�}��^�+���7����+�^�q��m��n��5C�my�cQ	�ݰ���2"��oF�1�wA�;U&�ʠ�2��������,�P�oe�3�<�C`)g=]�-�;��v�.���<�B��ר��gZE]��l��PV"�}ֶ��]&ޛ��
����.�d����H�W��W�^��lW^��yG�ie�cz1�AA�aR:yR�:�<�J�뵂X��tA�Kev����\�Ug��EAML/+�&jc�Kssy)�r�O}����H��*g>n��gb�m�]q�����q ���VUls�O��N`஬tv�kuTʇPZ�zY~�Za�ff�H֯7��<����Crn�Ul�P��{�з�q=��aWT���oY��E	f�����%�96	P^]o�xGW1�u��u���� ��>7r����u6��O�X�{�r��f�}����rׇ�P:⅐r����䱣 �ioO����-W��Jt����;�厏p��g��#��n ��~�;��U���vx��]�@��K�)��F���K�=�u�l\tc!j��=.�P�ywW��x޿.�Gה��l�����@ȟW�/�'b�T��E%��� m� b6��a����$�0Ox�[�S*�����1/bS�٦��9�%�d�S���W�YI{�.�s�/o�A��c��%��(��==�fc�:��z��W2��p��J�t�Y|"�1��鶵����\Z�me�O��w/7z
�H����&��V/m��Ze�wGrA���k5>�L���(��V^^�bi�}�y�b�ګd��j�K ��{8�i�[]2���p��A��Wľo�v`óz�h�+iҫ�ȝ���[��Hj�ǽ$��l�S>]�\bT�`�:����tXvE>ݑ���B��eK�X��;���͚
����u�&�6\ޛ�Z��͎��;�Ё��!�S��ڋr�dc���[�ӭ���ܺԴ�^�t�;=�^��]c³D{�a k��䶶bW��8R�;�v2�����"���77U�u��:�(�X�Ч��$)���._l(R��wc)�5�m���V)Y�4��F�v�.u]h�{�j/�@�3���+o�ES��@�ս����gtv6�T��1��y��Eҵ�^WGF�B[z�v�/��[
t���HG�A�����#�Ň���e�>���!oHCrmj����A�K8i�_e,)��ӭ��	��݊��5���u�xT N���l:�8B��e;���]gZf��m-�#��\�N*|��t5l��q����ח���tn�#�@�G�pr��-(2�#��x�(�^��X����#|z/5�uHAr\��+2�X�HNV5�Ʒ	Jrh�͙f��H{��x~%\;�˔���Y��Ӣ .b�'\=�^��2��Gp�O{7`�mS���u�pa$�A$�T�1θ��N�lh�1NwXN��c���R�++�)tZt��[3�[�\n�����!���;���yM��lJ�̇+�G���p�8w��i���n彉��ݣ�lI�ͻt�!���猡����ĝt�y�yݎ\�8�V�ҧ��0e(E�Rvz�]7 !��m�Ef�ɸ �S�j��0�vۤݝO�qҦnԽkv�����o>m���c	�!�F�od�!�`�M��lu���vФ4c��w�B��l't�u�6���[i#&9y뢊ݗ�>+�;s�G�um��x�hڷ9��������%�;r�w^�=�;q�zv��m�4s��0�vm��d�^��g[1��]�l�1�n]�b�WN,��`N���	[=������	�|k��ya�Γ��!�Ss���ǵ������8v��㮋�v�qZ�]y����
Z�s�rg�m��5��S�ّ-�^�9��s��:,���uvM���U�ݭ���t�݀����$^��OVS����#�W*�v���O\pMF���n!�v���t�<mƹz���qQ�kt�%�^�zz]�ݵ۠�cX�w]���0���v݅�h��;m����z�rr`�;�]=W�d�\6�8�{O-�\�͹���v�";�N%�7׍q�8� ��d���Juۍy�q���n[�Z���֕�I�vb�[��m�$[׷n,��ug�-<=��FRGY�"�n'Y.^�\�;2�OeNL<���!��t�J��S���{����u�[q�m��"#��nNƣ�u������$Ҝ'[�^�p�#vD���;j������pk��q�;����l*ܛ��v�kq!e��m�6��OZ��FH)5v�r,�����
	�	S���=uk�lh�wx�����۝ۂ���[+��Ү���(c;V\�ㅹݞ���qE����W��m���X�L3q��Q.��Ấ��m���|j�GO�6��pA�񰮗ۧ��8�]�bv�l3��H�]���Vl�,����deݹ��sl��;J�l�u%�K�cƼ]��q��5c�y�$�;��Y�N�������C�R�n��t�rU��ix㣹��pq�2m�넸bq�[ܼ0�CM�u��W]��h���=v�p&J�9���}��ی���t������:[�<����;=�X%Tq�\�rsGd��Z��&ɐ��n�@��;]7����d0#�[h�p�n�f{b��vk��A\lۓ��k3p'Vwj�pr�5����?��P�u�M�gM�0�V�
������E����?:~ٮ�8Q�\U.��'��X��}���Q0-gzbB�$H�SY���1h���;s�k�J�:՜��`-�+���ґ�#j�o���&\��{G�����x�ޛtgZ/ޕ�k;��V��(�Q����u�J5T�Kq�jw`˾�$X��S
�aT�3�J��3]ݪP�
�/q��pF"�����fզ�"�w�^ӱyE�@�,�T�V�����_P��X(��W,��"�W��%��{�ײt�,�o��gAgT�^�;�����N��gr4
/�C�n��vq(�6�.$WN����%<�N@X�uD�n��T�x��g�T�����[žr�K�f]>�dc���El�'F��t�p��2cR=M��V�������nM�[��$2�����{R������tڝ������O\9B�Nr&�K=K[����jEx����5�1��Өf��j�������m?y��R#0�".H�h� �O/V�����ܖm����Z�5�r	�X�nPh_;#y<���bk��}HJZ�7��r@O�.��9%J�b]���֭�o9��s>�k0�R`�tfk�=�0�b�C[r�C��[;vꩥ��fsbo2��E\	m(Jf$�J(�n
�+"�|�=�w�Y��R7�[�-*�9ۻ�ugz��)���%�h��o5-�D���M�\׋5��qoL(8��cH�g�7rfxm�E�p�������_��g�rmetM��c�6&_<�%i,PN�l#	�
��=�Â��2{�lyaj(	bAqT`x�u(Ӓ+'��1���,E{i���
7Sp�PDs껣NdV it���<aӐ�:GnH+��]wvZ&sj�h��������㩡��"�N��{N�Z�:�m��"�%��n��5��C�.�9��u�	�;����{���ε���"S�����YQo)�Ӝ����&�c)����'ݐ�A�Fv�~�7���]��F	J#���*Wj�]�|�ټ,�s-���b�3�fx�� /U-5�>�"o\�u��$|�i&�[9��M{��tu���g��R}� �h�
�&���J�)�e�}5P���rL�o�9�u��7�RT�oi��y��2�VdY�h�rρ�o8�����U�j]X�r�P	<�2.���/k�Z��Pw��>��lޏ!hG�2�����x��#��n8���n��{;V��kjҞ��(�'���,�t0y�Pӎ��Y����jqt^��˳n��ĻB앙=���&$���-����xըEj#Ზ���y%�������;)����=��������j]��]Ԩe�(I��R%kw6��3�ۀW0ND�y�L��z�:F�W�Μ�=V
R��-�����5���a�5)o������s+��`<t���vrVQ��)��X��;9��Rl��J#��3=�:��m��廛�Z�=��ߴ�p$�I���wu	�mxwV�S�JK��c�4-oagW=o���e;j5	Q( &I��T��L>�EV'��۹|ޓ�Ev���6��f�$�^�j༻������LI2������u��?}����������֙��*-Vd�0"=EQ��� x+�+��u%�P�bA�S����\����h��}ݤ�'�_I�l}�4S��0��kjЙO���In^$F�oQ�.�����v���q���Ͳ����ˎZ��-n�E��|�d�IgI|���E0����,�;To��xqX�ϟ���*VnG�9^I��UMS��Eb΢X�p�*�LH��Թ��/~�5��yc-�X���7@�۱���In:�Gl띧7�lU���H�Z�g�$t�^315���V,(B��_�g�
�x���U�P�O����E���n��:�\ږ��O`Y�%�)r�0�d���\uj���V�2��,벛��.�'`�T�};�{��7״�)=�ʀ��3�*{���K��u��0��$�JI#�6�k�R{{�#`�w|�h��ϱ�����A�d�Vo�K��k�hJ;[{C҅�inU؎����Q��:��Br��@dI��rz�ߏQ�L����*�Q�>r�-2O�{L�f�`^3/�&3F˾s�.j1	�������w[ٍ��d�3'fv�,�0�s&
E#���ަ���Ue]�݂9�w(\	��=�9{�~�W'59Y��1Οn���R�x���cw�Wb<�6ha�n��K7�[�m��n��(Wh�K_�5n���*.����m&Ue�mD9`z�Ƿ��`�٥���z��I�Y��m�����8�]�!�x�y�m�ͯgn"�'7��kv<�����V�nf#>���q&�N+a�͋��U��m���Ѹy+��V�\�+s���)�v;W.�{:S���]�q�G��Bۚ�����q�W����f7��۪�PL�	�f �����P:��Fמr��j��Q�����i������G`���3��[\v�)`�c.��8�v�%s�u��<S��1�[]�ڶ!�=lp��}7\r5J]jN\fG �'��Bx~�}:4��l��ko�t���[՝����d���Ywrz���C�yD�����S��k wDt�Q	�c��8��q6r��=i�&r�㕫�s��rBU�VM^�3A�I^ޯd�b�R����-�[=�̳������`�3��,�ә�ʛe(Ӟ�[���
�A_M���Y� ʵ¯���O#S�Fs$��^�i�SV�Cjokپ�8��$��
'$C1⎳+̧�w;�;i���8]NO�r!M>�{�Dm{ˠ�'s���*JjK���C'�:(�.7�"�-�#��s������5��!7AM!eq�fa��\<lLǍ���`��#҄/,o�?]�q����^ʧ=�j��&���>#� �S���:��]�.�x���*u�G�]��m���M�4Pm�HE���G�N�W!��U�w��]��|6}
�mEMwZM�+{�oڹ{��<+eў�V.���ox$�vǛ��dn1���gR�ֻ�7�A��îe��5z�
�K����/y_ iԄ��z2�澥É�*[��u�#�+�bsl&�Z�'.�.�����*a�W��7�z��|k�k�Ln�AHp�h63eV�#a_��TS1�Q/&�1�*J�t,�'�B.9I�:�:$�6�^�;�DQW~;��t@����+]7�}&��i����s���'d�¬[B	��)��,5��bL�V�ާ$�6 L%!q�;}�3�tt�j����#J5K1c�ڌuL�G.캃��rB%W3�gF��8��83ܐ0�j��L>��/l�V�}�y �� ��ղޭR.�7N5}�m*�dJqSg/1k��fV�2�S�o��ySkF�,g�^n�E�7lm��L>����%(�Q�
rF�y�{-�:�u=k�u�Nq�ek��[4�\U�R���F�r���;Z)��l��7�n�	FLW=���,j���}�br��l�ޕ���v/9�
�(�7��xx�ڌ��aC����WC}��g���ك�=����mA��O�
~Ÿ	�Ů��s(�{%�S�<.OA�8�=���l�4鉓*�h����7�V����=�]i2�fX�����Q�W��2����\���Lnh4�@К�>�y*!Й�����5�VӃt�yG���4f�i�kPj��,�/S�������A�em\^w�/���ʳ�2iP2P�n��y�3"�Uy� �I���N7$V�Q2Uµ���ž��LzJ|�Οu��1��q�#dlƹ��֓�Z�ĉ����La�gҙu��JG"F#%HzvW��X������0 ��e�yO�;���CJ�rڷ�E�zdOI�����"U���z�x��,�_[��ln������n��$,��z����:�^7]s7ا��lU=5����z���{����Ha|��!���!Z��1�7�q/x�X���ӕJ�f٫�uyqrF�⟑���E)m�{�8r�5.E��c��9�=@�YL�Ǹ�H��а�)��ۆX�y�g��C�d��c�{�aѠ�;�����vBJHRL���YY�_W
	�Z,`�JK����$����i�g++e���J�]$�U7{������=�@5g���NX��d¹#�:�|�r~���*�V�{�ʕ���P2f;5�73�e�z��s�2;"{I�'ʗT��p���}ެ���P�]���)K�mӽ�����w�h��mp3�\E���ôk��sDԀ�BT�M�ÎI^o�BGM��Y�~6�V�0��fv-!I��:D�]Y�e[�3L%��$��8�Tfϵ.چJ�v�;s��k<q�m��q�OɌ� ����ƃ�Gk��Đ&�gFA��?��Icg�3ziV�[/��vh�)t�nPx�\�j[{L˨�,��L��� ��Wz뙨��:Vv����%��Ę�H�qo0��E	잵V��2���~�GOL��պ�K�L5.�ݫ� =F���\�h���i@�	����$Wp0A�Uuuů_j;�F-*s/��/�M<��	 �kľ����D��4�'�u�.K�:�6o��b�G�b�:��8�p��&d���K��z��xntV�����瑱󧘃�#3U
" ��{=m�{���S�u,sj���R��r�.��䮪1�k�J���kY)�S6��YMv@ zc�:6���i��j#k�vŏ�J��h2�fD�۽rd���L�L�o��y,�gߪd2�,�9�v�b��"m�Vg;3�c-�*X�b����8-�v�<��B,l#7%dPK�o1�躁�n�m�٨�N)f8�y8Q\���\;�F*�R��&��@	�D���\��M��	�:�Y���ف�6�m�[ָ4v�e:x� v�Fw]�L�{���n[��e�!��e�L*�Q��u����e{=���u���nC7\���Gn'v'D���ݷb;m���a�Ϟ+�G-��n.A�8����]ۍt;<P���y�r]v;��{uX­��R[8mђ�[�1�﹛�fM�OK������2,[�$�G�m �l��sP��c:c�C�}U?}&�j�~9��=W����L�N�e��dh�D��.�U3��%w`���9J��qq��PH  ޷��̣$�1�4\*B�=k�~��eu��,��閭y��bz@>���V�P;gs��{ܢ��;���)��p��o-=�Ĕ1�J�7dgc��U��\2�\f�����Z��ihs��z]���,k�>v�
4J���)$F^߇�-�1H���pՆ��]ܹh]�c�8^]b�X���^��6�qy(-F�(����K��X9��7}���VS�@�f0�#�m�y�&HZ�6�RCl���n-r���r�7�u���hz��t�dtY5�4��FuE�錪J�T^cP��*_j�7 �	1v�a�<Պg�ƀ4�v��O���g4�G��=��z�`�{ؼQ
���������*�rGg�E�:�ƾ�aB���^�7}3�5|�S(�~�����%tw�˾֚�FHr4"p��w aI�8�x)��6u0MR��Ip�����ݗ��ǧ�	����Ҹ��,�Ap��-�z���V
�����%�x�mi�d庹s�:9��J[�R�^�����K����KͱQ�^��sDf)z�4�{��'7��μy��7q���,D�G �ͥQ�9+�l׆ZjsM=LT�
��;w�	�o2{�5��1p2[Ȯ�N�k�Ϋ�H{��2G
FdN*�fȄ�Ԫ�"F��Nm5�o���p�� 7I�^F��>%*��<
����ez=�Xʿ�/B�0E!/�W��[��@�}����]X�*Ry���� ��y'0Y4L�,�TŹ�>�C��*m�+��E�L`�h4�v{A��<�ͺ���F��^��a�˯�m��ע�{0�aJˌ���ɮ��W�|��jt]З��ё�2��a���6f�"yvV��EG9����$�a�\Hل��'ñ\��g<�}U)a}��C��B��#J0{�GEZPq|.\��Tj���R�X���X��)��v�,`i>���ڍ9Q�ʛi�e����oܱ����`B;hc��Dz�g?z�0���voK�5w�+R��[�=n�]/o�Wb7+F���V�=⦋}g5	}\EڅZU�̂���ր�d캸�o:��������F�
P#�Zk�Ų���VH��JjdXұ����WN��g	׉�l���^l���8e��l�al���j���!1?kꡃ1�$�ھ���7��3s4ѻ6m�����R�f��횷+L��S2���&IZ����N�.�(i��`����Z]ev۳�&�U3{�u5�vT��є�e��E��ٷ��O>Bӈڲ{;L�2�E�I�]m�[�}}�bݽ�Me���NFL�����^��}�(-����}�ΥΫ���Q���:��c�;ؘm�X7�s��v��Gf�Ի&L<���oZ�N͂�sغ�J%���x�-m�k���;\/�-E�KȐ�U�|;z�����NS���fU��]Xxh����{��^�7��Wu5��#����so�M&��w�b�e[�P歠�5�rTI��{��՝(���n�5lM�w����/������N��'v�/����ɇ:�f6������Yx�/���Gn�����'�>.n�o3��]�I�q8��C���[̂V��9�
�h����@�:c�-�ǲ�M�\�w�����A��j�\��c�WV�:obA�� L��:z�M��tcx����6���'o	Y���\�S�'TcC��y�3����L7o��QF�GQ���l��Z��ߘ1:�7G��Wdny��uw~T��E����BDBqFԑ��F���D��}��e�׺�]"�]W�"�Gu�U����� !W2XpZ��$�\�yP;��3��� .���J%#X��/!a��[�s%0c��ɾ�5��<�;�N�+nz+,l�C(P��4���P������uE���*eg/J�Nd��m�k�j����9�t�2抶:�5��Y"�@�2ھ��_�J�ipvDi��jxݹ�B�WD���K���j�G��i���Jn�L�	�ߖ["���j����8�J6��3�x1�]��@���G/�@M�V��������؊�H�`�6��U�/,�a\�n�8�J��f�M�2dBXRC�M&�[z�~����m_P���0�B��Շ.�ŕ*c�}x�i��Yvn�s~��l�'����VY��@[(8"�#�Q�݃��}��nQ��3j�^��%��(�
 ����y8��Ǖ��{'��u~Nfo���gG-�K�9�*��b�s�+��v଒��P)7-e�F�.�H��a@etږ��F�O[(�lo^K���67�;4�;�#�C�����1�����1��}�Ś��~O�&
I�g��kPu�s��:�'�et]��$]�y>O ^5��^\�s��ywF��\�Zh�����8���.2Dն5�Lfn8՞�H�	[2 >v�F����q�su���l�]*�ԑ��h�]�ާs^?���t�WR�Pʥ"�O��$ۻ�h�S��\ԇ�������+��J���Ҳ�˽W^��#��QI#m�P���*��P�M��qT��@��Fr�<�mƥ��O��@����n��S����f��맇ӹ��>h�Yzk��nB�R31#*ec<���z�L_�Ȗ�'��̄�{4A���[#;WiW�Mݬcγ�Rm�)ZU9�I�����e�&�0����kF<����Z�W/<�{+��Qu{wE�cV�p��K�6��JNF-7X�T�˺B��Q�H���1*Bґ�/ا����,ʵ�Ϧ��H��L.��<�]��:���n�X����n<��ky�,�@�}���_�}��z��W��3�ysCӺ�?����:��(v-�-x/�n��=͡AM�'^�v���{��2X���?_��O���&�\Q�K�DxW�vf���UՓ�n�3��\6���)ۋ���*mv�z���G\Y5ۭ�Om���=�6z�Y������3�=�b�n8�7nr�%���.2�u��V�"c.68��*����[�Ir�G��.���n��v�՗J�qI��{X�hs±�zu�<�#pϬY�dx6�玸�Ş��\S�N�NnMCƗY�!�o:뇊�ڈ.[V�]��o���ԛIZ�	gt=�N��&x�5tG=�]��rh6�!���!�7!͵_W�tD�C� q}=�S�`�s��]�b����D�b��
�1%���l��u	^4������Nu�T��*�[;��KNyw���&:�G�f��ڞ��9,�I���
�8�3����z�Ȭ OTq2�$�<�V�/q���,4D�2��E1S]�PvA ��`Z��0C�S������6X�35?��zu��Y�p�1�%�#5���=ZN�H��2-4��E�R	�����//�i>t�EH$Ghn��s&��ݜ5���DE5�[j9;,�>��Z�!��&H�RE�,�,Ɣ���{���Z�*ru��31��!�3���u-Bg%���`��4���m/c�6lO�)ڸ��%��d��&���a	
Q��Q�s��b5<��<푐����c��^������QA	R�E���T��}�}�mHTȩp��c���m��Sa\UXpiP�^4bܕ�N�I�grz,ZQ¢1�am^}Ud����=s[����ѓ.��o�j��5K��}�\����s��b����ɍʁ0�(��8��w}��g_j,���w�ɚ�]:�$� ���'��p��X=z>Q���feaȨ$�P�;!��{�E�B��2b���������D�Q�#C��ƈ*��@��=61�MEh��SfⱩ�MŴ�a����nq��XGT�dVS����$��Cܜ�Dp���G����t�1��>��v�Ju�z1�:�^�a��\K��J��N⩓�;f�rl���7�������(�,>������pG	mJ[��: f��lNU�·Խ�*�t��]�d��3`��}lfL�u�v{�T<��W��
�*j��{��O�;��m��� M=�����y��Y��v���*2u�/M��6�i�#N��Eؠ� :o�ӧ�BzW�0����Pp�����$!���V�7����*�=�a���7swewE�I*�����%$H��&��қ:�ﷷ��-q�5~�����O���GqRCƀKʗ�Ou;�]��m ��b¸jH��r\���r��{*��7��]Mۿ.���׳�&|���%�5C��ۊ�,��w�c�J��4.we�#ח$��^t�Y��|D���ε)�8¥����7غ��6|�p���Od�}�*�}�.�����	a6$j#���©�#y]��ك-����9+�K�6���V��0[�C #;[w��꺷��1�:�����(� !	�.�VPs�j���0�v��a��z�^�-al���X\U<�Om���ڐ_�14�m�Gn���Ƀ���;�s��=���t]�{GiI���ص�$��qۛՁ�4�~~��m��6�@S[q�bw����+�A�P�X��%��`]Ȭ��.2�Վ��Dʾ�T9^�*O<Vى�e�	�j�D
��`�\��߷��oǟ�dUfD����i}�dp�)Ks,dkw>t�D�:�w���3E�|pB������]}S�n�Q�{����&���.�.A��/_��Ui�t�k��J��Y�l\.*u�(���-���5p`��D�}�m���`
�ev�<O/KTZ����"��%-
yB���s��wr���7��Ji��ܵO1c���]|��'N�V��h�ʨ�E:-m�h��U����Q�M^��柨/��!"�{�X>�$�PE�"r����_���q�:��؅9�=/
���B�ؖ����QY�4��C�b;-r���[X�������Q�	�"@�)`�	�ڹ7`
�o+7.e�\nt��֮kVzn��\,���N�I-~۾�]�[����ES�W-g�����vj8w��.���c���?yv�6e>5��z��Ȝ�@\M�Zn��7e�?\�.�M_D�˶)��ћ���Xȓ
�f��'vl�Ui"Eŷo$i����eO&�ȶ��Xa��%�d)��.�%3�2.�J��'��47k�qGKq����>�6��9�.���o�����������ZM�	�
9�!��*���qUyMc�5���*��l��Sw7&"�}����8��$u��y[���oc�uz��G=��wЋ�B1�Ą�NE�o�w�nK*��ў�gF�C	����z8S~˽�Qk{�p���כ{r[�>�j�)�yl�n
��W]5��h\��8�>s;q�}�)��]K����X�Zr���r���*��.���ݪѭxw����M�JI�OLۚ|]���qk��"����M%aN|�`M�7:��'7zG�ٛsۍ�f�H�֣u�1�ֵ�v�Cۥ$��+���u�S��x]�Dx9�ۥ�����;�͟[�G��b냢�mذ	��n�I�����8�ɸ��w���c�gg��\P�,C�x4c��Z8�kur�c�I�cm�<�����s2�!�5iǮ���j�m�S�>�N�n$�v��O��.4�n�r�}g���<���.Suԝ.�I�;-,��X*�$!�@�'3�����K����{���L<M���Y8F V���� �6_q$1lzc��p�c{���W�]��1�^xp�t�2.0�K��+����û����ǝ��`s�P������w����v��tQ�U�i)�o�<d�@bL&��~S�|(��r��ٙ~�߇'�{ǩF�Y�!>��2[ׂ�c��e:�LD�ȭ�bs��.ɿ 6��M�"�]ew�#3Ūɽ֟Ys��t-տ6��^���P��1������i�,�>��Xl�0����wjD������rD�fG$��e��{����7ykT��H��qw_���<=A?Ťܺ�Sę�ʩrZ��,�V�@�~�S�a��}�^Ą�s���/#@�X�����苂��<��څ�d20�	rASS�{���Uv*��إ�
��U���� ��ř����qV'YN��M.
���+)*�=^iG�Ab3p�b����n��VQ�m,"�)��n�퓆��v�c�t��e�e�����#f#�Ӻ�p;���҈4����yE
]'-b�-u܎�7%Q□Õ�ZJ�Kzj�uK��c#��A�0�D��}d��@DJ����Gci��WKI@<���ب���튳s�Zyt*�����6e���h[�^�]���W�iH���ۑ�T�OG}ܩG��T5f�xkr�s�a<x@��ū��0䇕�=�W��SsM^��ւ"X���e.���`�5	28.2��=R�K�<�ܼv�JB�p�n����c!�,K�cD�lI�ȗ
�]�ƶ�$�������АqnͺB�×�Lۥs�#s/f���t�+�v'O��q:��X�U,�n��w�UUߟ���.]L1yE� n�d���4N��C���F.釦w%v�ֲ�zĵ\�c�S�R���	%�z=g�u׵��B�EH\a�*Vu���i�MY����nͼ�0�|w{Y�rP7=�9-/��ۄ�y~��[3���Ȕ�jņ"esk9ؔr��f�z�N�]@;�l՜A���㑶Qᚔo3�{���a6�jT,ݣ��m�����T����b��9�l��lX�G� �y���̝�<کzə�ޱ�3Z���Z�^r�:�=�W�3��i>A B	�|�EI���&���E�����c*��z��l2�i���L��s*}��;`�q>��ћ�ݑTc"�
�[!��"�p�F��z_dw�0� ��Nw	�+����x�E�fx'y
�t�n��%ZƐ��P9s�l���iά�iJ�S<��7�� AD�`ÍuΛ�vw]Z㛂p���c���L�rR]iIhC$M��+U$�cһ⳸��+3ηoF��9l꜌����3ڈTJ��Y�9-�LQ����R	 �Al^�f�\�t4��i�<f��!�f�EY����ŵ�2a�xzk*_sS��q�z�l��z���U��3&�	�.Ȃ����9������G�<:g�傭4}ȶsq�eJ<䝒�pjc4���*���՞SÔԶ����M���0�pF�RD�w�sU��G�ޯv׃a]t�x�����T�_D{ύ;ӭ5����g��̰���B��n&�C:wu0�ɥ��**�t���vnv���&#\7�k���\M潺�:k�� �nL����a�nʦ�7�Ę
H�T)H��3��;6a��-���(��פ�/P{�^�h��ٖs��D�s�C���ͪ�z��y|gm���gfY����ߧ:/j���؞p�Fz���cj�ӫjLi6�w<ݨ�A��͗��y��0�E�͹�6����������yO���u�.ԛQ{L�d�r���2ƻ�E�B\.m8��k���	�tX�a罊Z�b��̛�<^��Ͳ�g����Ѭ�J�oƦ�Wz�5�����6Ϻ'h��q��qJE�m�4{;,[5~>���]��`�<��23V�U�e�����B��%�����6�q�4�<GED&�^������Z$�y�jxj�"���I��+3*vI�[C��Uy<���붊L�+ŗr�d�%�Sq&�5}�͸i��<��vC�]�Svzy'�j��(#�/4J���8�d�s9\���/f�{�Lu���Gۏ�y�n,�,���.��{�np�V���mT�`u�`��n��DR���h��V+)�.�*E����c졣SOm�iH��wm��B��C��[�iex� �M���l;��jG�G+
���='P_NF�2�&r�uS�z���%�	q�[�K/��� �����quov�����H���K^5Q$/�gD��HL�jsܧ��;{tXk��6l�ơ���f��Xc©��w��$Q?aw�-�ȡ�vZN�HM��j��(��k��;��ٹH��i3m�땽��v�{
`�Av�A��m�ݧ�Bs^�U�VcV� zqVm A3V;!�d�!7jt0M��KyI���9�]���={�6Gr����%>����{��0�<��n:���;�ؚ٘oO<p�l�J`��in���;�Wtx�T�n��6k4�t�t����ۆ�q��D͆��C�2Ϥ���ZF�ķnݞ�ӻ˦���}�ޚ��C&��h"�s�����tC�H]��д�p3�z%twH��J��]�����F�Z [X�avs����2�	Kx�讗��.�>:嗴˃{I���7V��+\W	��SH�T��A����-]�X�j�h������N�}�Y�qξ�Ϝu�P���H�o(�SV�wj@���u<��vYFP�e�H�
��{�vm�߯fҮ��'#:%]���v ��o��*���nB�7�2
|8���(B]
��Y�4-�mЦ}O�2N�eZڋ$L���{0�k�b�uiza��*f��g�Aw2u�����d���Wm)cT{G+�8�;n=�����۶��l����2�]8S8ۭhG����s�Z�c�ێ�q��\���[	���<u��lV�q��q���u���sv�`ó�n�-�.�?__}+�C��mg�bx�;��3���O'��`r��;	v�m��19�ύںxu����x۫N������k�Dg g;�E���nťq�^яm��$n�Id-*΍�m7j�_l�C���&�����B��Nr��6�\���!�q�O5ԇ9qۮ)q��ѻ9�{F�r�QMm$�Lv�`���H��wD��(f,�ё%�ce�S�v;��1�Z����vtX�J!qq�'x�Mq +#�s��顝��{7S� ��d"��i��7i:�!R�7�ݵ�Z��cvIyB��k�U�9�e�M��,�6���n^|��}���OdM��X�S�9��š^�eV�b���HѭW�e�ySn��u�� Oe�� 3�qc� .{9�^�9-�ٳ �M��l.��s��<��=�V�3{�n�t���V�l�ͤ�!n\��݆�$�Ѱva�>�X�B����uېF���k�����.M�:�g�=mg�լ=�k;�N�d�pi�F�z=q5�#���c���9�;���ۜ�՛�n�Ht��J�>u�S����l� �v��r��qN�g�wRs�z�8�����r����rT���̒�[l.n3�c̼�ܬm���S�w vN�v{uƱ�`�V,��j�����t�a-�e��oJOSZ�|;]�m�^Ky�p/Y��Q�a��ݵ�ݎ�m�p�s�,ݲ�=��q�\mk������n۩獺�<��v��"Y�v�=�z����!p��vmٽ��q�f;t���_w�s=�tsu�=�]c�n�;�XC���КkKi�Ibї�r�C�vܴ�z��S^���x��@�d53/��I��yw�ɮ��*:�9͜q�''��[�����Gr�
.�ݜC��>׭��6ნ�8tץ����5��Ù=]K����]Q��!�e7n����%ٶ��q ���b�Y�/�]a-��+��=\lyګmK��&�F��aN�O�<!WH]l�m7\n�=�^U�����\�\\���6n�e�����M<D�s�bx�ᐩv��ע#b�������e���x���m���ozCv�����1p��]!�/�B+ʺ���OI�=�U)����J0BB ِ� ����.��[<���^w0軙�����c�6��5;$K�r�E��F�=d·��Jqoerݮ�;<�T���+3�2�$ӫ��}�/b7�^Ub�2$ډ-ϳ0�hi��]]K��z;��O_�����,K��C������P��(�Z��[+����/H�=o�о��N���Q���+�����W��˴E,�{��O^n^��DJ#ڧj/+$����m���Wy۩$���|,h$2�]�+�e���0�����.�a��X���ݗ�Dk��]�\r�EFj!��&�)�σ��qwd�j��=U��[u���N��r�m- �Fq��r[�5	��^?+㹔�q����#�9Z"I����h���{P)j�(;p�p]c;����C�}w��9P'$�(PH�e�]팩2�k�0�	5����P�!+�&��o#9�j@��ӵ��#�N��=/]N���h��pU���]� �y8U��>�&�EhXj�n��(�v��n0�(�E%���S4n�������Ʀ����C��7/x��^���@@$�j����ݥC���F4�*ͩN^��ou�N��Y��fE�����������te%3B�� d4jdI4Y�op��N�}�o<�����)/ȯ#��%�h�j��^=������EX4W`0�y��3����
$w�R��"���4|�E��^S��� @���5�ܝ鵻�L�*�v&mڞ>�ߘ]>8����2K�uz/e=���i��͖[�Ȫc����8�y�o<�ӂ�T#<��iz�Qۦ8J�-=�z��M�I9
ż�/�/�hv��xH5t�"��O�	���7Ԛ`{�ƒ��xY����6/y�Ia$eC"p��d� ��}0V�߫�����ؘ��Sw8QK��ɪ�
�{:�k�o(4��t;h�\09�p��Q#m9 �n3��+�{��M�<��E&ҽ�$���l�c��#��ŀ[���4{o ���J��ݍ��)�����e%�:OR��Q͈��:f�@���_y�ىԃ{�YB���?��Y�J��SU�|�``��Ŏ��G��y�<�Y\������r����:��G��Eͬ{�w
��s��Y�z[�,��#��-���(8���Uqιoɶ)2H=R�ZU鱗DeTW��̮\X��jɎ�M2��
�5�Y��^@��羠���&ێ�m����$�>�v�8.�&�c�����w�X)���o'gk��r�%IZ�iP��L���u�[��C٨�2W�����t�c���*{3E���/|�υ-v&�U���K-���EO7�0�>�f�&�����v0��1Y��&�e�؜���N�ގ��y��l��3%<�92uoQU��O�[�'P% ��2mڅ���vr���3�:��F��,^ xYг$�]�}�lT��{��)�ߎ�yƑM;@�P�$���fd����{�v�����ȸ����^��Սs�*�N-r �b����j�Auy`��4���>��˒\��=iG�kʻ���6�''c��ݦl�jy�%���k��T��x���7R=���_m��5N"�ǝE����_|=��UV*)u4����>�(\���j@��n�a���[w��Z8�0Y�o�^��}Fg_���ڠ3�r�����gҫi2S�w�=��I]; X+�e���]Ӟ[������uٰ��.���/Yk��V�`�v��7+�������b�����6����ؾ2X��ٷ��=�JI얌�tꇽ�)�	�����}�p�bJ�a���$��T	��rE������^����7'����O)Θ��^�N���ߊ6y��`��5,۰#�H����ͳ͋^"9��� ��qU��0�	��I��t0�c+v�ᚋ��
�}��w�[j�IVi�ǽO|Z���%[2�}�Yl% $�\M8���麞e�w��<�1�վ��yS4�~��t&�z��o}��jز���Qw��~35N!�:��y���
N$L��"qw'�z��Vʜ��d,#�u��	��sp�k^a��]9Xw��o�a3�k�)�,7�Qt<s��k��d���o.�V�ܵ���$��b�J[4i���/.�֝�̎C�J�r]�V1��gX�M��5��Mk������XQ�4Q:v��q��[�zE�Q�,�F�dg9َy�zy�v�耽-p��jqm���1g���[ٮ�<圪l��7�Ե��]e������fu����l��Ɵ�9�|�����s�bɩlt�c/f��Rۚ�4�����Q�@��Z��mջv����k=Z�zn���6r��W=qn�H<��hA�0z7g�CIq�,�e�=��f[����qD=n� ��G'�-��\C�z�bB��f��p���W�ܧ,��umd�c�b齦xd�g�5}�LC����"$�9�Y���.�z}��X�,&ʁI2D)l�^כ�O��5=b���q���A�1Jt�\�(K�. Ћ�=٪�V����2�����>�0���
��KlH�W��Hv��]堤"$�]*c�͉;�=5�9�=�:�l�D�$��T�\uVok�����%B�m�:��l]4J�E���������7Ƽknը�{�s8t���0m�^�%�{�'RS��R��(�J�<�F�	a���"�$��]�wq]U�m��Bz5�f�(4�p����Yi�G�ں�sn��@�Ƚ��A��ᢐ�Ls.�׆3U�/n(WѰo��o�t�v2ۧ
�z��'q!��Z�՝�KtZ�6�����![�������
������j)�]b�ŋF��@�O��]�{�=�}�o��l���@n��o[%a!��18��Y���l^f`��h�s�j��F)>��������l+�f�k���{ܓ�c���9��
\Kn�4�et�y�;dV�j�4�ݨ)�n����Q�D`d��
�l��VreL���v��8B��qk�e;n�al�e�}T5){�͞���\���I_<��׉Jֽ���fEV�
�O�ɡF�%>,��Ͱ�^E}[�3�t�]��@e�T=�f�XZ�������!�!%���	O\Oj;9c���㗥t����V�^��ʔ��Ԣ�϶��/e�;�ѴrV�2���y*�D�4�b���2!v.�	'��y��cY��''G�Pueٛ^Ŏt����K����~���ٔw��[��½u�g<��{�s�g�٭-�s���P,RIrYtD:���{E�ٝ�����v絹2b�&,��ٺW`�Q$F�����d��Կ#�+�ӏ3x7ygU9�\��N�c]ЯF͵�3����p�Í^op�< �Æ"ۅf<	�c{�WH��(��C�a�ʹf�,����Vu{8OeP��}��0���2O/�|���/��/@��*eVZ�V���m_��H�����,�"����ۙ�nu�z����������]0ݛ�[$�W 7*�����F�t7'�Yee�n���Ckkf�it�"3��F�:i^ި7���f��1Zz*[����i���� e�
��'��X�˽�X[��TǦ@S��8���ʐ���Zϻ�o�I�{�E���8w��$��Z��`2�UN�s�:�h��'UX5D��L��T*"V{=�p3$@���#��oI{=��wp�M�W]Ա�nUmv�'����IU�yM�1Zo{���w�isɠ��m'�;]X9���ߝ���)@�������ã�:��nzu��q�1Rg����$����������]^{����l���n��r�l�yW���U��H�Ҕ�Nﲑf�Z^8��HH\��[6o�d�o[D(��Qm[�M;��L�����i�"b���R�l�gh���v�mi��7b{<$�pR�>Z|��	�h�$���%HQ�9˞���LG�Zr�>m�u�I�J�Y�f	G->bL���k�E��Eˢ*)��n�C$�nzR ,8�.F�7��=W�V�E�hv����{����o?wu�=�\�Xc!����Qۅ-X��C�(9	���L��wf��Iwm�Z���s�)�IO��'/�(,77wY��J=�h��׆�n��X��)w���V$׆�+����I
MG�5�U`B��^B<�g	��q�L��ױ�ҁf<l
��j���Hw��>�yU^�qU�v�P�2�HF-zp� ��1wP��:�KV��8�+���/����rF��2�0H"n{xeѻ��M���@��srz�#UU\v^���.�8&1�*�ݛ%Z{14�wlj�N�:�����Xj)�BiHn��V��$�:�6��;.W���L	R�y�)݅���M��dMX�uMSr�/�jf*�ٖ��7a�e���rG����цY[����t��rI�㤔��T����:�_3��c��C�z���W�]�P��^6��mA!-5!8CӢ�_��>L������^�Kq��;�U�h��4��O6����T���];���B��N���1f��L�̋��q us���v\��7pS��^t�4�3;&s���X��u���U��6�Z�������i;,f7�-�=W՛r�dђ��O��sEHj#C6��}�3�b��oT�-a���s���<��n���M� ݙ@2;4C��g��q�K��nzw#�6����.�<�K��e���m�sd�V��ID�E���;j֣[� v1�6�y-T��F���9�{c��_�n�ood���]`��x7i���G�T#̓���\Wv��#svSk�t '��=��z���-t�����.��#���m�ώa:]�ۮ�2҈2W���˵�4[M��u+�b�jíK5��,*�ᄌ<�LC�ݝ,\5���y�r7a�n�+��،7l����?bU�?��J+���6��qL㩠�X{ñ�W�&�T.��)��5��t�x`��e�6K�<�lf��5�=t�B^<}�����QQ�'���4Uѐ�#$���ۉWb�H��_Nd*cM�=�B����JIH�Z�*o�#ٺ/�R�f�!�=�,���u�q3��IY��i=D�K����M�lQ��Q
Bb,8\rS��slfS9L`��W��]�F]�uoA�-\����nz�tr���Ev;빍+����+�F�� n��Jq�c~�8�+T�
���7Jwxu�O4������(�%k�P�g"}3���yy$C�����[��nޮ�pQȅU2ژ��0�,�lZ�K�ܥי��㝡��rnn)��=�nCg<0RH��v6�L�䚆;��1+l��؎��X�S�l.�:��/�^���U�「}��]�=GQ�0�-ɇ7Jf��u�=�2��>����X�l����\dc����\�آ���o����o�ͷ[�L�veuh��M!z�,�4"{���Z�0Gn�9���:�A�R��|Z��`*ɻ��`6�E�.���B�mÞBh��	�����X}uw�'��5K��5r�1*���g�wY!7�Z��o&��(�2,U������&.�8a12� fd�;q`��YuA=��]�����jX�7���u&��[�"
�J�o5c�s�z�}[��9����ՙww^y��~.@d*!m�!�2:�Όj	>����S2G[r���a)�Yvټ�`_�k��'!T����m>�āHeӼ�.�/��	Cʠ|L�yx�V^]��F����y���!�v���7���ȅ��]���RU���������.c{u���X�UJT;O��d��GUh�t�N�w݁�`�1TXhfg<���VsT�օ�JQ*��8M6*�%X�}��݋_��u63���&5����B�:j��6*���昧�Ȑbg[��ёw�ud�{霝��\B��ȅH�9$��^y����s�<��)���]f�0���ۼ]�}��r�����-iz�1�qn,+�æ�<t�V�Nsˮm����[�w����GP*A�}�i��Γ���6XJ�;V�0^�=%=%n�)^�;�#�-����V�I��5v���d1w�X ���¯��lBR�5ԫ��p�,�ӳ��ґ6WgaU���m���V�s�;WQ��y������ M�š^T�G�͚��(gM�F�zJy�{UY�������2r�ݍ˭3�TX[}�f�[M�xD�Ea�%ywt���\�,�_�) >iq�uuy��k�Ey�:^1�ȕݍ���/�v�Q����iձ��a[��W�",Q��3K�UΡ�j�ib[�o����3��hpD�l��s��Yظ����
�W��M]M�2�q������s���;v�w<=ȍ:�t*;�rVx�z��ց�~LB����k�|�7�P���B}A��U.ķrpwƮ�dT�i3I5�f�xM<�8�ӎ�M��q���W�>_>���oM�8����յ:����GJ���W�%f�<����n^��^��!:jx"َ"�m�"����ʍv��[f��eM�X-Cژ�� 86\��nJ�@��������3U�]�
�r�{K4��z��|��o�Ӽ7�Q|��Q�سK0�w!:��,I(�r�(��]2�K��G6ɒ̨��*P�/@��`/�"��K��ڹ�wH]���E,N1m<�d����ו�{s��1���{5/e�{i��u_jO��:��[�Uw�;����m�Cqe0�=$5�VZ�-��^fq$(���>�&�v�ui^ٝ���t3m/ �A�dsvè|�(��y{���gr�2�+4#Y�0NVa�t[�r�B������� ���@T�|����7z{T�Z�ώ��fe刼�:oX��Þ<�Zd�����t�O�d��!w=�����wn:�<q8*8�Ƚ�*4�I���ga�v���T.ϳ�T�v�pmp��g��sm'�E�Y�H.�A�i���uuk���绝��$������"��v(K� ��q�;�%jR"Z��2�ŘZ�h�)	x}���wOް,�AɒJdEXD|��u��� l�ot��2���ߏQ�1C��2}�HD�cOK^FV����&"�}�1Qܬ};]N]wj���ƽ2���q�!��J��$���n������l[1b�a��\�x�X�'�n�X����{��n4�pS#ə���ޫ;��=��	�Z�V ���	
5H"��B�aUE���+�vk5�{ol�P�f �4IN���kHDj^��u��j�E�~R��K.lK*���w���f���v0p�N�JkjX]��Y۝`v�b�5�����Y�P{"�9b�����<��*p���5桽��T[����ij����0��O��F���,ѳɽ�Vs^�����gU�ʂ��~>�$�L8E)�Ȝc�����E�e+:�����f���<�q�퐱ʈ�US�rT���=q�IΚ`��*d�]�ݶu�f��TS�玹�n͜#�&�6ue&�~>�7l����ݨ/q���;�@�,��Q[�j4+`��h:�1��`�9���עIHv�aNz�yQv6�'���8���J��#���Z�.�[��:�8��}��b1b������ݗ��3J�RG�������Б�Ӌt`��qC^�$' "0ڂG#wS,��3���s�sLP��B��b�R�16� V�vMU�s�q�+���/�)x�.�s�?P}j'���Kc�u�JP��K-��M������ݱ�c�Ag4�[�%�̩}�އ���.�Hԉ]�BϤ��2�ּ�˰bӛB܍�s"�,�Սݝ�H��H4܇�~`B8*��t��F���(��w��tˤJ�=�ɋG9�b�SlT�Ž��'�3t�S��]:W�vn�C�i�RyŹp�mi�3q�H�Z����cǙ>\�&�ä8iPc~nvU�2�Q��eiA<]�f����l�jF�.F�p�$��ڦs�Ї�G�����o\e�y�9��c�{wU�>���\۳�;�)�q��s���۸0p{X���#&�s��`v��;Xy���z퓔�nێum���������'��:�8}ga}�N�k��v��{su�Sm�8:j�v�Q�<��ݨ�����lI���kp�zu(i��4��w�6;/N�
NrD��rtcmɝnݧͬx�n-���77�������^�S�i:��q^\�m���sX�mW+B��:;4�����������_���t�X��8��o-=�bT�S�`[�f�u;ۙK��,::�Ᏽtgsl��[�s�D!�1Wh�l�D	��q�+�ˡ��<ˊ�
��Z�H�q]3��b�
�jh�
�KSYd�ظ�����qھ�0fw-����[εD�!��8���x�וy��wi!��G+o��w�Ytkқ�缕���l�^5m����{�,�+
�35�۪�(T#���Q%`�&�.8�3*��wi��\�7�����qI�U�B�Q�+mTY��8j��J�R��w��}]���w;��)���l;,!B��^�Dԉ�J#s&f/1d>�Yy�a9�ܻ�&v¨��]�n!t�r�)
{+'��V�l��,n斊 ee��̪k���4Ԯ���oK��w��:��!�qIA�*�n�dF'U/�,XÊۣs��պ4N:�3{R���6'gb� �C����&*�O}�`�����u0�f�Y`���;W�m'id�:�%ȡ\�U�ّ#G��Z�a)���i/C�	8ʐo-�(:��y���w�����~��$�Zg4�Gy�_ݡ�ᖯ
��5v�����fn�w�T�u��E����[��`�o+��<�UZ�=9��!0U�Z�5�n3d�����J����|M?QY��;������ƈ��b�
���9��_�R��R�Y!8��,'|W�8Go7����^�Ƙ�W������V�[;��L��5��F9JeJ!H��$r�"�	hgr�S#��U�>�Gy
������Eʣ��B�
�����`��wtt<H�E�n�Lϑ��c����������ս�=)1��hљY9���jz��>�
k��K2Ow`��Va+�=34d.�TX^�߮y���BQ��
&4KB$2l���T�u�}�������859�ֺ��b�sldq��&�p};\Ԩ�y�-������
!�t;H�W���P��i���˽�C�p��R
���O$#ί��+Ψ��e�$�)�Z4ф��;lr���s:e�*G�]
��rs1�:�$2�]A�A�.�y(�5���E�/���c6�7����E�J(�P�B%�v(_��y�"&�_�].,t����)G���3���� �t�n�*�̫� J>N�:&�^�2�����Y��mb��YW@����9v+�X���L�4Ǐ�GrZ2����F��9i���&@���BC@��p#�Q�I�ܧzk�o��<%��:��x��Ft��4����P�e��R:�N4'�O �Ԯ�d3�� �MY���o�4��P_�;c�t�#�\�}�?A�����f�w��i�N|��FW�(����t0k����6�oκ]��eZw���s�ۮĘ���<@��H�[��Kp�ee^��=kc���	#��Uk�����a�
f��V�$�P��d��ؚM�\X���'mAj%��A�xY� -�(<�wK�x区�l����j/(�;�E>��s� -�Ⱦ�!�w��y�vp�@fEMT�+EN71XH0Db�鵆v����6+^xh��Y�]�ȟ`�ۍ�Kq��	
�E�z�Vc��qW��o��e��x���>~�vܔ�c������n�9	e�@�6�fBa�Ԋc= ��B
�$=�+f>;�$���/f��6m���N�V�����^�L:*W/VZ����ir<�r��
	��a��@�������v���<����(Q[Z�^��������vx��Q���j���|�ǐ0/_��9l$��F��_��}c�]g7^4oփYy^�X�k㉃j�ҡM�Ӟ>[[N��w`	�0;�1�֦���4ݮ�[�~�'lB�8	fE�V��ymW":��I�wa��u����ß�Xۖ��u���S����׮"S<����`F�U�}���UI��dY�`�К;�]|1+'��;D�v ��$3Y��+4}��D�	��-@܊�R���{E�7;�L�B��ӳ�ds���W0��Y���	S�M1�[>]O-=��v��/OH=��׶��l��\P�Alz�����u\t��1F�yl�zD
ȥ���*>Q�w����ɭ�c}�"�ưʩF�%�ާlڨ1 ������0��A�$ZotI��咖�fɞ�	f'*�ž�}��@!��Z����Ƞ�r��vC5�T�-��z����s=:���T�_D���y��@��p���� w�9j���'*O�/1�d#nxZ�ɜ��hR���	l���w�kf�k2��d�;�b�R���V|b�(�/i���H+�ۈj\㛒G��pnA�:�ش���T��fpF���³�f\̭δ�8~�MU[��,��]��B�T��v9cW]uD��q�W����%W��p�(��E�񹻢��`��v��������l��r����qv�v݈�^��c0v��ܕK�6A��gGgV�s�Fn�h�C�z|o��Y��x�@/33��Ol�u�2���`��n�Ev|�rv+��8y�\jm���X���p�ղ6{nWt�T��ٲq��{��.�\�g��@ݕŉՉ��E��M�8��q���к��s��&�F8��g�!���}m��m�%�R%��4o;�0#��t�Jq��&P��M�J'p<��^���H7�����3ۡIzDҐ$����Y�{��X�O�1�6}�-���� ����g.��.1I�W�U�B�&�mrƠ=�c��[	c��X.��!q>9��x���H�l��K��|jk��}��ERF+�ܛg$����N�2��!����!d!sƻ�9�V:�q?e���g�R0نKIH���`2ǨbI��L��A����Z45xe!\}��Z�J=���n{qo��������i��N��V��!�(��������9a�͚���:��Q!x�a��ŭ�v��t��]EZ�3��[�Esk�@ �ݱ#���3s��|�̒0ȍ�c� Ma��;&�ON����:�uδf�S���\�0�n	� �WU=c5_g�]��eP�`��d�p\Q̾R��%7������\+��c��s´�i2>u�t�	2����@���p2Ғrq������حI�ö�1mLmW��-)ͱ�?
�u)�m�;b���
l�ϱ|u�/C[u�gf��;��CW+:�];,��3�sS�����C,|�)ֶc	���VE��+�W�o�����{��P��<ΞU��>�w��=�~W��-DYPD��ަ~�D[zW�F?}[;�Y�`��RO�>٨C�w��wI����@�������qU(��>���~�핻�H�m��ќB�D����XX~�Xh]�4��T?���xme��ߴ��DVx�e����w��%Z�������>[/�u�a�qX_&�BI��
Iϻ�6V\n5߹�۝�&_�h�^wv�X�N��c�l�uO�/I�ߴ��K!�S��As����47oq:�-	5�	#�G��.�j'��&�SYB����n�=Pn��v�%�%�9���+�-���#ű����?�jR�WKP�y�q�~̒M[=߷��_õ_^7w�W�r�;c$������ԟ/����y�*�k�/�ތ�Jd|L>S��fJ��y�v&c��V} p��C�4e�<����c���߷���m�M����d�3�bOrc�9]	����zøE���۫�����ˀ�$QE $���'�]L[c���ݵ�-`��f=���%�g�f��C�~7Y*�ݒ�b=��<�6�`�L�Gn������m�z|c�>��Z�U�c��ޡ/�+����JF�UrB��~V�����O�wN�������ۚ�.��F����լ���S�%$
8��������[:r��>�*���P�t�yI�ǟ�gF.頑��ӟb�b3�h��k�V��; W}��U4�V|,�|.YRLco&݀��=U�o�3����z�]��~��51j��m}2��꟯E,�]��ԝ*��������LD��*�Lzw�<y����N�g�ֻpv{��Ч�C�ۣ�ܥ�W�����H�Z5A��Xڶ�t�6}��@�v�X���]9��?J�?���s*UU'#��y�yѤ%K��o�1�^h'T�@O���m���G�tA��Wg�D	�@*vm�L��T�cԾ���c@yѐ�|9[��Td��ڐ������ەk���̙��+���V�t��������~q��a!�P�DR�[+׸jU��#�u���jѣ�Ԙ�Ъ��&�G�V����q$�;��_�bM?�~��Ru��h�oj�&C6*�/��L����P��%)�}2��<֧p1�!��e~�Ñ���u&��<�}��/f�C���U8��F:ݟEu!U����N���jn�J�%���[۬�rù>��А<��K�1>\�(��v��.���24YPE,59�Αݦ+w�����%]dݺ�&�сo3ȣ,R�<�7�;U�ѳ�}{����hxV:��C�7�~����\�@���(!�>���w/d�󝪡=���1O6�'EQ��#��oZF�p+w.Um�j�����7�ٹ�h'Z�[�@BBl[���ʐ�0"쑸���aI;;�#�������ύf}r����Q��λX�^�`|j+h\-�Wu���p�-n�>���;��(zd�����V0�l_���};Ї��J
�"M���i��'ʳ�b��?/�t�����`N����Q�.���Ln]ϤQ!�����Wi5c뚝흣��c����+��?|(�}�(�{:�����MB�IɊ�kĀ���w~�o>OF����_��1~��[��㳢U�`�£����Y/bUf;u4��nv��Yp���]�g��#0@��DĒ^�yt��a�If������Q�'����y-��`������gV?!�W�]���]������W�B��~���.1`�e�ù�Z�Iwwx��|7w:���Ɲ+�E��)�jM+�y���U�r�����ƤB%��s��s�Ӏs�%����ĳK33�x�bIff�bIff�K1$�3?�Ř�Y���ĳK33��Y�%���KbIff�%��Y���ĳK33�bY�%���%��Y��%��Y���K1$�3?�%��Y����I,���f$�fg�Y�bX�3�<ĳ3��Y�%����,Ē���%��Y���b��L��~�~�#�� � ���fO� �e3�¨����*�%R$�>�TsHiUR��v�	UEz�Z�R��A *$��$���(T�%Qym�          �   (         P             �      @ ��텶�l춏s]x�P��m�;��q��]�ĵ�^ ����*�mN^U��'s=�e��n�uw�Ƿ�V� oY7�O�����x�{kIJ�F�IR����﮽-�j�7�m�4=� =�Ͳ����;s7�M�zy��O�ok������v��w� �v�ݗm�O.��[�ݽwݯ^��3ܣ�
��r��[��}� ;�         ��^{��U��g�t��eQ��M���w;�n�v�� w)�7.�ږ;�[�ޫZ޵��ٳ��y^�uQ� 3���m���km�y���܉�UB���P|@�:>����k@}> ��}4С���j�� ��ǽ�M�hPq@z�1;� P��}� J�E>�cУ�����g���h���|@�4>JK�P����        ��4ҏ��X}i�ִ����AB��ҽ��XP�z/^ �����o0��1֚��޳��B��-�a��C^��� 8z
 P�3�s�g��ܠ�}	$(�z5�|�]�j����w������ ���s;w�}x��9��0��m�y��Z�\��oZ�T7��v�273�վ�v[��xq��w^{w�}�z��|O](��@J�)Ax         7^�_OMo�{����y��dzw:��{:ͳ�y��A+�� 3p�w�G�MJ��ޔ�3^�ݵ�}�{����[=� =��5뼷^mvWNx���΂}��{��h�w�^�AW;� ���������H{=���w����-�!G�q���5L�x ��jvם��=��ݵVn���{m�U�wy��{v���EQUR��}| �      �>�����5�Q��G��sۯ;t�m��{�[��ܭ� =��RǼ�H�cZ���{m���۞<{�y_\=^�����Q�� w{=)һ˾��m����ƻ����	$(��]뻹W�>�l�/���|���:u��� N�P�6�u��!B�u�믎ހ������>!��
�� �:�6�7������׽����o,P��|Ż�����w�pS��کR� ��d%)P   �<�i*�Ɉ  "~�T�
T   5O�$
T�� ���JT��j~��?��k��ڱ{������|V��֯�1�go//&}��Eg��  �}���_�I$�"6!$�P�!8I$������I%��I$�DA�I(Q���^���_��g���o��H��,��q%�v�v�s�ô��a�Wm�S-t�@��a��D�k��1i!5b�e���A�~�[AV���i�4���ʄM��@���ލÔ����E��ʽ�x��dkѥ�0	ueS�N��]<��դ!W&��s��C.ݰ�k�Tn7���;��P�V�!��ߚT�-������ʳw�7F'
�[�a�*�R��p�Ek��*�lJ�0��g�|[W��۹r�]
�#H�y/j^�xtPC4b�`�̱���/f��K������{�!VH)XL%/[O&��w1S$��ew����j��p㊰`�;��ͼo2$#��Hw�W��mR)@�F).����*�`���kɧ�,1u�X�L	���ͱc
���b�j��
7B�m��b�N���t�ܨ���Ⱦ��7"�-TX$߮�˕��`�����
�XTr
eMj�����'m"������w+B�+5-q��Ͷ2���{ؙy�K��0Ƀ�/d-�]Y2�X����!�]ԣ�ڕ�5!�%�<˳4�	��9u��dktI�F60aь<ī~V�x���Yx���I�XNӦ�۶�Z$̙��{m��0 ��BV��Zy�������u=�B�͠�x�U'iY6$z«���责��K��s$�3p�n����I�R�E��Xd�s^�l�)�Ee ��Œ��+,��,=���i�5%��Z���:�p��.�����U��6���ݐ]B�V��=��ͷ�齦^���;M	��q�G�<����Uhۗ���	P���E�pk*L�[R�kqӡ6�Wc\lvi��
K�YV�\p3V�a5�GBT	�y{��EZS͔��5@~��#K���I�A�6��U5�Vm���W{.6A�*mfO��L{VB�+�JU�������C�D2
Y��[zD��X-��qӛy����`k��z��e7�b��ɠ��
X���;�X�w!f��Y���i����fV-c6"���I�K�5�},�ӕ��4T�]ʑ-{7K��O�F���w�F���:I%�Q�̶�X��� �W���u�l������َ���x �bݸ�#�������y�VU'�B��[OFJ%���2�LnS���|�]�Wq�4V분�+���trnXĎb�r��	��l@c#N��dO9>�J��O�e���n�Ut2j*����!k�ȕ�)]��-;��j��%�oZp���СD0��%�7%�[T�h�Y��D��ض�=�!��4�4M����a�k�60��,f
h��е,Ve�z� �W�)�W�i��f,.d�cA�������9�dug ����,2�v�T$���<%%F�*�qo�K�]Js3'�7o�Q<yxP4/8�-8�mb���l�y�kB��O��H�U����i�J�E{Mk�/:*8T�l��Pq\9�l��Ԏ`$\6 Ɍd��x4ef�yn,f��dL�3���3h*0�f�hЦ� [�-f�Yc@�SMwCʫ�6ml�!��h�*ܢ$I*7^�Ҹ��+Ե��;�^X���۳y�9�4���[y-�a�YPې��v5�ХR�ג�e��0�ךی����V����FY�а�X�NĒ^]���j-�U#ְm�56[�۽��n�R�)i�&�,;����N!f��ٔ�������My1^�J��e����.;p\F�8,��V�r��˖�����s&Q�F�4��Z{��H�{�D$<��Y�e����xL�S��Rm�n�p(��x6]�f����Ae��(ۗE}��(+±:ݖ�N�V\��-�vw0}`�i��CX�,�fi�҄W)DN�+*���ak�CF@�#F^R�q���X;a�(�h�4�d�y�W8)��65eRh[�����c�hǀhvD!�+5+���(2�j�+N�J�Bn�s���m/�[J�۴lL��n�B�����4V� �z�#S⣧��6+�Q����ۼ[�H��0�ӫ�M�IAe,F�ge)a,b=4v�M�Ϯ�+��%��^��K~��ouqÌE3U��\Q�RĻ�`��D�D�*�7!w��S�nUoԄ�"���Iw&�kv��2����� R��կ�D�9@rZ�f�&������T�J��٠UH�3h����PO��ś���g�9�B���K��mj�����v�^�C����А�#	��.�r���D�C-��Z��lޡ9�dc\�^��S�BC܍����/P��� �qvb����u��j�#EXS7�3e�7�����_"kSwr�Z�!t�!T��bKN�.#��(VB�:{�����i���?<�IT	��_U6��2v��w�o/�U��9Yz.�9Y@����Z<@J43x�oV���
d���_��������B�(\#H�:D_=�o	�H!V���v�#*aF�Y�j�7Y�:ꀣΟQ�U,�i��|X��%�N�n�%���p�Pıs(ի3�f���V4Ή6Y+1�)�w�ƪ�h����:ng�O�y{q�3���լ��خ���Zo�-,�C��4n��PE]{�i�B��6K&ܩ8�捜��beCQ@zM�0-��܍ �y��r'V�յ�d�M��7Y�MiU�9�U6��U3l���K�/f����¦VԷG31���%@dz�����w��xX��1�eJӛN�b��6r��/�ЬH4F<Up
@K6�se����KA�EJY)�wQ1�Hi�5 �(�p�s s�1
H��^�댍w�Mfw�*â�9q^��̳�����MՌ�y�ˍ]��/k6T�F�MS�*0̽�mn��h2֬�I6]U:7T�Zܨ�c�,�"֬v1X���M�z�%�Z㡪h[��Z���p��X,+� �"��H�76�Ħ]ֶ��`�1b�Q����n�^��e��efM��ѫ�*O���1�V��OZV"�,z+s�Y����qF&L�CDX��W�q���1�c���X�#�^��]٘V�SM�LLsn�U���ͻ4�`_���\l��!��ө4��l?d�4�J��]�)S�u�����a×P?���Q�5f�$��W6��^�S(/�%]Ի_[@d��уFV����n@:�]�5���M�FV�f�VY��bfgѐ�9�k���{)ۭ5R�)�N��NͭO`�^3�g�Wb�(t���ha�f�y'i::k�ޔ��9�1c��X�]��ZՋr��z�
{J��e��S��f\�i�ڒ^Ҡ&��7��cjX�57
�*�������Ck 4�"&5a����en������j�8m:4�y.�r��yr��Ѥv��d3����vQ݆��C.*Xn�ӬBk�vNn�QL��(Yn�1屆`��1f�+6�Vr�Ť�݊!���[#�)�^����x(�Zv��9-=�*VlRЫt�	��["i�u���ؗ5jٷ�T$mT/:f�re;Ɔ7@h&�`ԭ3��*"Q�:��1�3NP�xաN�i�܉ḑ���[���De��r��1�6e�)b����I���N�)n�?hT4:;F��`���4E�#�ݹ�¢�e5�f�"��+s� b�)��6O�X��2���"��չR�pL퓖�1�ZF��.�:�ه 2k�
����! YIY(��yYs$��d��L���a�t�e�ʽ��j�5����v@������=yX�,0�^i&-�A���#{��E$���V+��+���#�o�̌jI�BÛ��䶛Y��l��yI����g%'�n��U�]A9h�^��E��AsE�O�-U��V.�{-�K~�h���67m8�M 1Vŋ!�7/ag.��*��I�H�-����ie����3^�]IZ��Ks]��`�L0$m�YzX�������KkkD����t�<�
6�PƯq�ʬN&⬖FP����ܽ��6[�"��Gf�$EB3�와����X�#)%Y��V�1�6�T�7��ة�A��,-,��h��'JȨV_�7l��I�Ɋa*C����nT:(��k����r�oP���j`��q��\(c:�d�A�ё�(=ҕ��U�5����d�����{���F��i��������է���:�<�i�����h4xeZ����-DAV�oB����{
	�M�:�S�D!;���Ǌ�Y�L�5�1�+1sc�Z�N
SX��\yI��Fk�Ugv����׺� K��(�������d����]m�L��I�
����C6�#��b��:�D���� ӭ+YJ�Sl� В�f�L��&\r����/6��Y���i�#�-��Bx�m�RT ��*sfԅ[�x���m�TK�{����Y.l��]:h����2�)�lXn*���j��V�^�Bj�sס8�R�dVo�0i+h�>�ʹ�+�������,�NI%�Q Y��f�`�3$h�%��t`����cJ�ڕz-µJ�]bß
cN^C�GSr�d����2�+%XS3$�$�U)*ǁ����P/�[�)2��L\��V�CAD�"���ۺ���Xwl��91۸V� �)U���g2�&���h=�nLٲe���ºcce7I)�`-%��I�cV�Ot��(�B7q3[��M����j���7�]U��q�@��[vE˒�]�{��`(�e�T�m?�%���R���Z��t�5�H��C���cjR@�n*�A��՗GV���c�m�d$h��Xf�n������OLV2�3�V�lE�-VT���D�v�f��Z�	b�����k5�ne��(�'/tF�J�l�:��p(�f�fJ�E<�h=9s~k�Y&�q�T�[�;fL�탭GV՚G�Ħ
ASie�jCB��u)D7(�I(Xo�i2��0�'VQô�Yl�l�夞# ���ݍ�l�t�Y����c�,��� գ��ZXAp���GP�݌�I��f��Ϋ�iC��fSe\tP�fѡ��\]�܃+u�v�}�gb����Vnt��M`5�n�+#��Y9d�3PZTû��֫�ք�є�5�Y�7Y����R}�h�浶ƴT.m1��#�F�6^���&�-M�m�n�^n=�jD�XV�c (f%%TƮ��b Q���sN<kmK͵5�H�@��]�QG�leђ���ܓN��S�u}#KrMËc/�Լ�8��p�+�^Ym���{ oXB��{n�)jc��ܴ(a�X���T��l�oNP3�c�Zv����E�t*�t�.ۉ,�:ą4�ɍSXy�
EF"n�!
-��佽dSA�;$ͥ�77,k!Z]�r�	d8U�wa�v%�5��ب��e��ZCН2me̖#���ӿ:��,�)�pH��)��1E��\��l#��Uk&Dt�U%k���W�=�Bq�����;ӛ�k)F��Y&D��X�%�óvlm�z�F62:���TЂ*WW��Gs(S�s�kZ��r�kU<���(Ս�����zU�WL<�v�l�I�â�M!i�15Rb���e��B�։��34���l.���N�dZzȺ�j�ދ�,7��X�خ���!Bг�n����#NR�L���6D1�+u���X�����	�r��r�VѴY�Ϭ�G���և�Y���CVɨ�S��bFr�z�e�tk:��fl�"��Rj����IT�Aq�I��b�u�V<2�Ti�v��g����V�q1���b�M���?������.��6�-���KF�cp�s�W�����h�Yj��6c$lj$��_��t_m�I�O!�2���NK\ZTəkZ��X�,e5�!�1�JAl�k(�r���B�V*�/Pm���%%vq�u.�r�2�ܺ�<cZ��u�uZC�ëY�9����%��Z�up؍kG6����Q�:��y��T1�h�f�W����F��	V���4�[D��n�6]�S.k;�L���mۺ��lmk��d�d�xF0����I��i�,�$�B��*T/0�z�\փ���5!f�m�63뽉�xM�
�ǀh*����G0�1��e�-�J�+�M
A�Y�m��nS]#PH&a��p:�ͳ4D���yj�Cv�ȋ0+���<q]�D^6�#�\�LK�͍2�E]�|�r��*�@�x�Y�8����v��I��M�!1Yr=A��T�`�;�2X�nn�o%M���FLqYz�^!�]gQqث��|�$�}�gƖZRVո�L�*޼R�.[qJ�e
@�77�u�û{8m��j���k�RO��f&os7.��G]fyj�4�62�I�� �"�A0x��b�������i�����P���0���ڧ˲Z5�Tܶ�5Ԡt87FI{������-�w��i�����S�^,�M��J���������$�cA!��&K�o0P�nƃ�cK)A�X4Fa�t���H3{�,i��죆)Ou��ukU�WF���r�m[��MQ'oj�m���@f�:�m��^��h��MK(޺ߖvA�w��6�L�lL�D7y�PB�e�1YŮ���t�lOVȅ����؊|-ah5�ڽ����L*=��#KE���˴W� �\p�-�s,�g7m�{y�!��p�#���P��n"�2,ru�b��h��_�t��!���x�'�;�Jt�
%���*mi�V��-4���6�+����]%_rb�Pб���-���;H�F�4/����i��[-d�q�,���?r9"�=K*��LL�MUi�Ţ���t\����0�y�Pj��'1V:�(wG�m��������*����v��j�iV��e\T��v^YZ�Y�)@P��MNԬ�UUUT����T�m�`���m[j�K�[m�UU*�T��l�����̨[j�t��هI5*ݶ���-N�Z����J�]X��4­R�l�E�6���Z]k�� ��g�FR^>>>���$\ם�5���X�ӭv���kytoxA�]s�c��N6�.$F�b\s�8���;mFe'���^��m�������C3�٩��G�{���3�v�dY޳�����7s��c57;��'���[�O�|g�kt<��bf�.������S�e;c.5n�<�Ns���u��؏=n[r�X�b���A���6cra�'&�#b���J{{����;-=���ͱ�k��K��n�dMZ�e����z6�f�`�.8�ݻ�]��۵�]�s�F����9q[ce��vn�9�ᳶ��|������G���S/��i���M��65�/8\�8���1y�M��
۶b�9O)���Y��Vz�q�up�e�cuu
Sʶ�bv&LS��l=n�9h{H�y�p�n^�����N�@�f������\�=�5۪�]��{
��}]w�Z�e�fEw]��O!��g�[�6�m�bK�ݱ�ez���{gtI��v��'cvG#u�9#AZ.�Óƫ�@m�{i�����K�ut���I��d݄�է��t���>�3���]n���r������oM3��n��z^ht�^N^�5�]�k`v�{q0wD�g���0=�mf�k��&�'b�/U��rv۳�g������y��]ѝ��v��ڄdI6(�o8�k^���PNn��W��<�-��tÔћ�[���[��i�b�N�`���6:��G�m��6�]��n7�Mp��z٢��¦��7*��ێq��{@��l7m'v� 㱣�/&{ ��5�ָ�a*��Fc<g�pt��B�ל���+{v�KW,m��T8����'ۮܟ)�.n^o瓸lv�n���5љ��v�=��9��v6�6�F}�
cVpj<ln9D���Zժ�]�q�`��cov롷%���-�q�y�f9���]��z
q�a�b�qQ��ۂ�9y��(�(������8���Q1�8^�wE�m?}����Z�_v�\�T;�x5�;9�"�����b;v�i8�v�tr��ܜR�Ƶ�;��vf�u=ʺB�ݍ���Z�[�����Ɏ�Ϯ��\M�K\!Ko\��W�nNf��Sb�7l'd(�hW:�M�Ba��]%��k�v��ضsM�p��cOq��o������`C��跇� ��`����a����Oru�n������:�Wv��m\��V��ݺyn㵣D����Y�v�s6�	R6�iǡE�(�t�8Ơje�"5���㹢<�<��q���h��z�6����}�����f+c��Dхn�;s�k�۴vus܉ =��rRu�5��q5�׭�H�����Pӕ��x�n4���BC˧d�p��v�����v�zG��E�Ɖ�;o]5��LY�9wv�#��F��\ޯ:U�n2[���к����ݩ�ӑc��v��a����p�ps�5�{���{N�8q�`��
^�;bQM�;=�؇�#����x}f�eF�W]ΐ�s���y멶��a�lIdV��^s�\^ø��������yn�]��U��r��g�7nb�Ƿnѷg��ظ���s:729�Ty�v�Żͫrs��C�RC�w<e�v˃A�c`���V{n���Nu,j�zz�y���aXx�Q�[!n��2�C�:�ЛKj�`�����ܘ7�ہԝX�;���\\�: .���z�x��J|i^M�^��OV�d������kq�W[d��CV�n�:6=:�6�m�ny��(b��kGhR�홥Y�%�ffF�ۏ"@���B�ɷN�lr��'=�����Y��0)qͫZON��j��xֺ�Z;�P>��m���1��y�w���k!����Q">��7eƸ��{�sq���';���m�� x���kA��b�.��9e˭�v��J4�ҙ��v�6�v���ݢ��r��y^�,������*���g8���Mb_n�^���ܤsM����WD�M�o���=v6�cq6t�v�1�/��9�7'�;=�v����'O�
��pp7�����zѝ�]�\zmq�hծ��Ka��l�&1�9<�aY���Pd�\�����gkpXc\�g��ֶ9-�;d�5z�����Jy[�=�������M���{V)���޵�-�M������Ά���Ύ9��<m�L��$	���wG�^�v:���[���F�V�ﯻ�w��{'�g�Ӊ�x�S5qyꝓF�4�F񝍆�L��Ns�B(�n����ga�!i.9'��$�N;z�r�[.㳹�]�1��<d2{0�9&��n���r��LW��F�j�6�m��b%�ϵM˹+���0�1��|��:��S�w��t\r�c�on��u���S��Y�ۘ����g��{ﯢv�{v��8cE�%C'[���7��y��I�,{unv6wG\'o+�o[�^#&]����p�q�6Q��$$�g�X˧ր����]��h�K2G������m���P���[�nN�v�=����n��� ���l����\��]�:N(O1H1f���>��IlN��we�x37f�Tk����Ŵkg&6��jN�;\�g�f�X���M�8��#��%�p����huƹ�cq
�S�s��i��u�6�lbz郔�pr�pv�vs���h7;��(����=��izp3t���A��h���:ڎ�ݼ������Ӷ�k�c%n��t�I5�8��r�cm��:Lb�/c�y59�{u�]�4<�%�pe6ۧ�����L���.:��!��:|v�z�!���9����� Nn9�듵�;��G������u��]U�of�z���v���7d�3�����1��9P�5��57[w!Sg4l���ۏuŏ<��ۧs��N7\b����WE펮���q���-�ܾn;��n5��:��!��8L�cX�b�]�l(����g�V6�s�j���a\�m=n9.G���8�����M�u�0
����lǉ�	�&;;rQY;Y�����$��ȫ�M���-�3����N*�k*��in�̇-���&�vٺ���Q^W����-x�v��܍먺,�!�΋�dW�g�I�ۏ�v�M�]�v#ar�cm�m�hݹ��y��%`��И�d�����Hh�\�i�1�� �ۇ��k�i�Ń�]�co�j�vU�x���y���A�s�]ֻ��;Wm#�X�=��f��p�7�����m�G�G����v�.z܉EUŋc��ku��Nx�룹x�����=��&h�s��۞NNNɈ�;o&�2�kv��+�$H<g���ݼ�ƈ��s��GXy
�n6�q��k�n>~���W(`�9:����fv8��)<�u���g[�qoZ���qq�^��lg�u�}���wf8Aۜ7g�ʴXu��=N�j{n�	̸�9��vƬ:bQ��NSظf�F��v��r��;A���bz��S�݂y�Pun�����#׷el�01[�!��{MӯtWmnSc��A�xǃ����=X�.���4�t���x|����ꌦ쳠�۸�=L��p�`����ɺY�3�,�j�˞Ӆ�T*nn��\dv�}kb�m�c�L�[����]��lΐь�.���a�W����^�Og�����ch���ucDw8���Uꛡ���}�}�g�ǈ8��S[=^��9ch2v2#b��v�8���g'q�=Wt<���;��
��.ld㶹�;)�U�ʆ<[R�Gˍ���M+݋�+p����4��ĩ'Grk�yi�9蛢�a�r�n���OO��n7r�+�z�]>��贼�r��O8+n��]ئo""���GJM��Z���:沙��sgl�L�S�Y��ƵѠ����枳I`.V}��q�Mc���W��Ln����{ք+�e�t�no^�B}N�q�=d�9�v3�z�mڲ��i{Y�X�q��m���r������w�"AZ�L�b�܊��x�u%m�iH���k&ghtY�۵�h:�;�dc�n�[	1�tR�쥝��Q۪{)n��;n�Y^m��;�ݍ�ǃ�0>�nn-���V�-�\秱�,�w[c��ۗ���^�oh���[5�E�3��3��q��|�n��6�gv�ҰSw[/^�	���9\3���M��<�ӶU�Ė<���쾽�͊7/�;̆�"�9�8��絛��ۧG��ڎ����:�.��{3@9��㧮���:듨��a�NM�l��f5&�ێ�q��gm��{���#��[�N^�#ۓ������S�玬5�m�ONݼ��ء�A筻q{M���J�����X������r����d���6�ۧl�*����7X�Z�Llwon��uÇ7<�%�}��f�ɹ�ݺ����8�G��X�)n�(yu�n�L��s�(h��u[�=�t}�1's�.�g���`yܦے[�� ����9�8�ֆ,5�nݠ��E:��61r�I��S�*��#�� �݌v�]���ׯmIeCme6N�v25�Ѽ��˶�2q��<�;nbIsg��0V\��t�=rt8v����pQ���9�k�m��[86g`��b7/�$�ƃy�0M�6u9�ϵ��q�C�_V�]�ή��Ɨ�'���g�sո0�b��=�݀z�<�;=��lgm������L�x��XU<�7D�n^2���nv �i]�uu���_f�v�����6�����<
^۬�2�){���T��@���ĺ�F�c���7g��JLuôa���~??cg��u�ۛ8�ü�s�[&�WN�{mt��8���ݥ:^=Om��퉦T;���d��M����ô/u�3裐ݷkvv��W�r��*k�T$�JD/�Qj%�Q
"G�BI$�D@�D�K9����t��k�y��P%����P.Ǭ���i7gZ2��Su�..�hݷ�\�;n��>��	���Y�a��:��Ǜ<�ma�Wm��37!����N,u��dì"n�i�=gp�c��t�r3<����؝v�+��v[�.�r�\��i�^�*�cFÓ��g�V���x�Nwg����gƧ�����gC������Id^ϱ��ִ���'uv�d�����8%�j����qy8�u�c�v�����*��Z6Nf+e6�-$m�];A�4�����9\)��6z;H������-�zn�����qr*aVw*������N��9,q�n����[vGs�g�b���q�]j��/^=�0�f(��鈷0��z�m��v�@>q�=�6�In�oS^=>cn�g��qx8zS�6Iݰ�w!��.#W��xݢ5(WO7���'�ס�n6y��ݺms���8�9�x���nv�G8#��X�\��ra�;;Yw]��I{:����dn��w�X�^��šS��N�b�H귞JZ��9��6�3���u=U�|�X���ܻvq�v�q��c<��\�w^�b^o;����N�-��g�'=($��9�)�-L.�멻s۳��cvyz�S�m��kn�u����cu`�<qطl6۫v�Ok��;v�UnE��lq��痗��r�-�bm��\!��c�f�����4�s6�n\��fv�f71��H<i�\�b�d��=k(��ت�Bc%������n\8خ���<���Up=4C�ۮ�=���vMN�ݧp[���^g��#�.5�f�c�	��ݻbK� @��vmm����ӽiۇ��{tmy����
��8��4F{Vw���A�ݯmŹE�d�8�K��3��}�-oF���X�n�94��x���z�ӷ^��\-�[v�zr>Hy㭗S�s�/�.95��¼]k��m��gf��w[i93��v�)���e��x6�N�@IHU1T�IV�D(���b"!B
!BJB���D(Q �%	D%�"D(H!BP�%�$�%�B�﻽������m��stj�n44��[���"��o`��jc�7���9;s�C�d��k�V�NX��5ڣ�2l�z�ݘu�S���>�S�8u9Mp�Z��&N�\u�=]���h+vܽ^�rr��A��Gꓳ�<x��kl���$읤�z�w]��{]���g�Cש��h
�<����utjy���Ϸ[Z�9��\s�7Z�v�{���»!��콗{<l;۳���.��p��q�.=�����`���m���������"��3R��6�p.��i�ۜ��1������k�0�^�����H�X4�`4Pd�̰��s�kf�J+Ƴ�T���ه��@>����%�����t�w�;e8�|#�H(ZTM$I%X�v�M�e��Tb����V{�h62�W����ת_��v{eo�M���R��6�<��M|i:b�h��~m���w+:�[�>�;���1�li����$�S׷$f�'^��r���PO�.�&ŕ0\wjQ=tJT����f{�u�����W�8Y^�,w�A<�1����W��lsP���m���_C��m4�\W�_ۇ��w��JRtu�7]cC�ɡ�^ۺ���Aϒc�����:����(���`�J���r�W��W�EZG�z�t\��t��I�nf�*����2�kYxfu�l�;<F�@���m17&�o��kŴeX��V@�̝��:���K��J�	��̬�9TB@)�q̰BD��ѷ�43t��_b�n���隌���-���Z�Y���aH�J�~���זְ(���2g���	��L~�GN�ٲ@lw<�@�'F�ʐ��0�D�A�o��Y�w/L�^����9���M��[�z^o\��MfO~'u-o��FfQ�s��,�g}�E$	��HK*�Ǉ��ͬw�d;9�ޫt� ��s��]h�)�~u"�[�Q�wd+FJ���z'g:N��fx��1&
[@:	�`������d����i��Ă���{:F�fD*�����.M�G6��X��JU�B$��v�:��љ�W]Y�qt����Zvv�nΣJ����9�*8-`6,0r%=�a朐v��MiaI��Cx���l��r�>��wq)"���Z�Mۥ���v��{'	1fg{ty�k&���7�,��?3L��2�	���s�����7L��#�R����d}�3Q�l�J��}3�wI.6}z ��پܽ�Iu�#e/_�j13L$
HM������l���G?"I�3yA��s1�|�X~�(ߣ����v���p����/��g�Ӆ�[��V@�E���7����M�;�qلh�m�(s���`�*��vA�=⬶M��c0�	�[6��D���6�U���78%�$��RIa����J�Wi6����G�It�#��y�%%�V	� R�U߲B�]���6h|��%�c�����n9��e���{�q}+aY��Ƚa�>t���l��j-���L5wIZMR��Ž*����kR�e��-b��*��s��3�K�v��r�v��N�R^x��nJW�BM�v���(W��Yia���x�mX�<n:U����n�:`+�et��P���`�=N�xG�.8?��jQF��Pj� ���'iF�B�p/F��$�@��~*�wM����t�Ytl�A����/5��@ֲ���-w	�̏��-�i��n���m�/�c��(mח]�`��(�y���w�~��Ǔ���i��p9tt�]�+s\}�td�) 崶[Ns���ت�ÊZ'1�t��X���O[R��X˞3n���i}���	o
��ƶ���lk]q}c@��K�
�f�nGY��uFm�gl��(W7s
�X��V�Nn�rݭ��	��I�w���T��� �=���R:�Mﱙ��M��|q�]�._Q2ͮ�x��ku�{Tmx����=a�/��	��;w��G�Di��'l��W�_|��nޫ`�][qC���Չ�m��K9�c�TD��dvY�������1~��6$fbF�K�3�Lt�*u��v�����n��������]����z�s�j�@�2h�H� M6jS/A��Z&�{����z�fz��ZQ3�70	�@�T���v��t>�s^L���'F������ 
�Y&��ft܅��p)���h�%���8;����h���Y�<�$!A�Q��G��#Ӟ^�"�g�QJ�hQ0.�.~	oC����y9c�R�v���ބ����3�ŕ�m��B�l[�3/_�5к�ACc�� �QD�5�	5��e�H?>\��E*ES
��Jb�Y	�C����en�+�r��%�\=���@H"btw��ܓ&^Z��|Y����/���.Ƈ*����-��Y|�ze!I^.�B,�36Qs7�^1��$�V���v��n�{ޠ �p��za^��y^��.x#gs;Ζ�ǎ�&���'�7\J�=q���y�	7�.v�P����;f�b֋���n4���G]lVh�냋7���>æ(��<�����fz�quˢB�z Ovz��h�3�p���D�\Ba����p=�rGm���m�];�Dݭ�T/����Ŵ��v�W]c�v������+���u4�h<��9�gj ���{!��V,=�qy�ۂD�;,d5[���5O��H3O�p~����܊;�)��o��t�x���Q��R�Wa5����r�ֹq�m5�U`HШv�A�$�GM�ķ۹����|]<�:�Q�XN�%�u�該����}a��RT��&���]4���k%�6�	U�Y*ҿkn�Ɇ�x���{���۫����G���ń�[�����L�� ͼ8�5ݦ�4�S��*i�g���F?e�.ߋ)�y���7�ͷn��zW���i����ޡ�L�a��g��*��^H�"�RA�i6ۙ�>�����O�ny�^�� ���Vc�N�0p&uF�\�u�΢҆O+���I�Z�:�,�r|7`:�=�ٺ�n�	n�rH�uź'���ۢ�;<k���mv+�&5��pDj����.��yX�#[g��ըѵ�6��=�.�1P�؇�S�[2��i��W��u��_c*I
O�u��·�򖙟G�p�͜�:7':����U�nff��w�m�q�laԞݛ��:#|U[휃�SU�yi�:��C�'%ٳQ)}�o���u�����<�~����n7���\]wK�ץ�������$c��QoKs���p+<�n����.V�F&=M�_�sF�Z��?'!��h��aH���Uh2Z�])5���7�&jI���pi�\�v�:�c�~�
�^l~z���BZT�}�<x�q�XMudkV�v8;�c-N���A�u�Z��Hp6B����]������3t{&:�6;�Y5�xy*C�Z��<�7����5=�]�n�S�p���]��ּ�#�t�l]i�9�ギs�Q�n;��$�[�-�U��m�7���k�9��^=eoWL�Ta㜋��!/wz��-[!ޙ��N�
Uj��U�q����׍�<����X����[���{�h��|3wX��S����Z��;=�����AX�{�n4(-��B>	4K-"�R�z���C=z�ڭ'y�iζ�B@uՎ�� �y��Kt����*dgJ�Q���^*���Pmּ%-�º��h�l�v�!m0���'���QW��vhmx��t���7���3����)Yg��m�	ҳ����r Β�T�ʃ�o؄wf��rew{*T)��n��[,<�`���۲�7)Otk@ځ���*9�*�M��%�k7�\AL��_���Fֵ�){vY�����^��F��'�?=�4�w-7�&�q���/1��|C�6��^�����fC;��nf��rS㨺�'��jwg�]���߇t�im���'�ɏ�~\�-u^ӓ��$�mi�w�R�Uoe�޴G3K���.<�H$���B�*�zbG��_��Z�]����Fn����d�̇D���~��q����o�zV�{V���"�|�/H*�
�4�e�kqNA"�n>N�<kۛǵ뵔�2N��{�W��1y-s�����WA�N��d����T��{�ky*xނn�{e�l��w����_`δ4'�T���V�v�^gE`�A�[_U��&��9hȪI�c�=����w��_h.�7�w����k�C98j�b�p��v�r�^��a�9]�������6��~��`* 2��cV?[���yn�O=�������&�x��h� T���@fK��m�s�&��H|�{Qk=&�sz�y�>�jҶ�E���1��]�9���� ��8ּ���m/��,6�%�SjW��b1�3"K8�g��TM%]���<��"�ko��X��<G_cU��7ΛP#j��E!F�Q(�4	����D�un7o,'K�x&i�w�\�r�hU�펺�V#����Y[zb�?BXj�\� �USm�V��I������r�2���YD�o?u�o�B�G�ç��`.v�g�dNF�[Uz�ЈRʅrPL��f��ŕ�E��v���J]p��)R�����Snc>�c]晚滬���]��l�耊�[8e�Z��/a�M4�*���ޞ:�evz<�:x81>W����ڭy��~�О�GO�MF9�ǖH�7{�s
��)��qW-�}hy�Ǹ�L�u��m�_B&O!a�+j��񗰘+�u��=/@��r�!;6�.�GN͍�A�Tus�&��O�b�vg��`��qx�������ַv:�vn>v�^��N�۵��d\�ͨ�\B�7bb9y�뗺tr�#�:�tk��7Zs��N�I��2:�E�0z˯/6���'t(��9� 1��N㱭��%����YD��nwC��A�����sx.w���1
c���)��㭹�Cn�OhX5p�Uv�&��;Lq�!or�b�r��Nյtl�;����.��\��x�Y����?f1l�3�F*Y�����ӆ�ڵɻ���T�5�_��fb� 8S�Y�joڅqƨ��V��8���>��P�^���W��r̲�j�y��gb��)i��)���z~
���=GX�[���2�ln֣��i�iW�u�bc+f�NȍncX�	�W.1��em�ח�ϊ�Pb�TJIf�s۟joc�������Kα<��Se%S=�n#�$��/vK=|���v�,��)@QR�+�RW����:�L�Қs��3~�^�Ɇ{3�$�D+�Qc��jI�p�逰���g��ZvA�u,@y�n��n���uG�1*ŋ�[�b��mkV�-�@�Y޽@d�v3o���q�H$�p�ȏ2��n-�=��mԧ<�S�T&�_�����)�<#2ܧ��"�����D�*���7w]s��]�k�̧�:��ˋ��Rrb�V��b�4�fB�9)�&�G.���n�	nU�nk�/��l�ʱ�7�lVqK�P��cr��3�8��8B��T啍�^��b��̃Y�]��,��+6P>���c��[7�G��1{9�r�̆D荣�J�^qa۽&���R�|��ݜ3�I%��r�"�j��=t���UH�p��i��z�7w��o�,9��E�.�F��[���L����g�W_��Mfc����P����DQ�E����uUl�.A͝{���i�3���`�������o��,���.��G-��߶�~�(����!�I���;�D�wh��Z�Ν��M՛��hF�q��C�m�#֮8y���[��}m���r47���{u�o�
^�=ZOr@=�?U2{�6�7"�	m�J��]|���,��U�աρ�ۄ����	��`��<�B
�˕|�]���#��C��J�9t���4�:yn@�q��;e���U_�%5�@̽Ǯv��"������[U��-���&G�C4+�"Z/ʲb�.U���(����҉)T���*�G+rBM^7d��:W�R���q��� �!��+ u��8h0��+Xϕ���&R{�x����Z�U�b	A/4�y�J�ڎ��V����|Iy�0mie���;ŧ�X���˜�w�W!��ٽ�I"=�l�i�r�.�(�f���:��ʤ���S���t��[� d�m�l�B�P�su`Of<�%�g0�+L�D4��wS��y�4O�:Bb�oQ�n,[��Q�B�b�"
d5)�N���M�J��J��^d�-��E��F
}e��1��m�@Ү�)8K�æ��[��v���{�������ħ*&��8{������qΙ.Tb*��L��kX�gr��R���Q��f�ы�J�y*%�e̓���8���d�T�����n���s&p�)�vj�վ�:u��s���ˢ0����={�#��w�Y���$�<���$3�lϲ!�Ef��Z�2d��ƻ,y���X�4�Z�HY�R��0��e���G4\+p=�$�si�὿m��݊՛��ә;�������{�Ejԃ4��7����7	q�Af�%̂�3�,�ඳ"�u�5v�gw�'e�ڔ{�{sp.ySd�'w\�e��]���`�ۍ]XkJp)/�^�ş�:T����W%6�."�x,��>Hvt�j^����B�,�	u���#HY�Aޣ�ut�a�]�1'��Gta�@�7*��v���}��?qV|hH��pǃ����v��ږ���2A*�"A�	�y���<Q�]�L{�d�d.�l�SNm�Е����O2�'����=|9�a�]��`�l�<��J%���pL�2ַ���tw9�.�>>CB�%*TgC�R �^|�>�af��>��`��P�Eg͔S ��(�!X=�d�N��:���1u�Ϯl쵷��f��-v�v��U�J�n{Q���ٿ���)���E�0��U�o�r��C-z����2R��3�v��G1����5��_vt�z�u�t~a���l�Њ��Z5�σ4�-t̩)�V>7���7b�Ub�󨻄�;���mK=��_kS��tdхX�4�m�߂Ve[\A
�b�"�e��k�-�+Fպ�w����4���z��Z���K\�^=�G#ھ*�=Uc�����.,��̮F��f���W���(1�%6Y�s��3�eDvt�ދח���w7��� ���[�5��1�V��"��Iŵ��'^E���n|<g^dg������+�p�)隬��q4:+9�QUy��s���"�	�ڲB�-d�a�ֱ�u˕�+��h{ �*z�Z���ox�M�|��y�{ �>�B���2t^#��m6L�E�i��.��َI;�ݭ�+kv7m!�� �W4]��Ο;�f�*�l��i�+��m��!��z����7&'C�z<9�>�a�j��ś���v�p]e� d��5�8��;*�|q�K����v��+�8�����oXy�<v��#�ڀ���������E��<�/����%����kz3�uv�=ܙ�M1ެ�5U���;W�D�@y.����ԉ�o3��Z4� M�,Mo��"<��^�H�N���{����M��7M$��z)Ǌ18�\�>��pe'|Ѷ�(1��L��x;p*ܱE�cK� kģ��f��|e�N�\U:䦗w���YW��<[�et�R�������Oy��*�4:�3^��٘N�v4����rn\/7�谫�7��@�v 	�3J�e;��� o:�6��B�	ܱFj8X��\7���9W3f}+a;S���T;m�jd�t��Xyޣ�ݞx9'�.\�s�
b�d�a�mڶ�u�Ca8,�`y\.�.�U�bŝ�؟[��;`s�7��N�B:��ssݸ����l8�c���%�ڹ�1y�kh�-��CXw];mTb��n��K�-�}�����Ã���t=�Z�p�Jn8�ƭ��m�s��M���i����
�s�痶-m6�uwCvn�긣A�e��;��Sc\����E��:�}���9M��Qy�x��a�@�ax�`�}:m_��*F(��?�7fS
�W��F�76��z"���ssr��cyò	�h�A��{C����Qy�Ů��'M���,eI�b�-�&�'�ڏZmq�mO[��ޜ���y�g �p}��n��v5k��eoN�L^��8�lp2�um�|.�������.�]wx�ք�q3�o��>�a8���vKے���9e�.�OgKB�b>�+�`�[��Y����j�('��U�!�&ĳL� ث9�=~Ձ�������"~B	�t��n��y�^>y�zd�cYK�NOV�zo^z�_u��e�Œ~1�L?&�Dz���B�4x(&��hOg~�������2�skX5���-�>0��۪㵀y��^ދ^�t��9�"���cM���5R�hq�f�e$h�5�t���B�W�U�d��۟k��W�U�+�mD|i�T�Ɇ�m*�,rq�| �'���3��Q�����~׾e�e�Ue�"r�d�B��:y7��r�+w7�./�L�-B�1��k�F�r�[���[Գ>��$�d���xMȷǼ�Z�\���ֹ2^K�>�ʆ��2�L�N�$Jcvs��P�a�Zt���C�yx�
��u�^�2���+ZkRO6X���c�٥޼�dEM��Q�KV��e����Ȼ��"��t�2�9����{;r\����fP���v�d�9�x��y��z!=��  @�������l�7�I|�2���I���HB�4�LLV,k4�%l%��{h5��4���>��-t��	��J�V��+
�ތV��k�R7.�[;V���f8�m�Y�ט<h�E4�>6mݫl���7=��:h�3���-����*�����M�V�Ǣwm����t���!��LH�)6�G*j�o�5�[�I�4�mKZV^�����;�U�Zj4>��Y&Y�5yͺ�zjh�X�׍���A:@r�Z�x��̲�|gfR��O��Γ��u�l�_U$�XP��4�I�M�쓅��\�����f��W�o.�2�}���1iZ*�1-5�><�4&�&gH��Uk=A��/��+.t�V�f�]`��:�$$)m&�a�l�+�W���t/.5?@Λת"C�v�A�������z���X
aQ��η��n��}�r��_���m� -�� L�Ka���j��~��zo���������	wB��/���Rf��Б�m��w��9�s���e�^�~��}��P�1����u����ҥ!�l�w7x��p.Il��9�{zn��̷�k������EDUhJ����aD|J<IҞ!^��!�(�K��jkF������SQ0���m�],!�����hl m_�б�g�":���u��63����ip*���}�3]���Nv���G7Z�Y~�[+�z0��g��)�cx	�Z��
��~��kqE\J�Ϡ-KV������oWo��ff[��V�@�ti���2���ɱE�6�/@#7�<��"+�ɐ,b���*j�[�l�Gc�x�x����z7嵨;3w8�d����l]s:5]����Ҳ%�tYK2v�uqn[�i��򖆇�/���m^(���˚�f�Q�]���tu����&�%z�II.�l���F��������O�4�6�"�Z�y�����ir���Z��,We1�[�*ˎ�8�H��ٰ�:	���u[��f�q)ۜ�ĉڹ��x7e��݉��qr��mC�������/�Ӟ�����TE��}e�_�w��2�P/΃8��^r�x'���+|0�j�넣�ך�#3�s.�.�5r�<��.�r�^hi��/�Fq-ep8�7����>�N��A�OY�ܨ��}���[�B�Aa��xr�-3����aD.�*�6�b�+:��.�ɓBÀ���:���)(/F�Y��ʏ�0�����6Z�`)�zf���4n��u<h`\lU��z`T<^��.��|+��(����X�����ۻ��,�U8Q��)�~���y�z����Ɗ-�d^��_��[��C&׫��]w|n���<���\�d�������}�Ȯ�"Q����/fS��ͣ�.Iw��J�x���ۀ��]C��=9��(�Oo��$�:����\�G��7�7$r5hՎ�Z�H�ե�f���Ɓ��vݎ�u�]���׭�����k�톗g��ث��Z��;�o�w���f��L%���؇j��pWGbM�-�v��ݜ�.�Nu�=���Gm�h�^H�h����Fu��kjӡչ�6h��؃���;�ʺ��8í�L�C��s�A�p��)�\nVv@�/R��]ݻ0jt��Uv��ݹ���ד���~����G�YaT=v[�س
���� y���ݭ�ك�bDnj���rf��/�u�C��fͤ�3Y�m�S�����{d��{ͣ�R����W'����<�"����z�yڶ�w���'uz������V@Y��{e֧9p̠mSZ���^��d�v�ܺ�˶������
�e:��P���f��������4�ř�R����E���+�ɩӹ׌I��*�)�60�u�������;��}��$�1N�ٝo�&����N��J��}�'%�j��{E�ɝ��-�ǒ��RD�4䒐��s�g�<�-md�i�z3�Z˓s7q�?�zE�Sjs�LRݰ��M2�-�z��{S3��R���[u����>ti�^3s�yݝ���v7B\�k�g��(:x��t���5e�F�C�We�On59*�f>M�Q1��]�yh#j����.�}ad�D
5�>/����[�l�aOqG%��r��[k!-�{�r����]量>�;�����,wƝ]jD�j>YN��2����\�׀M:c��u5X&R��gV8h�ʸ���̈nr炥���<c̨�M��t�}��ᛄ߷�<8n�0�e(�7��to]]��fo,�|�� �&i�ӵt�Ƭ���d
�>v̛w�����4�Y���2��u4s��Z{Qx"���*��z�;u���}~��o�Q`Thk"��m  >�2�@Ц�GP�����]�S��T��A�@	m�9��2�<=jU��sj�yL�E��_x<���L����y�5~Qλ6У]ylMc���I�k~�suKYk�����&�U�H��U��' nn�۞�)��r[�Ԯx�"T�u���y�]��me�jM�ݪ��R/��<�Y(�k=Y.݅��>r���U��4���lZ��s�1w:�=����nz�	۔����ᡌ���8����V(��*b�����#�.��~N?0sp��q $(b@eJ˂I\|,J��I�K�лZ�;X�;!�a�Q��+sD'J�7��Sn����gg4�W|���2��� `���ܰjs�4�Eʯ��Jr�'�z�L6������}����Ե3��x��^Q�w�M�(�#aI]��P������^d�GhM������)S��qׯz6���#�i"�xƇ�D9�S����{�!�4�_U� "�n���S�X��t�y�yb�%w�q]#� �C��Gg�m�c��1�ʍBV�U�=�b��l�ӡ@gT���O`�v�p���7V�&��x���t�5���[�n���,Kw���?���W�����iU���^�[
�+��^�����j�1��)6���u��>:)+	N뼶�[-qL7A=w����[�S�n�ܣ<�3R����GR^!��t
�W���jť���u�)�	�J���Ƶ9j�n���8f�=�=�~��^��s _=�A�Y_,�sW%�Ow&r���^�gԆ�I0-&�e�W[��+�F^tɡ�	hn����~�!�z�쏈E�ú���������|�>��R��Cz�r���E��읭ʵ�h�&|��;w���B����G,M����8y-�q����a]���Ϡy�k:�`L����݇��}�AY]j�j,qh�P��O���XWn����S7E�v�ɎVy��vF�y�TDu%�V�u�C���^x�j����cv07�tM4���Rt��L���y\]���˩6Af��:��%m��>*���vZ�stm^����\^���q륗r�a�ʀ���K=�^N_�� �f9��𕽝�3[!� �]4)�_���")��s��X�7jO��K�I�~;u�8<{׹��m{,�{i���-�;,Q�Qx{kv�?^p6��˴��Mu&Kcd�Zr�;��2��6�Ao;���8r�z�GY{��>�b즁�#w�Gz�r%�xx��fЬ�RJ�nK^]��o	���<C���qU�{ƹ�$�"����h�`.S�[O3�$O�/a�я�.�5h}n��e��Q�qGU�W�����=f�ڛ(�K���Gt��z��N��{q�G��f���Me�7)f�C>��N����?(�KywZ玳�J.�)��<�s����,<Η��T� �D��o��f���_g'��f�#��`��N���R��	v�U<��V��@A�H�.�T�GZ{ێ۝#5���AlĲ>���;M�<:�f*�U4-�IU+�Zxf�7r�	�$�G��&��˩�!�~�0b�}x�
G�؊t�;84C�6tȂК��t�歵r��v]#6��;{��\�m�өu"�yԷ{���u$]�*�=훙;R�ǚQ `Y�b<˰��Θ��g`:;zk�¦H.�6���7V��i�^����q\���;BЩ;6��_˓X�[x��$�
���&�z�t����د��ۃ-%f�I�5�F	K6owX51��\���ewbЮ-��/o7�@wv;p�n��J�4l��{��S8�[S�KX2ƽ�A��W}r�l��j�#KR�$ݥsw�*�=��Ӯ���)��έ3Z�6�5��+-e}e�@a��d����3�G:��kK��Qu�q��k.����S����v6j3S>�\����f̒��V�+���p�uJt(����X�q㭡|��m�R���|��1s����K��%�ͽ|���EaD2�.���0q���<0G�.��!�E�PGx1^���J��0Puj�'D�Q�Z����ҭ��I�0<��v��cT�4A8vnVY`��K��yHvH��r�Fh��;��}|;�a�Q��O�ٰ��Of�ao#��_�6A���n�zUZ7��\�HYJ n�k�* �b��;b�2�eZ����[9Z܎uc���<�녪=��&3�u�=�z�(�����kb��0�6����s�鷣�� �,��c�q��\ܮ㱺y�p�8ͱX�a�;'[�gu۶���4�ݝ��1����`ɺ��k���7BvC�QPrT�pv�6_^��k�>�mRv'Og;6R��j-���������9<�\���uO����g�.g�R��7h�n�/[�9�'o=���q���.������9:ڶ픭��{���}��l=q�&4n�'%�lu�V8��h�a�F�mu|�8��؛���Y6�[r��I�ٻ��Ў�T�[í��n��;=�:�:���ѻ��u�;n��z��l=1G��km�H�\\�P���`{��{=ն㾒�cm��`���������3���ȷ�d�O�m'v��5������f��7��]pɱ��.�;�僞�J�7��sp͞L礎�D�8����c%xH��M���:�m7�t�;O=eG�=��S �f�\p�wt[v�	�q�)�g�����_h�݀���v�-�����m�Z��`��.����;'�t����g��#qC]�=%mu
W���a�7[�q��uݴܻ�n���7!���q���.����S[<��qԼ��p�d�z���Nt�h�Хd(�/=v��Ӻw:�n�)e3�s��r]�Ɨe�*3��F���קi�w��qJV�,���dB�Rm=:�v���C���-�^ܓ��dL��y��[7[��������`��+T덛�N�&�%7.�Ɖ8�]��Pct����<ݤ8-�6)U2t�Ð7��vu�\�d�g�W�m�<=ezl��C�eς���w�`��t!�e����v�g=���N٭χm���:��ںxk`�X5k\�Lx�;x��k����q�q�#��N%"���=�����Ε�0���=�ۅg����w�vn;��9�z�ؕH��4�/k���x�m�4p�dٸ.ū�p�z���9F����e�g��Q;�˱����b�o�/�iw5��8�	�m���v�./H�B�-�����Ч���rq��o[��y3c�C�%����P�n[�a3<G��B�;zrt���&{��xمɷ7t��{yvOl퍙��ۍ��k��� �h���{f�v;��Wa5�L�K:��z���p�;�W=d��؃WY�����G=[�M��S"�n���R@����vcj����v����e�%�Rj`�ٗ<]Zf�a�t�h�r)x��^g��;ypg,}�Hl���h(��C��uu���L�9�(͐_hM�f_��sw�xп,S��i�#%O?S�}ť�p�gM�E��)]![���E �
a�>T�=.{�ǽ��iY�TF%�sDi�*�6���9P�m����� �M �*dR��A���W�U�{������9v%c�[�ed�/T��u�P�~PMn�����׹�;7�eҠ�hU"-���P���~
��&j���<<L
�]7=�P�&�v�ەR���S��B"|��*ku{��B��Θ��am�N�Ѯr<tq�����7<�Y�ηE2�ɐ�\R�~�q��+JG�pz�ܮp��,�fs��	)'����-��\(�%8j��i�����)y5�F��*^���s���z�3J�E$���"z��bcB�s=sf�r����a����zI4cWeK��.�j�=fm�\�����[8�cp��}����nĳ\}�ໍŏ��;�)��bz,[�0�`/j�%Y�A��s��aM���M,��V�����J����i�ږ&�+P�@TUI4����*��s���Ȳ��y�X��n�*��5�]�#Ѭs�q�=yX5�^K�,�+�B�vY�vY�}�ui�?a�V	Ջ_GJ1C}e�$��p����]��A�}ڝǲ�zw-G������)-"����S�l�Oo�/�mz5W�}Y\,����Gk�P����i&e�_�X��I����L�W���k��ã��Ok�5+Ͳ��[su����X�f�㮬�(`x`.��l�]��|3$z���+i[�Ȭ��@G-�T֬;��M�Mc�@7�u�rc��u�FAie���<@D��;bL�0e�ƺ$}���m�T<���^�4$V�y��-ͺ��(,L�[u���!�����.������7B�f�JңT��ҡ~�TW�AM�r/�od�W�)ڟ ����3cڋ���>B���]v�8+�S��V�,��U���W���f��7��'P|����������圮b�Z�^�jx	�,�yN2oi�����z G�s�jM|>i�H4����[W�}��m�i��N�z�x�W�sgb�(���|���p;��^*&����V8,)�+�p,�L=`�Z���e$��<6������fp�GVk��FOu�1��Y���7t�弋��5.�c�<���jO��e�~:V+#������������Yb�����`{!F�V�+;�=bXe��pbg��0&�^y��̘�4��W�Xzog�mE���7�U;�3ҕ��@8"Lh����-^�3���x�<�8*F�&� 㧤%]��M��t���W�e0Ebwٕ�:7a�Id�ٜ�!�ږzo�=�^G�vxt�d$�����m:���kL��\���\���8[~�ۡK��=G�)�6��I��V`�K�u��c�.��H]UR)U�[t�"{B��p��S9��g��ky�}�2/*�oy�¡۴��V&�( �LǸZ��6���1�e�FS���}�32��P�e]�uy1X����䵷�j�9�M=�% �ak#o�v�`�6�f�o�A��x����ۑ�F��\���ˡ�F�m�T�l[�볼e��^���>s1��J93G���Ƕ��˺,L�Z�P������1���T�إ��{��*���<t���/'/��M��Z��&�M�it�%rn�X$9��nt�;�ZԿ������-Nu]z��xgZ3I�&b���}����Z�3�.{=��1Z4���A�����7�;߼|�O�	evS������9d�Ukn�>BlCٕ �.�y,+�����z���N���ik�5,�[��3=4���mЂ����<߽������ز��jy�>=!��JRmƘ���a������Tܛ������	��R�H�A�%+Ȫ����*_�	7�q��7<�;T��.��V%���y�G>6F����ͬ��f��X�"VE��IJ4�jt����1d9�=���9���L�l=�%*Mx���0��v�>@����S��S�e��7�6�tVNSH���6��AF��) _=]{��!n՝$����d�R�޹�
i��tպ���;&nC�˖�q!�
��6�o�?��,KF��p����:���=�]��7Ey�]nR�=\Ї�n�;�j$�0:�DC١^���=���`���Z�R�	);bz+,��u6�s]�瓳d����:��v�Z����v������ovv�gm�w�r�T� ���c=R	���՗������˛t�W���p��)�v���ɹG���@<����Xs�=�.�ܛ���s��pspi�=r�I���y����6:���^������"������mP-���}��Ǯen�y-�S+ŷ.��a�T�I%"�����q�-A3�=���~����R��R��-qbv�~��Հׇ���Wd��Xw% �ߕ�5� �۸o�1�,-Z~�H]���=%�\`-�\4�PQ(��H�of��{�ڸ���#�Zv�y��9E%Ԏ�^���9��/��-�����rުu�<n�0R�IN�-j�-��"ѽ=O����K˱��q�Fy���
eZ�����c}��7U��E{�tK�,�g$��k�P�J�4�`&��DW�b	���{��i�B�\���v�ɬ�v�U1�������o�ԭ)����D��7�o}�:H�!��$���t����L11�lu��/l�=_�k���F�N�@��VT �N���ǩ���o�������/8SQT|��հ׆W#V�\��]@�h�2��[�O�����+�JڜR�H�$@��W���OԽǳ2ȇf�YU�_���5��j	J�n�A�T��%X����Z�i����ѽٓ���6��(�v7��O�ڊ�Z{Y�m�Mɰ�0d�8�-ySs.tu%`�o�Y��� 쏮�b<Ή��o��8��]��j��L��ۊ�ߑ���	("��VH:���9A��aZ5u�nT�j����`{^}\��8o�q���͊�����{yn��[~k�m�zׂV��'7��� }j5�U�Ž��vk��l<?x�\�,k.�� S8o�<<sf2�� �4�_��*�6Z(�o׾.�7�U���zG--�}/T����<wό��_����wl忶⡜��b��w����=u�y]#�,�s�u�z�s��
�g*] /0�O��N(G��	մ�����ff}nۮ�"��dk*��D���;�Ӧ�C޶��;�kv���l^;�7��Z�i�=�5�X��u@���!A]��'6��&}�bfs�J�#;V��5�2�n��X^��������V�l.d>&ys��o5����էo(<�Y��,�H�i:�|y"����ͭ�{o��;��gN�l�	��<�vc�`��ӓX�L�ڽN�K7x�E�㳭7�f��{�	Ն�gw&y�֦T��}�)�8���b��V�1����֝7�uJX�cr+�ڵ��慴��KE��a[^��8�e&����e�A.�ye9[�h�I/�u�*�����t�A�S̗a̘j���H��ꅶ���(:�.zc��j3��X�;]��y�T@��0�k)�J��vA<��eq�;����ry�����SቻeCn*�Q����U�*#�g�!.J�;h�:w-�Xɋ���e��
jFm���8wj{ڋg�y��Hc<k��@���v��8(���U�-�B�זH�wū5�/!e�>e,sᒭ�Mڲ����r�wZ�6v�.b&s�o1D<��E��r�K�8��������� �mH���<�$)*�)�~0�|�܇|q�+�V���?"|��z�xY̊�dZ�q���W|ߞ�o2���Ǥ�좨�GP  �٬�f,��~:z%�h3L��l[Z&-�5��S�u��Kb�i���zR᪥�T\��6iďL����˩|�<8o_I�J��5L�1f���-����q�t�N�����{Rz����!���ݘ��M�O�S�i ��t�����׵�
aҼ�|�{n���B.��u�c��'�iA���i�>�f�ͩaaZo���M`V��[��<=D+�7�R��l� ����aHw8���-9A�p�z�,�ĭ��dj�
���m���YF�.>�ierL��1��rlٌ1W���Q���y���'��m�g���`]�MK���-U�J�-��9�W�����٤Mϗ�^{7��<Z�I﷤0����3۽�<���;heߥ5efv�N�o��2��m�����(TJm]����#�B��1Y�͊��VN���[l`ۊ��!Xؚ���~{[�26_n��}�	Z�7:���ߪj�)!Wh�!��<�+P��j�n���8&�8��1E�U��e�e�z��;����k�u�ӓ�V��SZ�a���C�m2�Q)�9z�粚�s�-�*����3]���H̲��{ǲ����[���(�@�0)�����zB�XN;�v7���@�����,�;ji\�G0֋�^���;�(�r�I#\͗ه��g[)6��,���Ň=�;��{s�m���/
n���n����<�kBV�ruۡ��A$rS��f���ݐ9'Vy�Q��޻Z9��C���ͨ����5˹���cc��#��	����a�wQu�����u���=��I>�9��D��9�N�ڧL����ς:�v��\�7�ڱ��k�2�]���]�1�U����툁Ⱥ��m�(*���H�6��m��$��2l�k�	�wV+o=\v\�u���L�A�`P-�;+�w��}?n�g}��QA��x^�Ǐm�]7�mY���a�2���O�PQ���Z|e�ᬟ@�%� -��3;w�/֫���~^��b��k�U��O�b�D�#�xYCͅ��v��u�gV��S�ME�"�L ,5L&��Ej�� �{ژ����FB�锔֛��r��$�ۨ��x�`"�"B�;��<�Nf��)��rI�i2	j� 4������~�GY�pў��n�b��UK�=w�ORU���~|�����5gj�݃(}Dۇtf��Lz^�w�gƌ����[j�y]�V�̫�w�kITe .�p� �����+ְ�J�M���[�Y˪T�\`�;r����W��\t'ꊣx�V*���[�?�?}۬��j��7#dۓ/'^��;���\Hp�Q5A8�T����Nx)��{_����oM��wE�Ĭ��������9˸Ԭm�$��{�L�����D�Q�
�$����,Ph=��w�@�������m�'gS��u�颕�ZTX��9���
��	�;jz%Ubrɗ[�K��JF^n���~���)��V��{ha��O��^{j�|p�����4<�X�ץ� ��D3°�B���,$��{o�m�2���yI/��Vk�V�c,Ύ�p#��f���-lY8�F¡�-h���dV|�O��*+��i�Ulg��P�b��{�n/si�RH�x�g���=��SŶ�ݏ�%D�C�^�I���=������O�"��Sb�Rt�g/\��x��9��z߅z�zY	��l>�S��B]�$(o��/4�D'����j�?VU��ŀ%/6���~D- � �"�A�Rl�b��;.�Nv����]̝�����8�իn7)+�՝���F���rc���ׯLM�/����o���]��]Jf����0�����C��c���îfXm�MWt���lB�9eZ�奫s�fvw�Qm�&�cF���B��ҏ���e\���.�����:z���Y�݄�2/��e�w�S N�`��v�DW�)s.Y��̮*#�z5��5���jX�\�k븻��{��f��-��9�ݠ�O]�����T���7&�#�Q����rz���&\��4�|��Uaoy�����ELku����2݅J��X���㦴�̝A�:�^��9��%ˆR�B����M˻f�a#����s�J�5����Wy-����;�C�
3�9��DŘ����RYڋ~Q�ҕ[7g;8@�@j����NP)]ؑ2x��z��!	����cBGx���3XE�M��6��:\wůMT����m��s*�
��4.�.�s1�ڂ�e�[���t�DaY(����b�%�J�yrv��v
;�N��J*Lz��yJ�2����>���q�>E�=b� &b�ү�%���1��RC�,��k��v���m�U76�LWX|0;�{��=�Ye龵2`��d�Λ]�� �����ࡽ���tw.���g�jXٻ3�i��J�oT\��:I�mN��u1Ccr�;bf]���|�J��XU��9�'�4�F��F-u+"Kٝ�o�C�r�a8\2��� HiAU{��sf\�2�n��J�US��M�T���ϫf㇣r8YY7�݊	�r��KnZ�h�1L��Ɋ��6--�	�q��`���!`�����Ja�u:������KX��Ŏ��w{�S�׫�狸��G��$#�G���&���w���ӫWl�5i�#q�t�\&��q1&օYGo4��G�ot�j�q���E��ۊ���Ŀ�P�J����5��_���1:U9�&f��b���׾�����6��v�G�l��T+_w�����-Xx@Ţ�q�s�i���=���=P�ey��4�w�w�k�&v�ä�=�k���Д�$���r��OҢ59VI^ҭ���,�斃�)���{����]z�L*�\��SƘ��U��wᬥ�*��V����"f�J�\��Dw�s�<Jw�LR �!H�[/�}�n�C��5º=k.ƙ��iB�������\����RїvG�;��+�:�:���c��^P�����v��
��b�S��/1-!���
L�� �cN\���Z\��Z�:.
��c±w����t�8������v��/�|{�)}��.{�.]�|w%�g��K��x��/ڱvT��#®��o��ր�1c�M<Eܹj�uE���0TB�D�R'.9���k�y�ٝF����럅!��<aM4!s�}�μ�+�N:*#����������.�o�K��\rB���!p��1���p���������������_y�k8��M[-�ͭ4>	iT�C��*�?���Hຈ�}p��S�~��Zľ3-��N�ɗ%�W>+<W��%��'8s�V�_8��L<���M+�/����8'-.��Q����/���*�آ��BT��h�\(F���[��w/J[Ĭ_q���;ϖ.��K�x�����E�oخ��+���²��0�=���xEGP�Wn$���}����k&�ڝ]Ni�D��t!�=	�B\@r����>�9�J��f�8oC�X��{;�������(�^�aN��mW��4� �RAO�1}?ef0�BC��� �@��j�5K!}ֺtV�)i��O��}�����O|-�Ef�
����i�kk��V_۸��#/�T-3�C�^��h,��4��{6���dX��ƕ�j,�e��<��֕�M"H�jDGED'�o���_�����85G��ji(�ue��c��{^XX<�+�z�L���<s�^Mr�˪:�B<D�|"Z�`������g�mGƻ�Q�%[��?9e�騡9��%G��n8N�~u�Y�⴯�w�N���+9-*:/�f����ປ���{�İ�|ՊȮ}����ĝV[i���\iV��~´5�����ت��h;��X����D�^ʅ6�����.x�2Z���DcZH��0�/r~��v� ��0h��R�!e����иtV ��n>v窸Ĵ�C�����9�U��C�J�$��]M���$_��qg�f�%|*�bL�SO�>s��p��9P��f���_��yup������_H�i�o
��ŖES�so�k�p��:��M<>Q�=`��/��;��K�	U���}*� �E�����81���;Ց&!:tD�mU;��Z�>}�މi_	ӅG����Es3��IX�`��o��~�!9������k�Y���(K�[���)ODP��9����
Nc�����R���߾�Z�4N\{�)�>��2>0S�۹:���ϫ��9���7��5bd�Y(�oϟ&�I���,Zc�+A�︳
��ĳ����*R���<��د2ڧ�����T��s�c3��+t���N�"�b�T�ׂ�d�W��H5�! CQK��y𙲭���n�7�.��T{1����n[��D�)ZD��7����uk����kymqz�q亰���.�V�v�t�y�}���T�)ӌqVM�����}�۶���e-�\�cnn2�c�FK`sc��91���2zƗ�K]�7]s�v Ӵ�ݸ�"!�/��:qGU��q���,h�E�vZ�;l�k�map`�wj�5�	�^fr�y\=u�Ϸ��rg-����ܝ����=e�W>�v�d�j7��`t������G`Y�N��n��d�0���W������I���
��*�8�'-�8�J"�"L�P��ޖ���I1nԫ#��b�D����+�a�'�f�{;��nv�<.����X�f9�]�o�i��W�),V}�a	��/�:��jZ��֖3F+:a�X[��%��g㿞h��~�����+#�+��v��iX���ۚ�:oD��S
��YM&�9�)k߾v��:�C��"\�r�A�}Ϸ�H�@K�8����S��j�z|~�X�Kڼ5�y��Ub���%���|sݕ�\���E	��_Q���}�D��]"J���ϝ�K���Ib@yS~��'��T�ƫq�WL+Ss����篆cR��)��n�Z�i�H�s3���ӄJ�d�R&9���_����	Zu�VҜ��-��������y������x���;���ɵ�8B�$雓�-돲~�m++\*/�VB�?��~��J���"ݒ+n�fh�cwޢ�.2v�9�X��1Â^��w@���`�Z��ϰ����e.�\�
�.z�5��~�J�y�"��Q*���q������~���!R��Di��TK�X.��+K�H�Q^k��*��b�'>w4�uM*�
���Hf`�}bd_�/�k%�����;�i����1�������s.󹽱�C"U��5M�:�%�v�Լ�4=�^�ƀ���TP��_q\-#E$/r�8!������4��D,��߾�H��s����fr���O=�g��H����W��=��p���6$]�ʶ�SbS�:���-�*�SC�1i#��Y
��5K bSO���j��*"������c�Z�����LlW����F�:�[��v��or��Dn�m��8,'P�䨵��"�tԢ��\�L���{w9�@Idd��E�*���B����K��iʉ��-6(���k�)2@Tw��qX�8B��,���ش�M�7���hp�
���cͿߧ��ԣC�:I s=��[�p5~%�'%�D�w��G��KJ�s>����zp�)9��XF9�����]�zaab>����������RB�I#�smZN��/�=�"�S2&Qe���\P��wܨVBdtW���Hv[TQQ55Oat��T|Q#E}���ҿI��L��#e��`��$��V��sk����%��G%��cg�*�5M�h���D�����/w�,�>}��ZB��\�"���!V�{��r:�P�1P捅��)D,���Rv�
O}�r��p�Ť}�o�W����äe�r���Vϱg�����v'˚0�gu��|��u:B���
����ͫ�"лy0���#���~���S�a0�� t�,���N�m�U��ry�;=pQ�c�x��K-M���}1�`N�KM���=�=�:;�z>��iO3n��.��`�x@P�R]�}�b�޵҅�S��H��Ea��NV�7"���wr��^�&F�ک��p��ÿ������H!Ø��!O���-~}O�$� u�`K�m~����vC����Ş0]�.���]N�W7���_/%��R�;��Ӑ����X+,@����
k�wŋ�gdI�*�ò�_ۉ���w���s��z<O �������,.ZԴы��YBVy���qV�ﾛTh��K�R�#���`�'�(Q��DַϿj���)rZ�_<!�Wf������"-�g˯�}���	�-�>��0.d'�N���h�9���Y�h�A[�;�����{�}�8��;��F<���dIb�ӷ���f�����Z8t����QmI�h"�xn������bQ�7��y�{��u�M�]�z]uZ��[�| 	��V1XǟV�ű��!Q"��,�=뇼��Yn����p�|��5۸�yWj�]sx�o��[8����@}��M�G}�r~��X�*���/��yT�TD��H�#k�R���ң�#��"�(Z�Ϳ��m����}Xss�U� ��*(^�����̟�ߧ�k��O�ýk��#��P�;��+]#�.�謒��FI�ܣ��켗�nآS��2�iò	��\i���G�K�u��<s����ѯd�;@��������iDy�~�K�b��"{���,�Ҥy?vn�"A��Q
���V�ks;^��ϼ�t��R�0���]#o���v�L�4�Y��ȡY�wꃹ/�eH��M��@�R%�i�TG��^o�p��lR��5J�²����Y�5\)͘�:0������?��+���2J�e+"�S�QS�k�f׳J%v��=]���KH�g��*QB��$*\���4�E��j����x���qã�b�0G�>����L�����Ж�RTa�o~��-�NWA�x���]��g Vm�
���!9��6�8�����(�:.C����_�I,-�O��ŷ���>����p�]�K��͡8�R����X��M8�r%�jm�sd_����*y)t����\Ɠ����E>I@P�ұ*�<�w���şk�zuՊ�ע1ͼ���'!st.��W��΃bl�:��4�@^$E�[�lN;�-����#Rߐ���s��}�h���:+�p�����	ls*�R��W-!�9KV<!���
��}�^y�5�dY(�
_�Х ���l*��F�>c�� ���O�~昖gj��i?u������U����j�f��BnKZ��KH�L�z^��fE��o6�cP�v�[H7d%��a=����m�Y�-��(�j#p�������x�U,N��q.���j?��CQ����NB�fʲ�iy<�Ȳϭ�;��<Kz�[��,Z&}�J�Mg_��qZ^�T��B�K��ϸ���8$�B�F_yɵ���:��ۅ$b�znI��eJ����p������CF��,0���13��3���T�,\� �I�D�����{�ⅽk�J$�$J��!�{�q��B�~���H{r�!���ӫ��u��U��o����v�}�����s�pT�e�k��3�*�Ȱ֕$}�Z�Kq$|)c��5X��}���\���/�}6��_Y����k�Mߦ0�r�'�l�ж��X��B����ۍ�BÎ��?���o_�=�ҖJ����Q--�y���7��Jc�p�{�\-ˎ�3���
���E�&�+>9������U���v�B��R��d��{�h���L�hX<\��bG�����YS�;$,���V/�0��5���,�]�z��)'��S�j���bM8'��aB��cK��}3�+��Agb�l���w��ӱ4��]�߽��.��8�P��5d�Y"Y����|-�ڡ�J���E}�}V�GD�fW�i`S�H�r󸵟1����'9S�F�D�\p��G#�+|�H�(]�v��,�G����pf�����>�~!�^o,������[HԾ���Fym�a���v�v�ܷ�PH����9[S�jDA�26�rq�v��� ul��u���ɷj�.x�u��0H�S"��c�;Ǟ�k{�h�wkEj����6{�yt�w6��Z+K�]m�gv�Tsm��n0�8���8a6sr�Ǡ8Ÿ���(y�t��ۍI��v�pւ�uF�<n�!v؉�+�oKc2G[�qq�v�ܝ�.s�|ۭ�O�ʽ.��.�ۗ�sv�Zo��^l��O���^J�ƙ���O���.�N(��p�M^�dG	���g�Ed_6V�Qdh������|���{����T��E���p�d*"E��iiP-p��P��<)_�?�_~���U]l��%�{١n-&�1+>$�%�L|�UЁh��,D��}���,�
�On֜�U�K��}Ʋ�}x#@�p�5��K��ر"^�B�>��,OZx׸�!~��n����:��W)X?}PF��������疀��椕X�V���ܿV�H���~
���j�iC̘�y��+�yQ�38��\9޹�������
ut_�-�?s>w���³�`}��qb�|ޔs���}ʐ�E�4��>�K0�z�ͦӔ-TMJ%ML���8G�e��-��-�|�xF�ę����w���<O
P?��"ڱ2=y�&ԊK���@%uЙ_r���XtJK����/�缟��%��s^&F�$A�e8r��8(ֿz�����p�V������ڮ4E��%&%:�s�}8�Aç�S|b"�T,�˷�����9�k�Y�6��}�ZY�q��#s7�tpC| V_�P�܈��9
ѳ�>-w޺�t^mS�����p�e�|�����rj����sv/>�%��f�{pvנ\b֋݇�#����k���k��z�\���.m���D���!XŞ�e��|k��ӂ�]y�D�JDk�W���q��ofq�=����z�9���^{ߝ�3�;��t�I����Q�D*��:d- �s
�X���[�>:�33B�	U.j�dp㍺��.�
Z�����od��*�W��>�!L��
Q���=U5wl�}���+���Wlpc4����6�Bk�[�8%_QcYj����˷�sa�R����O�xc���+}��/ݛXE��	�O�I��]k��o��8<s���l�*�2i8_O�j�k��F�H��_��Nֺ�X����9D�\\h�P�1RJ)m���B崂���K̿��4VpVX�ێ��W~�]��~.9�B�9����p[{G]>���Q�9��kL��w�1����f@V/w��p���ٺ>Zx��jC�-k߾����p������>�Oג���󯱜ޥ'�Y}�l�Z)"E�9��"�>��>�U��U�Ņ�
��%�LW���N$�vB=�W�T�T@U~?��C���O
���Z���K�>�GE�\tUn:.�U�|�`�IT���<�\�R��\Y$�����:�Fw%pAb��]�㾵���>��Ly�y����CX>�5�a��m_D{&���z���,��m�oOO
z~�S���;�>�C'pg������v֜����M���쑶��K]�LnǞn۷kC�tr՞�{e}�!7�E̹$KY��f}���9q�5����8i�>�eN�QB��c�5W_r�X-�b�%�����J�[;E�p����|��.�I�"�>�qZz����P��<�4L��<���aP��[+����Z�U�
?�{k���ؖ�ϋ���\mw+�˽�ML	?9�f�eo�F}�ip�C��p�RD�͉��V|\I��ﲼF��bdN��O��.���#'�PuJW@*�8��
�pP�R��Z[u>�*ƴL��^��p]9	�RX��֋L�n�ﳝ.��#�ڿ�JUZ�y�t���RGRL!�vi�#�����^u���<�z�EF��l���G�i�w���<���b��y������C��8��f�˥|ʿ-5�
ΉUO���Z|t�;�`��)�n��k�i+̚0��}�]�mm������R(V*�-X����)n$Ro�������_S����-זVں	x�qZi�B�|xU3�*���SN�8��o��g���=�^ͭ,�!:jH�j�lGҪy�8-߷ŧ�@8���%�ɵ�)�*Ra5.jh�ZGE$pTxJ��̞�3�VF��*$�^��ɅB��r�|��>�ֻ�g'�XE����!W���k�ڹ�8X)e9#m�j�����'g��g2pJ�`�D)���������e��qq���8�^*Ůrq\h�Λ��`:�J�]yٸʉ���1Uv�g��.��RPĉs�G|��J���t���]LQ_SR P��J��w��kVH#�����1i��u���Q�}esh\8��Ț�Ͼ�C�Bv���3f(���_��u���t�r.���h�p�-%bt�D�33F%���^�0䵢��JD����鑢��GFtu�up��
Hb��6�8�x\�V�\��r\�$L��G;�>�_�щ}l�Y%�� Kܿ���s���7�l��@A�q�5�,�{N{�VªJnU��Uϗ_�k�m*���D��߮s�!h�X�b�����	�S�(ڿ�7ݘTv�7��y��6����0�Έ�{�V���	�g�H����{��+\�"P�m �i���m&z����#&�NI�.08*:Eg���qE�� �ҭ���1.<ح?1��q]�0�WZ�E�ﺮ_T��n7�X��!e��qbE};<��0�~S����������J�k������6���n�*�)��dC,EG���'UfJ�ήN��	����	��^C�aU�>�.x��ѻ�֖#\|)��EvԜ��|b��}ϥ?D�\�S*Ym�>]u��:W�k=.O���an��Y�^ݘN��g8���x}��|-��+^"x�Q�L�>��V`�z��,�8d�S�M+$��qN�H秞���|sꖄu��dXS��6�G����O~�߃�/~=��Bm�y���,�ח��ص�v��aBڇr�u�c�oj�@�g�7:��z�5=����̊EfS�,ds�y\h�5(L�WN��Ƌ��_^�K�j"Dkҙ
�S�/>v��4�5r�������i�X�
�<�]����"RB����Xدh�s���H�AD�.�l`�E
�,�<%dQ�}����g�#����͇��O�Kx`{�w�p���b�r/��ia�2�훉HL�H�L0�˶�8�~�-aB��C���|h�����i��kK����+QU%������}�]�����zӖ�>O���oȎ�e@P�$F�`���k�ظ2$�=f7�&���Œ�{�$�w�e�߸���1���8g���/��iky�r�B�3�2(�2�z&
��k��$G����-6���xi��W���/])#�}�T�^�}�q��&`�VE��N��e`��,�UƗ
*UK=ܕ���?��\�X�V�L��nl����~W���c���Ǫ}ڰ���b^9�)�,!��,,K���u��K$���Mm�ؙbA�+T�L�s�g>.E�MR�[O�0�B�S������#���p���+����{3%E�J"���\a�;,�[�ڱ#��P�ټ��Dp��Օ
�%���P���]�?x��oɗ�'enA��stu�"ϡ����?I�k�N���Ǫ���+4k̽��	d��Ds�s�v�Ve��9�A5�;����>����-ै���B��0�*���d�f�4^�����q0p��Mpm�5R����%������X���r�O�`;V��w.�oi����*�Eeܚʇ��r:��ŗ�!=����+{J�,>��\�q�]����X\��[kaWN�E&�9��J�_i�N#wa^�1=sP��M��dX�߁�F,����;v��/n͓��`rU�#U
��˙��.g��K!�����z�{i^QVejA�M�Bܦi�������V
����V���[�c.�;w�V�2r�7�]k�YJ=w��s��N)X��	H�[G��y�<�,@4������ۿ*޻�9�W���q\����:�Zt�=��V��T�n
5
.���y��ػ�Ɏ�}��B��X�V�v�:ߌ�b�B@h�y���{]�pK�28��Ng�j�)�u�7M�7�!�39t9��{-��F��P!��u2�WeM��\��Lƅz�4r��7V�)d�흎�X��Sa�lꁘ�W9l�+�y2�؍����[ئ����Wb��k+.`O�c%��w���c�kF�nӼ��%��u���'3�Y�.���rv��5���۽�n���ZC���y���ۄͫ��� ����u�F�8�dQ^g\ԪR����wԸ*8�v�8�$���%&�v�]�݊U�V	�3v�ݳ�t�-���\�S]c��S^p��g��k��z�nݙة�Ճ���ݽ�gq�k��jBĜ�/��F0c��.�ͺ�8��!�z�殺/�qd78s��{��2�ɇ��r�:�x���)��L.1��S�G���v���oG�Mat�{u�m�8㓱�Ja�n�]��!�m�e��n6�vA�܆�����Y���^'W\�Ŝ�Z��sմ�m�v_n���wn9���ۓe�1Ϟ�ɶ笧<ޓ]4s��H��5��]����kVA�n�lc��5���y�%�u������ѐ�=�� �2��{ub�x� �;�`���Y7���96�T�ss�圧�7�����R.{�r�n&|��n:�G�{5�in�����/u�9���^����N��z��9��lV�ɮ�p�RJnx�Ǎ�:_ep��m��]���snv�ŭmwd֧�;T�E�aY�\)Us�7;\ġ�$e�L��{n�f׶�n�Ѝ��d���3�n8�9�9�;8�1���(J�gY�u��qF����v��8��0
ɴ�a鵖��N�-�n휝��yx��w&n����(Nx�V�.)�N%��z�ٸ���&r���lRi�m�.20���Y��=���n�ԧMs���;�\ő;sm{U5� �\�"&���(��J�۬���:������'�����Ξ�f;h��y�!s���\y�v���ջsF]�fδ`,�c�3�n=�b����+,�5�Ϸ6�x���ż"�`�cur��	�8Z�=�$"�c�E�= M�"��ٹg��m5�^�6��嵗Tk��*w�����nqñֶ��v�%�9U��X�8��[;69��qЀ�%��+������9g�m�Kq���8�b�Mێt�lQ�5������E���H����ψ:���+�-�)��:�;��Y�çL ����Ϝ.���	��v�T�X�\�����#����i
��"�ݳtvM��wmPkmA�kH.dwd}��n��T�sĶ��wU�ѭ�^m����N�BM����.{j�9���ay.5���+Ge��v�v�q�<�a�<���\9i�XƇ]���+���n#lrtL���k9� �� �oVK��"z{s����ں1���O������&�]����u���{S��Tu8��j���N�N:벊��F1�����jQ8ۍ�:�Rݥ��#��b�,M��X�m���4m���E�.�n��O_��/��p��ً��q6Ջ�fb�����D�ǥQG�d��]g�7\���۬�}_v�塀is��X%�B�7�ߋ�ٙ�l}rC(�P�C�o�W=��+�ߔ�{�B�k�������f������ѹ6~;Yf�������^�����}L������om������e��b�v�Y�픸��wK@��-�B�YB�Xt��W� 5�j�}����.��q7�,VB�f|j�]�'/аV�l�m���f���sC�Bщa�s�ゾ8TD�RcbE5�s�}�}�s��K�e_2�ɻ���p�g������Cr�L�di߾��hSY��O��D��[1ao����wm:r�@u2��*s4bVi4�t.����zg�������/S������FE��U�X�fˉ���|-��"�%�m�I]�J}Y�p\o�E$Q�4��R������`�����zP�^�(�4�O����6�mSS��q�i/���20�Fu?�{�\!1]f��L���+�sP�/�&مί���E��
�"Z
� B����ɴ����J� RE6���s�T��s�0���$'_d�i�_uӻ����U����{N�;�[)dk��ne�n���6���l1N�X���`��-o�x���G�dP���(����kD#�"�T�H�[�7o��z�Qr�E��Y3�����:�ᓇ�*���!�P!E������oy�$��3�I�w���A���J�z��JQSU�	p\;�a��Ԡ�pж�훅��ϯ�@3��*>ȷi�����5,X�T؝��eg^ɎݽG.�MOOn�>ݬ_f��<}���0	�ڐ�񠷙m���^ף�N�I�����k�W���)(\땘�"&���*��M��<C��x���b%��"�����8��Ls�����u{��/˰�v��މ�iU69�TZ R[f��Z��l��q�[�if��jЁ�͗�g�W��SL�.ۅB�_��/��N�@����6�x���O~����lK��9K�m�4@#���H�`+��Ƭ�|��rqd��P�����{k�Y� 3�o�TE��'褕b�N�"�NS{�>}�w��d��t���
��ցӆ�˚�VBb�p���n�9P��6�L!��W�v�Y&�����Z�(��&�8�������9��e��9��i�j��������x�;)l�k�x|4����ҳ�p]�y��\�B�*�LX��4�jn��1��^��c���xՒi�a
��h����0�Z�u�$Td�
ȕ-Q" �}�Z���ѷ�_��XT2�����s�{���N6l9�m���,���iu��q��d�x����7@q�˙�)��U��Q:�_�w���\�g�
˗��v��D�r\pTY���ﺮ;�s�"X,6�+daw���W��dQw�5�|����x��&�T�n�W7��kN��iv�g��8��=@�ڠQ�ʫ%��kM*0Ji�J��̑�o����
�~{�����|��jC$�n���j�*��@�4|,�f�]{���_Hb��d�łUodUϾ�T��HW8}�]��_\�d�ď8hR/���;2���� J�o��?�U�6�~ࣣ�&����\a�^��0L�بT.h��?zmt]7�M8����<�G=������qq�ݙv�F-���G��B�"����q�I�7�e9]tv[��4�ϗ[�
r�w�����[���_�d-<�ʡ[���Ta*7�� aDx�Ɏ
w�W||�vV�_�5qn�]ڢ���V����)���\*$���ק��u����ຌ���\8g�t�,Z��D����&o']Ɩ�`*"�j��;R��g���V�m���(��V%�V��ۙ���S�����k��B��\B�b)�|.x�?�G�4�Z�Kq-=�5l�Q֭+CR��d��}xe	t�'�s�1��7��{塞�mU����<Y���.zR�}�-h����"���d�]��v��I�>oonk����i_+N/UOiS��j�����a$��5Ej��Wi�u��\�ǩ���xN�������sJܺ:MS��� �6�I�l�0��6�j�!s��U���Z#c�b������p���* 7���
��:n&���k��=������B_y��+��z٢�8s�o��|X\���Ʌ��{T�Q�\�5��宱�� �}������D,6��f8U���d`���g���*�<�6�3�IP�����X��{��_d��,��9<�i|މp���T���^��H���U�x�1x]�����ߧ���i�{-|���j����"�2j�R� 8ԝְ_[�9᥂�w߻W5�Q������hʙRMY���[ٞӅ$W��}���z���O8�.��+!H�5����4� ���s�0��3-Jқ�����tR�V��,ϗ۾�wB=?^o>��i�ĽM1H�=�yR8/�Ȍq|j���c<�+L����.��/o�όko\$�H4�&�#�g?qb[O|6Ҳ(E8���Ӊ�O��ߤO�l���k夽]�%��}ũ���e�V
�*�U��b���u3/���Q\��X�%�Ƕ�gE�*�wnW��E�������L.��P��_Yk�jF�:@M*n���Ť��f5B1����"c���� ֟3���(R/u�e���'����g>{�Y����%v�E���gyߪ�
����$�Y
��Zz!�p�&����?)��|�Y��[=�Ӫ�b�@F��N<�L���Qc��^ۧ4W��1��m����]c���FUZ���M�~��+��q����~3�;�ƴR)(�Jtp�Y߹��W���¥�"� $�@�n� U���B�>�Uw�n�up�?P��)�Jm�\ꛧ��t���p](\��VE|�+�w��R]e�0��e7��X��D��6�]�`A�Զ��VF!h������D���va1iB��d�x]�f��8M��a�L�}��3޾���fJX`�f�N}�k�p�/��L����mr~~� ����O��Q���2؉�USUV�	�����E�OZV+(�{鴳��;�bb_sg'f��Jc�ߺ�*;�
��ݑ�ӛ�|H��IBWý�_&7�O�Ʌc���TEy��w�Uǀ�<U��.�P+#�l�']���+"��ii�{#C���1w�o��r<|4y��n�>Y�\���Ɖp�ݕ��ς�8zs�W��,#�j�\�*��ھ	j��|m*���++�Q�?o��p���M薐�XL+"��&������peU�8[\%X���L��%%���W�j���.��i�Eh��<(
`����Ǩ'K�}�:Mǅ{�\<-��֛M}�ݔ������9M,�*��z�����2Oq���I���-��B!%]��[�\��e6�� ��/�g`�{/)�gB�\2P,���(���U��_5�(�v�h��߬	^S�y����qd?Tᥫ��׺���p��nM[�Z��nv�
���zx���a���tl(�u��b:s�{�-����-n�Y-�����Og��/����#�z#�:9����=s�y�z�p��;�pS��d�[tS�aw&���2���P�=�:q�9q�qWm�*�M�N�ۧ�c^B���7'^F�Õ�m��-�vxW��7Mn�s��j	�`�κ��=�e�y�������7c�+��eK��h�	���мG<� �bडP�3�֋�>���2�]->(�W�T���;���:%d)"m�u<~�����izs2�]��3�/�i�`��zF
���j���b^7�����%�y�,̙ꟶ��R���o�^}H}D|/��!w�q�g�	�����_����I"�Ֆg�13�p��og��d�D�"Eo�jď�RU4�\5�n��9j���qw'�'�r�����B���n�6'����dR�s56�0��%a��5��s�ެ��t���%�B�Y���qB��L+!�Kћ��׫�d��@)��\,x�RG"���}sq�6�{y�(�֏����Oq��E��pg���1�o������_K�k��d}Ɯ�����(�ֳ~s��r)ͮYp�] ��[�r{)I�p��4�v�D��ٸ]!l�������g���莦�O
Ӂ��J`o�X8}��V�>Q��
���y��OF�R�U�#Hਏ�v�%B�&sﯗ��$U~�Ռ����멨�&��-�|>������bV_��>���8)��I?})au�ڭ�X�-8B�p��VJ���f���y��&Bu�U�K`"'���Gd�q�mڋ�}�j㰗c�eI�p�/m)C��eRn���/"�bVQϚ�`����]���*o���O}{IY$1_��WF��dxTB�i���1ZN���}�ʮ2<#Ϥ�(���6� ��n/?��]��?�l@!��!���I�Q�UT�, ��I���MtX+�_٪�H���n����3��7���2e�SѿP�n���x�S1^rSWvn�N�]� #m	��>쬺���O7����n�C��}�{��~b�-���W\�եG5�)��XB�\��?}ɴ�	Y�5%�0����n[����{�I��K�v���p�V���,e$�+Z����9�����͓W)1H��>>�+�-!v�Xs�N!��K��>���5�� L+ߐ�`A�v� �Ù)e�=7HR`�S��~xB�~�-n����x�v)F���.-~�����YU%�U������X蓦.�Y���>_o6��"ī�;?_>y�4}󘳥��*\:Ʌfq�h��-��TB�D��ϋK�hRq�Չ�vRߥP���:,�}�j[�4@�K��>��u�x��j(���ꪦi�|����V4-B�lK=�� ZK�b\�M�d`���~�������iv�N��Ğ>%c���i��|YQ��>*��F�R�B�� ���o;\7��!rڱYg���LZ�߻�s��[�&Yw��e���ak$�V��;�If%h�t���u���#�ͺ}�管y�y�=SNj����W�2����abb���;��Z��z܉���T�e�}�u\.?z��B�v%BL̿�v��)|����+�r��q���H��$n�˔�~�|����\R��	U&h�ZGݙT/����("��i�+~�ix8�|>�^Y��/��T`�^��;���jiŒ%DP�w�u�N%�p�'��<f80����k�x�H;%���u�_��~��O��⦪�ьە�Jfg��ԉԀ�Q�a�P�f �,���O�����Ԛ/�o�Y�Y0յx�ߦ;�Xh��n���5^o�<?�n��e�ܐ\�;���	�`��uZ���2�ܕ� ����Uٱ:��ޭ�L:'wtd�%2f냻�r����?>TB���)z{^��
�K�h���j�%����M*(Uܘ��غW����?i~k��Q�5YK"�U9NX�P+"���my{)�v�/$V�{�>#�ٙ�!g�cb�>�ϋK������,��}�dܸ��|V�\w-*,�-�
����O�>�s���E
��a�﹵-���,!|��z)��jj$�%�R��i,��+��o��~-p�A�(��d+�
E�������g��s9��x�z|%�i�/,j�� R+�[���{���O)�I�@�1�%U��W�每��#��R��j�Z�>�?w�ů\����`Z�/N��m�f0�njVy��tp:�z,��]��D�4�p�b����ڔڏ�_�K�,S���4v�k�f��-��1�-͘�+[���{��]!r_�N�*(� ����?s�W��#��/���@�"|�W�����ia�/m�Q��h�f�ZcK�?f˷	��!Z������D'56%b�}o��wE^+��<;6����"��4);��W
~�¢2+�P��{w��|!QWR�&%`B��}�ש�8�>����c��z���KO��qs��������턖�Gm�SSxy����V�8�l�,�P�9ӟub�8b;N,����ȱkq߻���.o&%,���ڢus�����=｝Y�8o[:F�BR*���X��i��T��1�ʳ�Y��_E2�(*�S4%1/�o��f&�p�X���~���tgQ��;K5�g\Ɖ_��pZ/�5�jkU��rU�d^���YbS�>��*7�5�y�K�}X����QU����6+>��;���s94�|o��a�I�B�~&qK�o��lYm[�G���:��O#%d��vVvW�K�3�|��
ɍ����"#Y��k�ع����?G
�Yc����ߏ�Q�`�	[Z��B�{�з�¢�����O�t����{���Ĭ���,�gO�X>l�_>�+-M�0�-pW�þ���D�R!HG�(/
>����ך���% �.�n�]W����\n;Xsr\m��q�g��nŌ;����o&΁[��G�uw����oe��BA�~,�Y`G��������Re\Бm�f��i�-��HG�5f	YDaYﳋ#��}�+�mno�	p��m�����s�\c�Z�
g"��C�u��ˋ�-!΢"Q[UTӾ��>mX����+!���;���]���/�O�����2+�E�ox�>T�J��>��<��V���v �+�j���J�e8���C"��wՌl��g���	'����'��G���\^�y�4���}�J5��MGe�K��TH���a�Ց�_ڭ.�7j�'����,Rڒo��W$֤�#~�k�����^!H�ü��v�T���`��J3/g�rms�;־%
�=C#S.H��zg)?��r�MT0�j�p����c�SgL�W����=��:���g��7�\���nEB�$_B�#���nq���x�(SM�.�%�~�����h�
�Ov�!U�,-�v���z�U�����9Ϋ��/�J>���W>=��%$VX*J��̓R�Ƕ��fW_+�I'C���k�ӤH���RwDQW����WW�Z�hˁ���
��j�TB����X�=���=/�ҳ��zB���Ŋ�i����_��j�@Y�hZ��߾���j���j���!$tg\o]e�]@Ύ�fe���f����͇��k���xI���C>P���:A���Nv��9eQ���x��Ɲٱ�YV�m���nnCx�t��3q�%;�mή�t�rI���p�J�V���j�.�z7g���{�a��ٲ���Ĵv^n����n@����3n1�uk�,�8���ﵶ��v>��G�dö���������S�=6ͳ�m�ϑ���h:l�
�9�����ݮ*�\ڏp�=t�n
\�+����ڻ���l%���p����7u�/��&Q�{j�<f8n��fsZ۔�5��cn4͛|�A�=�	YHJD������bG����k��p��7��	�"�項E�;1�~���*�}רo���������iP��;�$�/��u��\t��.���lO�����J�ct�-UQp�\2ڲ�݈;�J����K�ppR��V}���,�Dk�+�&+��h��4#��Uؖ��zӍ���8,7{ʠ,}����	p�Ɗ~$T}���1]�]Z���y[��~�yu�Z*7�������1Z����r�,�Z]h�����M��Y�+��V�\4��n�辜�P���=0�7��D��N-zF.sO��~��p�$)�o���؏����.�K���=�����tK��Țq��a�{��*!�.�e��./��9�
���z�ϝ�Y����H����g!g\tTQ�}90�Y.=9_��Z�R�PS蘔�N���L���?Z�I��qay���u����س!e���Y��X �>���v��c�c-5���]u�>n�Ӊ���>����p�Bb�#�$-��z_>���~��r~�+�+�B��z�����V����wmi�L�XIR*"�>���8.�,K���%4��W�{瑩��`�"Ez��a�8Cv�2v-�K֮�\�9�s�&��c9���u���F����*�e��QFK}�:�a+"�\Ɍ"�bx����W�X_v��-�y���QڟRY��ݥ��M#��3���$_LŖ.!_^���&��_\�k�]1�DW��50Y}���% ��Wm�\{�iӰK�O�����Y���S*o�{o�rA϶ԗ��A��R��S�EG]��9�m��Ts����t�#�x��:����c�����C-���m��=�)VuYb�ns��� _/:(��䪧}�m�,k�L�`~�qZW}��#E$.S�)���C��t���3�i���^��/�Mל+�W����G�	�[�R�R��0�$)��\��T`">���k��\k�Ɇ,1��*_f.~�>�Ԥn�����g�f�]��c� b�-��*C���ߚ�ť��[���{����u����?�D:ҿ��#��-u���VB�'�K������-��K�-�oU����]�$�ȑ�3J/+�U������ִ�rV���i_ܻV�]���,�.;����NL���ϖ���>.^��j~}8�:�\�E"t��ۥ�P����NG+���%Y�ڻ}k�,Ǉ������p�ӧ%ȴ����b����knՕ7����U��&���a���Ĉ�T�RO���kEM�I�D����$/��b��s޸��,�S+*�?K���:��������e��M��16�ıˊ�`K+��;d����;��]�%N�#�n� �B��.����MI\�sI<l�_-}5�rE�)��Wm�H�a0_}�#�z�)|aʟB��	w��ğ����7�{4}{d�&E����s�a����q"��4Q��1�>�
N]EH�j�%�`�L�!d��`��>�>����h����\���=ު,�UK�_	`���q_r��(XB�8����	��|�-����_.s�H��.o�j���@tV)9����gQ���<�.*����ɖ��L�9�����"�>�4%c��'�ag�}��/�H��"���߾άZ.�*��
m��_,��ݝ���j�5ω����'We
��Y�F���Y6s%�WŢ,���h�KhN���}P�%���o�Ws{��[���Z �{��$A�U��lW��6�u���!�+�����r���G�f�U�R�n ��:N�dQ���^������X6iF��A�5��^X�N�Wi��bK֝�3��#��!�Gh�u�wb��&@��6V�S[�577�o؋�SNX���9o��Dqvr��q��
�ހ�Δ�!�X���Y=�8η�Jc:p����m�ӧ�84�x{)έ���n��D��f.���n.�]�6�vD�^�Y����=LIlk/F�:��5ʹ�C�F���pշ;�2�v��
����8��]!cs7��,֔Ui����"0vn�}'@���1��s"�S���B]亴0l�-^�����M;�gG�X�q)wA^d�9b�3ȭ�ЪɄ^�E�5k��`ٸ�N�}>$��+n���Ta�*��"Mo����I�7l˥�Aju���6뤬L#�I]@��{��ْ�ՓGM�a�Z.��Az�!,<�hK�7Y�G��׉�P:�1��݌�+b!q���"Q<o��\�7���]9��b�-.W2b}74��q��e�	G)���e�JK�0�7�n
7��Y�i nv�uѽ�]l�7;q(N�z�%Yʉ<\�����sFmr\y$�tsiٮ0���RźI&.�m_���ob7A�v��w5��;_��V�E�{�=wC�1�13��b�/��U�/g�.S�*E�B��}6��8B�O'n#E�^�ch�q[��ȇ��B�X�I)��z>�X���f��s�k����,[բdx��Ҭz|z�c$ZJ���+K�mWe��B�*ZmФO�
��.�?��Z)������U��ȳg��^��A��w]�ݘ�\*�d���^!�����K�@ܱUa*�^o��ӧ�k0Q�]jG�Mx����rPv����p�����ߗ��}���H���Gݙ�F&�£�rw�7�|�/��Rw���R�򾯯�~�m��ӥ� �����L�D���7Nۭ��X�Z6��{J���.�6?�˵�)�����H!Wk-�X㬕�����w�s��8�g��ST��~��nX���A*�&hT����P��sK�k�v�,��q�4�Y&���0�U�B���yPM�������F<^���G1�z�I��/�<mOݫ��=+ߙ�$9�K�-G�g{�ߚ#�R!J��&k���W;�{,�dgQ*��؄΁ܳI�W!ol�T���I|�nex$���V=��i�K�Y����JD��R���,��x�56oJ��e��3,�y��vG�|�s��d5KQ�<�m[�5++~پ�/fJ���G˭N���	S������-���M���]�%;��ze*ݬ<��M��i��j��v�WLM���3�tU�����;�U������
�-7a��'��Y��v��v������[����Q�E��=����]��۽��(���{�c�5���+u������������=`rݸ�f��X�Y�A1c���6�6BA����Jq�	|s/�r�8���z���+��"��P��"�Î�s���4���{H+�x�k3���`���U������^�OT̛u�k�5��|�+׉2!��ͻ��:�;�P!w�7��Yx�������+� �gn�>��Wge{q�����T���Y!�4�K�qN��=�i�k=x�z���x��C4]�6_�UN��жt4���|ʹ�S��3�Ԯ�`��V�^��#��_.��f8es[�m�Vi��\��*=^�bi�b��OW3��𝻑\�'�.ў��㚣����G���:i�YHSo>���ZBc�z)Y���k���Y��mLe��=
�����e�/��Ϳ�O{��&�x.mB���\*g����e/I���h�Vf��5�<2ԡD��͒�*o��M	@�+;@�Y�;f�1M�ӫ��|jf��&Ԧ��*��O��t܃��,�KPK�w����{qa�')�Wnq�Sx;,v;I�3�ڸ{vvZ��!lƋ�lq^����`��n��w\���{�i��n�ڤ�n�S�n�r���t�/Bvɫ�0{��<�#Ջ=rݫv�[lL���63�ᳳ�}v�NZ��gû,1:yН���rń0�W/;�vT�=���j�:ƒ�=��[w �;j7S�u��Z!���k8�Ő�9�Ϯ_M��1��C���\q��I��0�-�ڏG0���m��$8�V��k����,J�-�U~~�7;g�^ؙ��v*�����z�1�k]#^B���@�m����.띚�x7�ө��2�q��{�/����G��S-M6ǆ41Gyy��|�c�*��6�����z�y`�j�v���-�V��V�=OTw!٦�mp�_M�`=�W�.���y�. �NˎeJ7�����b��g�NF��X?�%�ȸ,���i����#�%�rޖ��t^������W�����F+�s�w|�e��3D7�L>6�ȭX��:b�6�k7i*51ꛐg����X�I�jĸ�(���k��q��UVgyf_7ʃ�ʵ�3"�C����7��Q�M�c��������	��$V[�ny��]2k��:N���1� �s�.m<�u�u� LS!6'�$|%�u��h7���LOnB���[<�-�k�ks�Bb�-�w{En��5i��.�Q}����) �	�YͶ�i��񱗩�Jf��Qr(pĞQ���5�m������T�ҹ��!�$e�G|�y`<ߥ��M�8����C�T�� <�}d��c��9�r��^�e�W�@�t�9���t��ɝ=^%�Iְ�����fl����fO����(&�9%�O�ȝuؼI�����/j�7�ݒ=\�.Y�u.��WQ�S��G����a�b�/�T�a6�i�ҙ�l�}��(J�ښ�L�V�{vX�P�i{.��g��`�t'yJs����bj����V�i^CsƆ$��Fee��� 	t��l{����I�x6�B�"�w:lE^�)J��N�k)"|��-4�\�Hi����3�3����N*�?���`V�m(���Ms���ԛ�;0���l�g9PzǑ��'�v'J�)�U�s�CC3��D�����"���j4�t�i��~�W���c3��/W�H��Y�'��I�Q�E��`�׎�F�\����@�{��\l��=}�y�s%s��+	��ԖUj�-�7J,��5��^�W��h��`��2S]��޻�'5�~�P�4F7Ne���yn�=�{׮���8Q�\y�MAջڭ���&r���8CS�vUGDfg�-*����Պ�0�@�)֟{v�/-�M�]��F�B�/޽F��f�"#������&2ZB՘v�K���툾O�YŠm�pfo޷k�u~�]����c�y�؂xX�>u�W4_+b�y�߲�f��5�T���i:lQD�J���I@�rO>͘���S~��f�[�/,sҐ'~��������I�$p��3�L�EX�����yk-��`[Qb�RѢ���<!1�#�������gQ�=:�ֺ������x�:��=�7g��S0>o(��~\�]���`.N���z�jěR�p��nx�t�`�B&E`^�{w�)���`����n�L��n��}ʯ%ᶽYKG�z��-�;�t��y���V�v��;�
�����:'�i��W�4�m�dٗ�fiH�g��N�`��di��ʃ}�2��I�jEr�wٝOg�}��we�9rn�A��m�v��n��2�g��I
l��4Cb�)��˜�%�Y�J�фV�����I�CIF��l0E��x�䵐���î�*"�?m�x��F��'�m�6���gU���k�&&��ֱ{2�,�/]�C�v�7��2����3�ï%yf{�cĝ!@�a����:M���P�s����)�uً�r�8p	�?SL�[ճٗ]h�N�ѳ%�A�+7b���KɻUiL�zf"��=��;ֹ�ܗ
ʷ���e'%���:{dk�1���0���+�����!e]�~᭛x�5]���ON0W��:P��K�2��.{ކ?w��T4�,�Y�λ*:��|O V4��ڷ���ܲ/���E�H��aQ�jG��
l�jn���%,{��95�k:�%=i�������\|��@o4㫬PH���ƀ<���w|�9{:J(��6�[�Oo���Ξ���#�3f�<R�2ؗ'ŲHtS�g>��h�K��j;���Jo6j��������,���^n5H�N���6�[��^�:{��mو盿#I�i��N�J�p	�!�H*�vz�E��*���k���3�1׈8s�)}���&�'r�k.�I�8}h��cn�D{f�f]����x-W��1ԉ�C�@�) V�Y�dv�r�/(����$ˌ[9����Q㘲��đW;KQ]m^�E-�����ډϙ�z�ɲy5۬���
Խ��e���݋�q�����>�8;{E�YƵ̦�Z���ݹż\����W�8D�e6�;��٣ݥ�5ܖ��q9�^�'��:F�u����v�y.��k+���o.����-V�f
���
�z�7�h����]�m�ŭ��ka0��1�\Ol����	�<nkcl] �A��WF�Wk<�.+J'j�	�v/Fq�[r�7�B���I�i7�s����y�=[��cZ���a�����q1�!N�����4��)F�vw_���fWH��J�rZ�zF�`)��]i]I1s��)����1���O�����]��՛Ļ�]ui�RV�P�p�{��J�4��t1�$��
�����``y�W"����fV6K�ߟ�ܺɿ*1���7�9�W���3�q;�_;�~c��4Y%K�Ui�Սp���a
���<����"K1+e3�/�R�뵷Lgd9���_r�2��DG;�0�]��a����t �Qd�̢k�aV�:��] ��fr|k�3����a��Dk��R�\�E���f��3�׽�Ze�u)e�dj��wW<^�;�'EY���Z\O��3�1��:�c'f-�ٖ� W�$��Ε8m����.�cA����Xˮ֮��³m�����Mx�c(סXs�9���$�7A�@�[[��Tt'a(1d���qc1�{�+�q�Hm�ݾ�E6h�nj�ATe;�;N�b�N��Q쬨�.�]��4[-�jq�**56���}�S�q�;/��T~��i�ZY��i�5�y�ץ�?vd����㱖ryi&'ʜ�(���ay\�����'������fd��ߵ�Nk�F�i�&<ۆ���(w�kqAVM|��>.����"�uqi�}�=�ў��B��7�7u!����_�F/�ݖ؅����6̣��@[�E�2ߔ�~�nVz�t� 2�`6A��c6+�Y��s�ט���R�����)��q�ĽZ���<VTp>ASa_�~�m��J/��b�o9�����
q���Sp` �l�滌��s�a���F�`����0`��^�h6���/9���7\�o�r���T�J���W�)���j��{PVT%M�X����I��'8k�������kb���n�Z�t��J_��j�z�(x,f�ӯrNc��C'e=� �jo�rZ�g����V�
C�4@��}'��=���Z@$�#�C.�m�c�`�9�*^��y�T�(t��$A�MKb��x�3��*q�������"��u�Ya67(�Ӫ�a-�Kp+˃
W.�j�	��L*6�-�6���q9l�Z�9^K�����j�=�S��4�>.C����J�I�Y&�x�����g\�Ϯ�yd�e��/4�N`V}�<YS��G�~�1�g��N��y�m�5c��#Ʃ[�VH&�YMp��N�u���q;Uh�a��k�A��M��o5�1��ݙ)���o����}���m�Qwlku�33�������ZB��*8�7Y0���8����OL��֭�+n�vwFT.���a���7��%ͫ����㋕���˦ n��wy��x�:8;�zH��<W�)g`��}fcɮ=��ͧH�#�e{��Z���2��7����.���~ه�7d�r�� �sX/Ol��S����q�B#��F�j�ɝW��+ޫ�Wjx�#e�՘`�Z�}�K1q�=n�R��L����n������W����{]�x݉�3��ӻ=�q�P����T�)�.��N�v�{�jD'�s4m�)ՑBm�K���߫K`Oe&<��۳��)�"�YY#x��8p4S^�F�r�&*��f�t��9Rskt�.A��P�DK�j�S�SN�|���c�no�ˮ�/o��>�N�2.a���xN�K����b�L AA��]�e�׬b�^�N*ٴHj����aeWdZ�84(q��rm�7m����\Ӗ���pWo�����;֗�����xaV��YƸ��\�s�\c�s6�.:��-m��/)�p[����q��2�1���@g��	[��(�ł�s]u����Ӕ��O�\�����3`��ͺ\���V���Չ�d�գ���s �k��{ռ%��s���fJ(��E6�� '���N
P��4>���)���{U���=7Wd�F[-"���4�m��"�60Of�~6��=�x���ݱ5=t�w�ۧ �t�|��Q���/%�������TM] ��6­"Vq�m�� SJ��ᕾ�v6���X綣�z9	��:���Fq.��JVhbRJߙÈ�Jş�i�e�m�fmL)�o�������P�/S=�w�λ���v-��g!�2�����I���W����Ŭ�v�GI�(�+��7�O��p\�Po~���&�y��s8ۃ�.�(.e�;J�U暎�}�����ٸU��,�ʾ���:tw;X�*S�W9B�e�:��׎�v
'с����%�:Y��^ef]���Ǆ4{m�\��b��9:�/��J���#ȱ��+���`�$������&|�d�1�a�]Lm�9tJQ���@LK;�y�>ͼ���a��ݐLy�R��d�F�ly� �w�S����oo���v����J��ㅠxWA�[՜t�'s�/!N��72�1e�t��^�r���4�������Ty��H�]y��|��^뻚꾷:�BGq��}/���v6��!��!�NWO�9٨v���D�{'1�,�ڷC�,AN�����vN��Y��s�;�抲�P�sʼ���r�f�3����uwT���u�(7Iw$���32M�z9��u�j��R(���և3�ǯr�X��j�BXĭ��ՠ�4K��`���y+ r���Dc��|�|���C��P�/I56�����W�]q�c��o��r�]ER����uno	�y�z�G��M�����*_#L��:W/6T����@���b�CwG9�ܓ�K��V7Z�l�ᎎ�ѯ����۫�F>*������.�橛� �Dp$Kzl>L�c��f%FZn���K��;��S��0oU�폹����2��K���iA�	�Qv;��ks�j:���v��i7n29�@�*�s8�6�6�p���V���l�n���ּKn{nwu�pc]�[O��K��囃ݣ��秴�m���[p�s��D<j뮱�vs��l��d�3��-�W�i��NNOYmq�w���`�3ϣa��N�,Mq���1۵͵�]�3�s��}���Κ%�b�v1g��u��\W�I���5Fõ/v↖�/:�kpVw������5s��ush�Chx�ou�駶�n��mD����\�TIƴc�>�p&����]�E���Nv�kg��^�i�i�r�4'f��y�����۫r��]&�;��K��u׍�/G���zJ��66��V<m6�N���@�d���y�ۆ/8�l���-�FPz���y8�f����۳�nu[g����[F��&���q���t�%8M�:ػs�j�7#�G!�2�n�[�S�w'�8!����躥{'.c�n��naT�6���A\�0�#Ù6�ps���5�� ҃�1v�n���]L�g�7/
�ʍ��pl,<���〓�����#�ó��e��ݽ<��qm��n���DI�n��ۥql�'j���y��^�vv`�1<M�X�"՜�k�u��m�GS6��䶐;\X�d{m�۝�qn�s�z:�b��L�x���C�ϟU�l�8Eq��6؞�����Ŭn9�┝�Q��=a7�p�nY��tiĞ�b'q�x���	[�tX�a#�l�c��^�a��&��=<�]{<:�v91³��n��\�lۯm�<�N���vѮ,���k���\6�ו��]\v��O\N�&B�3N;��X1�q睱jK��\�ۮÍa���>�/n{&��n�\N���;�ї��ȘzvB�O�.��[��g�֙�9���\c�=fncחS�u�el>�^;@vwn�;���Tݧl�%λw@��&;`��;��۸��z��vˢ�g.�G��g��V`vwg����ؠ��sƱX�Vb���:1��>CV2;�x{a�烲���su�z�͑�.^��=��1>���^�e1��5l��5�`�ϓon7��2x�E����:� vI�y��,���(q%��,nzL�"Q�m=��ы6:�e�&I��+���x^-ۂ�睮�{�n�:��ō��f���=ng��]�- 4y�k���i�T3W[<Cʯ'[��C$Bݨ۷&�F;�"�z���2�`F%
%Z�ߟ�e���ʧ�s�����:'Ӈ9��1mΰ^���~��t��xl�L\4�W��ޒ�k[��+ҭ(�ʗB�����m�]��ލ\*�ƾڜ��UǪ�Z.�����Vm��{1���a[��Ӡ{��,�&䲛9�z�P�����hv�����f�ګtz�7�|�9��O:c�j�/c�kY�#xz�Xe����M2K�i$�E���y�</r��w'Vo]��s����oq���(�c* ��w���8k�^ul�)Y��-ݞ�E(��T�u�@k^KV�˹��#��k=Y�>ͫ�!5)2�s�ֵS��0��3Pˆ{y�0�q�P��x��A.��q� I/Z�,]�4���\�n�7[c;�A�n�������8������&��N��b�H�i��{�zS�9��9�����?W����n���ݝ� ����6g�C�����|������s���@r�i�H)�;N����2�����
�M���}��A=�E<g
2-�i�kwp9�ER6I�@�X;��O�ݜ{���tלl&��U�)g����'��]�#��	�j\�oeږ����6Ǻf��.�M��3M�
n���8��;6z�yk����iLp���:�o|{�-��k��u�އ��N��lb��[��4` ]"�2ۭɔ����6S�2zo��Ywh��Q�y���4��n95���':���C2�y�K�Վ���)8�bxR�DE%m^6�ݜ5Ay^V�<�e���| Лp���HjA��\�M���q�5�i�1!�V��eR�qh�=iJ苚ݳ.������C=�m�=�%��qO��0��֚)����Weg�o�a���ʽIL�=j��OV�RE&=�f��l*���Jà+ѷ^b*i
͵�Vk�b-�u���ez���N�ed��v��+ �zr^�qk���x%�2��c|6h��^����RMO*�|2�����0i�PM����*�������B�s�̘tw�m
Ͱ����
i�̍ʺ�����w�Pl�X�c�����ڞ�_]�V)p�*���-���ueU-3������©��W#jV�`/M�����Ph��cvo�ְ�]��1B��t��ꭖ�+2��V�����������ʝ\�k.�;�W7ϔV��7�o�<A��!��a���Wbg�q��wT�}b���yB���V�_XH�U������+�e]eǳ/9enp�:;f������ݻ��L��+/�g�`�0���pk"��cpS�~vB�Q����ۮ&R��ۭ�t�u�\{ku3����+Ȕ>����O=l��������ʑ�(?!�>j�:�6�^1Y�����ߢ͈�Ҝ�n˶���]�U�w��ʚ�!2O��ʈ��.Ѽ�*6�Z�FmXs~<���=}��o����h	�c��>����R��Xܥv�GW�2����l��W[�u��,R�x�i����6���j����~���Qo���^ ������������J)N�~�|T,Y4��h|�-���6���f�x��6�Q"��`#0���h}�Ź2׽�eo�NA��B�]�Zǋ��h��|N��u�euJ������U����ŭ�ZևT�kh��G�#��3��Q�*�;���X�$�L�[W7�ǥRh��S�_���0�ˤU�����ש���#���<��En�TK��,%Rd���g�inl.�V%�J��X�$��n{C�u�;=����<ڹs���2�8�g�b���RX��%Q��J�W��0��?�W"?�=�}�2kG�]�C���*�����x"����8��U�S{l�d�4��i��|��櫋Z�S:�T��yLxE�;*'3�-鼷�)b2�/_e"���K�NMY�	UY���f�4��(&�H�x��{������j@�t��l[AQ��4B�
�R�ű��-]vøH��R�\-;&� i��W���JJa�@�e�ILhݮD!� m�ĭ	k�<��`f:��sP[��W=�v �14K`��ί�V����;zB׻[��2ԷFǃ��L��A�H��n���N��;;�7M��9�_o�\_�%7�������ڗ�,����R{�ܴ�.��6�J�x -En^������6�߹r�-P�e�v���zގ1}Ʊ-Yj���7!� Z��)�Om�ܬ��:(�K���$M�-�I�������������1�Ɯ�������d�\�Z��;p��p\���v
TGh���;l��\�+�j��^�ql񼽓6�`FYI��x
⻎1�H��9�T���u�mF^wHaꦱmחd���vx�ӼV\�����{������M�;�7<� xv̜Ό
�ɬ�W/G2�Z�׃��޻6���s�Ꞟ5�h3�l����b����g�u˞�:c�xx��D.���5�&�K�+�wF����=�<jG������2]�:w9��eB�WA0cg��.���9��>�O����Gz���TTHTRV����k90�����Z�D\���9u�k�OR��#���^H�N�>]�#=�!5|�{�g�V|�_���e�M�D�-נ�DZ�xS��W.�z��exc��5/@z���-Wr���[~\�S)���m=v�Q�a��&�!
-���b��0�f
�<�v�4�}�{KW{�L{����=zs�@��5���Z>��O(�ބŭ�J�=����	AB���ڜ��f�m/�}6)�9�iQƗ5�w���Q5���2c
��˷�vϟ8;=�a�Vk��gS_z�9/���PVU.�8K��/@>�����ڝ��W6�V��Fs����Ҝ��+E"r��L�[��������Q���F89����/�Q��}�_M�����$������z�E��Z�t	�E6Ru�V�=y�7f��Q�������u{�6xqy��G����2)v��8�:g-j{��k�wce��$,��*�"�y�B����>�n.��+pdӘ"{Y�ɡJ�f |�6*� ;� �"�=�ݳL|��#A4�^R��⅕��&�V�O�뗠{B�� "��G�m4�$��2�����oP��Լ�F�M %25�8y�.��h�AE���?X�γ��h�GL����3T(ޯyF%h#uox��{��5�O�� �F׻J��M x[��^j�D�:e�Jcճv��nY�w�=�ڼ��##�%���8	��l&��.�~��Ӳ�f��J=�lu
��Q�hF���r-�]{zf�*�e��m�J3�5�t:�w]�\6�]�n�]��j�1t�7y�Z�t_�2���N}Fx[��¬���0����{��E(	E�z��A��y���Q{�L'd�O��!0�L7~4���S2��X"������OMR�����n���]E�z�����A
�h����ܵM����E�bi�K�E��$�g��Xȳ=�ܝJ�F<��a���Vh�r��:�[���憬 ��Iյ-�\�6�)٣���+�N�yk������o�hf�D��p`Ν���;M�(�a5�>�1Z�g�ݾ��퇦b��1�IP���E��n��;��;î����fzv�{�������v����/m�G�ׂ6�%[PEz�sW�����\ND����B*Z��֤U{���	�eF�ܘ�cs�}�=E�A�W:[�9�4؅
����� �Y��X�Y��-��4��n�ݛ��gmĤ�C��,n�����E�������ܻI��2�2�%��l<W19�
�]�9��x��A%���h1y�+;܅J�5V����USA�<�Ք\׮���"���H�M4��T�r�:�R���HZ<���W'�ѻ�3'��x� �n���b{3!5����y���Z�8|�J���F��~z��w�E�Z6nŠ}^~�o�Wޖ-�sk��7��1�:�\���,��,�Q�klӤ�
	�uu��gwf.�xilh�A;no�v��Fy���������u=B[o�5������z�6���s�m`�Q�k��V6]���I����Hᆯ㶰�����ɼ��̺9�7+.�K˜��VF���>�: ��N�!�,�`QE'{�t���e��7���G�h�]q'M����m�dP�Sp����v���3�ecVq*����Μ�F�x��[�۔<czJ}�aN�8��ڗnm=�����TN�h�Ҫ�8�pૉ�y���#�Z�����m
-L�{Ӱ�m�+N�&ϫ潷0��+p������+�	$��E���O�7�u��������'9:���{)v�e�����u<wJخn��V,����	2�e%�Ȳ�2������h5�Ս��o�2�fc�a�`��]�ʋ�-�V� ј1X'B
��v{or�e)H,4������!��I4�[����/�D>�t��3�v�랭'�]�����ch�ۚg�>�T��S�
���:��δ@�Ϯͪ�ˑ�im ]&�M6���]����^�>���Jט�`�=���i;���)
�*�t�1��VL[����Vb�~��.*^8#F��i]�3Q��=s�f]�k�˓2�Z���r�����S:-x�0�x�+��Lέ�G!�������:���- �ye�wW����]g�����s�$޷X[���ˇ[!��)�v����YW�h
��pv3!�{c�F=��uR���{sc��Wa�����0���ݪѨz����.z�۞�����r��y1ێ�j�;yC�U˱��&wv{%=J=�ͥp�{�72�ҁ����M5�w	�N�r�M���z͸�[��/l�v����ls�ۮn1{c�C��q��sqp���=���^g]���'F�Q����@���W�k{���B5V&ee7��L�h�x{�̉(�vX���8oIA`�!|f��f�����7`�B�
�ب0�	���pUR�mwfx��<���kS�iD1�܋����oFg�����~t�c����D�֪AP!�1�2�B{v��j������.��~�
t*xצ�a�]}Y��<3j�A,��4�C��2L�F����O���/]�VH橉na���]�lT��x���@{9�V��.���@���G�*EM�t�Li�`	=�z��zм��=3ϵ�i�}6`?wlO7i������B��m˘��kB�g��ڭ�7���j9��vdE�� QK]�S]���s��ht<v9#;�I��Պ�\��1a��ȝ����������!<��<BKKs��۫=.�?:�ؘ��_�y,W�4��܄|yX�6Oǃ��R �CtiҼ!,;2����ս[��$���x����������QOADt�tp���vK���ܪ[u�{ksLBi�f�V�X��,T���XǦ�ڕcXF�R��ߦM�S�nf��w�߫i5k���x6�$츶5x��<��gT�NJ(U��O-�i���Œ�>�DLK��� ��R�n�/���/�c!���i��;�ݎ~��sfjd�>��!�R����-��Պۏ3Ч���������\�[�fe��Lq�0^7�p���9:����V����h�‡��	6� �u�0�m�'�{��([�V{Ԗ�]=N�\��y� �H.���
�{X�a�{F4=rr�������[�����9�;�0�.W.k�O�/�-�'n�:�`��5���<zz]ɪ�h+�*� ��<��z�ة❐��;7r�b34�y�uk���7ٯp%�N���A�f;k;�+BFK�v�-&�K�a�����:����x���߇ŭh\]��?7��������{�Co5 �^WZ�Mѓ���g��V1��b(�;-������(s����D�U}����L��L�(�u-h4�MCJ;:�&�P���rt۫�s�vwi/�ג�Dp�2���4�|�P�(Գ[l�rd=����[43�N�/?W{��$�U��C`�]CL�%g�*`L����-���������6��M[��oyT���$v��*DC՜�u',� :s{��p�s�Hx�.W{��+�ֶ�X�qPv����d�&��<��q���}6_ѧ��=+5CUvMX-����'.�q����k� ["��J���X����(*�5t��[�Vk�yȳq����07t!r���Ǉ>̀l[�Y�����vN�Dv���u�ZI����srq�l��㮡k`�2�r�D�����!�}c.o*w[�=V�w��P�L:sb6hwq�k�!|���t,Bs9(�`��0ۈ���7A+FP��\W����;mEw�+ү���o<��8u,����4䩙���H���y����Z�N�	8��W!齹�)Qv��7sc޻�x��
��ׄ���99���2���<oG\�a����!���[�;5u��,�v(j+�Ւ4��bD�]t����fqU����ڸ�����7�]�*j�6�d�;|P�݁�j�gy�y�ػP���P��&�84.V궳���V;��]rٳIʏh�A'z1
�c�p���Z*��7י�f՘QQJ��T^�;`�4UK�J���ٳ�z�\y�:�G9m������W�,wr�`nV�J�i�K��+�0��H�{'�û�铥�d��8q34;l�buB՞:*S�Uz�x���r�O6�ܗվ��a��3�uS ��t ��}7�ORUo�;�w҈�|�&h�R :M�I6}[����r�pj¬��~�wG=�e�3��z����t2��c�� ���/�s���BuY�x4�pn����ut�f��Ou���ݵ+�]z]+�F��G��Κ���l�����LZ#�Z���7X��y�-������m�t�j������w�N��м��j��J޵U�ݚY��=Y6��.�sW����6�b�ϱcaV�����r����)��eJz��O��,K{�����@+ �n�mm]:���@�'�H|��B��>�F��Su���Hޜ��R.�p|��~�����t;M��`�D�W�)��^x�>"J��G�{;�v��lɋ	zzzJ���ZS�z{�G�%3��1����/e������x���ˤ�C[�D�R�S�(��@P�	���Ė���1c�nc�m�5.�n�����`@.�fR)����DQi����y��#^��@D�p����[nN4O{o���@jPW����,�J+�M|��H��Nu��aut��a�"(J��s�N�)��W#�N�F�ι�oh���o.�zlh��|Y-��l�t���9�d��,�Aߤ�.z`U�(U�$.�i7����4�nz��H�����s�H�J_�MYKV���}�~������-�j��z�Y2D_����2��.2o΃>~Uـ�rm����
:�˾+\8��R���F�$�3K�[P]���A,"H.*�2Y��\�5h�	�Z�3��}�!���-u���h^X�h\������hRLS��5�'Y�l��mΞ]�Ϻ��v���l������s�N���P.`��X��R
7��Y�SՖ�yhoW��Y"Y���������ˢ�]dT/R�AS��Tե)�ƆR&s�_3zQ$OaV*g�=��r���ۼEŧ4��F�)�h9��FQ�)��0ي:��C�X��fۭ$S�<#]�yP;��q%Ȋmr*�3�E*s��ݎ>�r�嶫l�V�R$J��lM��y�6�9�#ٲ\�v�OnG1��!���Ŗ�rv�)M6�t��^��r���[O����xM�[�d������t��>��T��rjc��$K�\���+��Z��mZ���ƺ�c�W9K��d�lu��������8yœU����[lx�\v�6l��Dw�H`�g�;[l9�����s�\�v)b��뵳�8��䧴�hQ����)�y�ֺWth�2!EU�n��S�-��k�I��شFiҢP�~��y���ROC&��]%�@rռ��t3����zХ���
`
M�I�b����y��z�Ew/��h3Eoh�ow�c����VG���{��pj;��ѣ�����)	s}�����J2I[n&��� I;LzM`U�Hĕw�Ù�<�(=.�L�_��w�O+��z-a�[�6���wHȩS��$�L��M�7^Y	�E�zh�^Y��^��Rv�����(�d:.�>�0���h� �[��'�>K9{�ˬߣ��m�V�I+>���"�� 	�X�8�k%Xzg�E��ל_�s`X���x�5 �P��s�oV�4et�c6��J$n&QƧ��4���5�����m���:�댜]�Gt;��U�p9�]h�.��s�j��w�[��`��b�5� �r�Z<��v�#�e�O��>�F,yG����z�PЫ�ҹh�AST"�M�sA���fC��e�>j�r�M�{~@�p.��c:����q��wIwT#�RWK�b���W�9�1C�.���J��p�sB�8w��ť�];rn��5�m��=�0x{�Z�̒J���I�eV�n����<˲�d�yѡW�_J�Z�-�ͷw|%�=u��LS�N<�Y#�e`�|����q9����򳵊�Z�)��#��/��"�,�ї[VQc���:�ٯ�y|vox�0Z�k��Z�s�%&��s3ڧ��c�g=�ۧe�3:��\��@-u����A2��h&�܆�^������	Br���]��zk�$�k�L��[��t]�7���z��zl�7�C��cn��j5q�j�ױ�qv�,��fw�m#��:�5��x�9�t7k&�֛m��gnKZ�6ԑ�*�9�*<�3�e���W̒]^u�K^�i��U0<�tg�y�lc���S^��=3��A��^���ѡ����Иǝs�m����O��˫�>-e��{���Hd�@�R�3H����{��n��8ʽz��к�3�*��ح�������[�|���F0�CB�Z�p��t�[Hm�CVl���'���c�W��I������փ�B`#�1&��߹W,��c+榟T��*>*��I�{��g�Wǎ1���՞��vN3^=\�k�qܫٺ��+�WJ�!0�<e�t�!6�Z��YLM:D"�Y����{}+���ı��dd%�C��fP��<\V<v���sǷ���ս�1k�ɾeζ�x|{!*B�Pe!(���u������X�����9���v�3;oc��H��Ue�4�b)u�M���U�{�f�ۢ�5mt��:=5�ћ� ʔT~��<pm�xߟ��J��h�F�BȫWe![��1'S�*��{6a��R��\%�]�����Ё��c%�i�B0f�A��^�e�f[u���O:���DL	I�X��A&7u��b�ȭY��5öfo�������~��t*��B�n��Y�_WVk�{}{�+8!�"�N��N�M���Ou���ʭ3<<[Xn�JU�%s3��X�H4uR�\������l�}����ܺ3A�gj��PY�%n�6����Y0<����j������x�H[j������et��"���{p�۳%{^�m�!>.�$�m4e2���o`zyҤ��ohy��aݵ��%h��5�L{��
�����b�[���@9fm=��ur��t3]N^��ح�i�m�䜖�\�V҆�ԉ��W��u�]��$�7?y�E���O޷�8���s�hT�|%�G��t�؇0{<(���N�o��z}c.�k��8q�o�T�rRsS|~VŇ�d��	%ůcmn�w!w�$���r ��n����z߮���OMn'�8b9��٪�t�(�QQ#�C�ZkޢIW�n�J��]ٗz���S�9���\�n&BJ�$:�;xe�#9���V(�~�^I!yD�J�l���k����Vw�&�*���o���s-�ؘ�U��ߙ4jk/:t�6i�r:J��ʮ��{}.n�R����1�)"��2�e1���h[>=5�O�j;o��WH?l���/�[�O��Ѿ��6�_[!�9Q_��1u��9�Ѵ������d�ÂW!�o���[��*�xӕ�h�Y-���um	������x���u����돐}u�lU��)#B�&s�(�w�dَ��S`9�1����bS���շ
��e���[4z;z�j�A��:�W]�|�ۭN��Y6���^8��Vݍ["�4\]Wkq�"\v�ܕ(��l�糱Pn^�ql�f���ɹ�㵱Pn�9Nwmon�A�NwδڈGq�\/�;�:�Hcv��]��]�۠��G�ں�u��ۿ�W���rgdx�ڞ�8����=c�:�Nٜ�r��mk�������&��.��y�9gI�V����%V�*�i�{����e��J��w�v�[�˙���qǄf]D��-n�Y�s�#�ſ��g)�	�t)���%�32�4N�ٝ���:�����LRXlu{5��D�N�4mmo��>���B����1!
*�:I7]�9˵u��YC��f�r��<��v}W~9Z������%s/M�NU�*�:��Ω���D��J)��%�WNVA�����Nԫ	��i��<��)g��9���N{wW����n�f��b̃�U8]��j�%��Vsmxrj�j8�N-V���ʛ��\"6-M��}�;��Dp+�p�B�	�ԓ��]xxVM�7��4�d�n�M��nݼ�y��Ү]���m��vxhō��8k �!F�%N�Y�O{1g�|�����{�*�LsN�T:TJ K��wX�R�S��*�Ko]�{u��zyr�A�f�#%܅��;Z�*伫�U�KMfkM�:oeke��ts2��pӱ��hݨ�c���6�Ϭ>#>X-'MVX�ѝ���Ů"�)��3�#�j��[��ƀ�c3}�9O^�os��쬘s|���=bʛ�q��5����s�4
M��
M0�u�hy��=��VS�T��33y[���F<c�a��{���]dۃxVי�μ��'B��a�4��9�q�ý�x:]������]0�*��Nx�J.x��B�	�{�6���Y(�M���,�;����&@%�j�j}�0�y4q�2���퐊�zww�o��&���2�{���V�ܫ����jg;<]�S��G��g�ڮ8�Md,�����'�c�0{=\h]ŭ���۶� X�]aQy�v�g�.�/z@��-ٯ�7�q��o�L�U}3�R�����i|�M��:5�K��!��K���%y�j���z��F��l��y�<�-g.�-�m�A�,��oz�����~�3���/{�u/:	��[S5S�>8qL S�Z��������=��5���3.�<^:�&��.ɗ�V�|�]!��^�Y&
���M����ދ#8��`<�ׯ�ov��e)���t�(/�j+4'�U��J9��6��⃫�?)��'�"Lyl/��/W��.4GEG�s�!ʒn��m��;]P�^��u3(vCJ��W�n1��{`��^��W�ײxJqeZ�ٴMP���o�h�I�~����Xf�RF ��J�d$�ަ�Н&��FeҸ��O��L�ݭݖ8�>YE�������|�-^Vr�خ�˻�fj�Oi_Gȹ@#�U�U+�5��`�:���D�����5�=�8��i�R4S(�^�ޑ:����b�coN�`W�ظe�%-���J�iC�mz
�b����(������˩�C+�f߽t�Ŧ�@�k$v׉��*�ן�,�Zz�e*A
���`�R�����w�,`~�*�Q����S�dS�&4�'��m�,��!�}H}KTvR�~W�uve.7��f�2��=���Jd:&��s��@�iQ۲��1y"[�]Ae�]
	���W�:ݍ߽���:,��{ë��V����(��G*$ͨ��[���Q��E�=���oXF�ν�Ah��Ø��Eӣ�cʸ�uC�ݫ闏�H늑�	�Z�W�S��ᖻ��:��)u�y/���0��a�ɒ/_=�x �p�Z�kۨ��nV
֠J�9e�|�<�C�Zo�'��S`��wv]�8͋>�(��w�ԑ?�6��1�(��|��Djrv7X笠���)�����Y4��YN�Bq��V��*��
@vW7���G�Lǧ+}�ǙK���3~UH}����L�܃&/_;ev��J�F���}�VS�hKy���n��Z�ͽ�^��z�׎�,\]��`w���m[ݍ����!`����m��*y���\z�`����#c�$��i�Ii����5����ۧF�+x�s�:��A�v�]	��u躊l2�n��f�K�S�칪.�	��K<�@(2N���e����ﺵټ�3J�Ӽ��z�8�Þ���C�˻��/϶�*�Mڭ!j�ew���~\.������Q�q߇-��o��s۽��\:�s*���f�Ʊk̄�^�6]>ŕ��+|-��t���G����\��}�7�-͹6�rd��gv�{��x$ޙ�f	�E�N�:���f�S���s��d�Ө�����vS�^.;��9u�c�A+yk'j^݂��#�M�D���K���v���duyJ�ܼ ��3�R,�N�	VR�ͷI��t��10������3&p6��RmS[5]r\��]lJ��h���P�(�����ۗ�5t�䎳��.!���%���x{S�3����<{��G@��u(���8���ֆ���-qe�A{\zR�oi �Ӄ�Q��#���ʒ���3�/]Բ@ވ��CS~��G٫^�L������N��s��n4��y̥�nY֫3ay3�rb�[����e�Ȇ'y��C�U�H�͙.�٭{rv�����S��+M�3����*R��A^�Ψ�;,�A�[2�W!&
�\v��9�2��J��V��m�x;�l6�CV���N��{EUq�n_W9R�uX��qk!Ԁ�pf��<�6+|N^���ޮ��*N.��2��е���9\!
�2q�ۨy^�:��.]d�B��7QG3�R���콣Ϧ�B3���]���΄@�p��w��bn�� �u�>vwn��HQ��>�Q�9-�����pe�����Ιj.�a�x2�DA�f�'[W�x3}+e�"ֶ#����w�b�en>:�t�ܺJl黮U���S{��@ǽ��i���Fu�.:�s�Vx;v�"�4��*��S�B�mܦ١�4��w5�3m��-�\8��&5�;��"���֒IJ�N�N��S�s�B��k�ڧjje�X�7]��uo(�gƉ|q	Gj+�g7z�<�[\'��vS0�vb����:�B۵��'�&�Y�X�r�[����	Ok�ݰe��vv����C^Ljq��6m�ޙl�:��]�$��9�՛���;�����7�F�p�cv��fJ������%˱�(�V�q�MRb����d9�2v���<���R�1���5\C$���/�T�:^uԣ�S� �R��gm�lp9}9����ш��-�� @p��w��l�{\{�E���议MϨ�!��W��۝��Q�S�����)��|�wf62v'Q]�As`zwa�K�`Bl
�1�vV4ۆ�x�ޱ�rv����@�<㣀�;7<v��/c��j��9|�}��׮/m׳=�%�Gh�=�9���9Aw#�;�k=�l�pg`�8m�<"C����=V�y�&��Ƴ�v�-\hl�L�=�G<�g�E�:�nM=����1�[���Aة��%ɫ�nحקĖ�n����[��z�W�.:�wfi���<w=��&ޮ7gz8ՠ:x�M���������X|{Z���'=Gs������y::��;�����Eomno\v�__�u�A3�<m��}�e�jͺpWd��{Qv��uڠ�
�
��v;t's֠��s��wW�쩚�d�l�!O9M����p'�Ej}�`�)�y6#�m�X��������R7�6z�$zW]umUත�ȩp��`'%�[=���Z 쎺�l]�.x��oA�ݭ��p<u/e���[���︶)��L�Nđ�����mݬ�7]�۫'P\�nt\&����v�[�u�n��d�lu6^;�N��ͮ�k��ޮgZ�����]meŐ�X4�1�tc�۞קq�ŝ�n��
��&�ۇ��m�OS˜է�����
����`�oF����3tvu�ڶs֚d1j"���uփ��槥��c��۟gm��/p�d�{m�]X|*���{&2��� vd�2�b�[��䴙pk�zka��X���ܽa�f��7��knN����հ�s�_Ln�.61�nT�[<��mm�=�.��bo5dI��t��G�U�s�K&R�<���"Q�ζ;�B�=Ӷܗ�S�WU�^�����:ݦ�;n���oWmF�1�]{���>�Ҹ��ݠ��J���d�g\hWZ2c�<m��v]d8n�y�����ڟ}�>������x�)�%���y��m����v-��L��x�#O趚����X"n��n�[D,�Z�=W��vG��e7F�f�4����0�M���I�y(��aR�j��ERe&5�w��X�*i��<-� ��&���V��<���>�0���}U[�)N~�8oT�
����~����0[n�����4	����u{KR)G��Z�b������OG���*�
��fT�6t�}L��M�	-� &�S^/�u`�����U�J����x����^-��z�w�>�+���[ƽ�+Fm"��1)"�WtBH�Y�<�C��vC�=�J:ǔ�~64��A�3f���TJ�W.�^.ݪ����$�v�ߨ�/W^�r���{@�vѪ�-���۟+�,l��LSӂ=Y�4�c��WRsunŅ�4��[M��cOZ~��|��S|B��:�~�(ny_so(Q�3�L]/�xγt�+mn�'�	k��{③�a6�ŧS�H�s�)[��K�0�\��{p8�X�9V���%��F`��W}X�B:Oj��[��
��|w*"���2�)���]�SR]fޣh� �'s���Uf�5d�ZP�{�ۘ�9؃��v��c�^�ޚ����A��y������P�	��t�Ae��u�o�=ae��U���k���=���#ڒ)$�V?`�:yX)���,�Z�N
�>�߽��Q1�S��chmj��I��s��M��B�;�b�Wg_��7J~o��bk��-:��+�K-���om��*��D	�AZB�����My�W�p��6��Hܘ����[��q���OokW+����U�+��g��������;�y��l�{�p���GU��-�s�%v�cH�㇓��5�k�Zx��ۧ�N����@'X�E�)1�A枷+�Y�Z��VyS}�I�_�[=(�4>�G�J�Z�6�9�6�x,EW��V$H�M2Yl�
g+|��O��||���tD��?��7#\���f�z��-�w�n�9�y�^��]�U�=�sX[O��e 	tA��Z`��?K�R��nT)T%�ѣ_��$��w�7�[5�^u}�HW-�B��E�ϯ���g��z��L�]�F-��FVp=J�R��ٷ�ҝf���(��PT}G�_�*��!�P�^)1�E����(�H��L��aӱt7�\
�z]̩$���G���2eg1�^�;	��{����.�x�+��%�Y�����5lL�(�&����@�ok���#�ҳ7*7I�	����sڟD��q[��U���W]g�2���;a�&ʚsg~���g�K^��IѢ�tS�җc�ac�,m[��\��몛v9�rv��y0�5V�(B'U$��C��y;�[�lש��q�X<�yP�n�/��M|U񔛖ar����^���c��Q'H6
D������[�bj��e薛�Sz�eN�	rQ��k��Y�ԞFHT�	R�z`�{��>�m�������4��8��G��Lc@���o�Y`]̃�G�[�����m]d�.� X�㧰���JDh��A.a2e�Q�n,���W��?��ҧJ�S>��þ�!�dR�[w�y�T��m���1<�� ��x_eyfX��i��\��YʸT�.�p:��4tG�)gMݣ7Z���}�{@�L2+t�E�Ң�n[\�Y�2M�j�j���|w��,�2y�~h���-ӱ��؈�77Nmm�l}ɍ{Ҽ���gl�3O�,,�{���
1�5�{ރ%ޚ��A�^�G��/3���1S��N�AQgl��S�'�Y���c��{1��`Ղ��ں���vy��e��l��T�|9�/D��u��<ó�W�:�V*r�=Uzyɼ�_vD���uw_c�6���b��1��J(;K^i�o"���I}�O�����mOlux��l�2\#ww�K�w�W-���|���Ux.ml��V����?3��r_�%bW���_#Iz���*L���kv��[~��@�h������o2�7��'���{��oA�o���T�#�¥h�A:8�qBU�p�ٷ�[��W���.C%�n�,��đ�|���UO!Ah�7�:+O��Rӫ-���hW�����g,�"۪U\����l��=gݹaP�`��"�Zw�)4]��5VÝ�Q��1H|}j{=6��'��t����}��i`����O>����/�e��UB֚�AQS�]���+�x�KBE��3�7HnK5g�o3�K�N���m���r�ӛ�m�$��m�k��GC��ps�0�iy�mAmk�|�c����G��QYb7=�s���r�P����z݇�ȱǳ܊۶gO�h��n�N�H� Z�$J<{<Q��y�v�u������<Z��SgM��.5��S��|�[@�M��^���@sq�ڡ�މŻk�tn���5��nOdj��y�;]\;V��-���c�e��ptwRSVM�^�>��Bv�ܽƶ:㮧t����Q�z.�cLn�^l��ߣ�ZM(~��&��pX���Ȱ��Q�T��ǹH��Z��jQT���V/��A�C�SL^F��|�W[u����n^*�??�2�Cm^����y�wk�zCU����s�x��T`���}�%�y�%� �$&�d��0?6�[k��eb�4OW_�Sp��3�c�E�U�w��9-�!�.y�N,4��g�!�&D�$XA [����:R�u7J7�q�պ�!�*A���@{�T�r�^f[n�s�X	2����s9C6dJI��ӈ�)"�.��k��7k�b�"��Ftm�V�ف1��ފ��E�{c���xT��]�v
5si�{�
Ѥ#cY�>�����P�$�'���}��Z���d����2�A�ӱ�Fh9��]��;]9.��#����ָ3�ܮ�cr��	E�M��WU2�%tF9���qAI�o�����P�]��I�Yu�n<HSc'� ���s=���:�4X@�
(6R����O'������&��Ԑ����6�HLA��m����ٕ�q�zɼ�R� x���{\����9c�Sy�j54�u���
�2녯w,��s�PjV)0	�ѡp[���
�b���<}��O�!��N��^CK��3���龼Hco��`���.���J�6�hS���y^��>^��w�&�ز �HTm�ܗ멻Sa�++T�����������}���9󌏡j�3<����yX�0ٮ�<h*U��b�<�x���"A`�y:��:�҇We�Pa
����>��Uv��	fAlh� �L��3���+�S�h�^���5�����#OU�6)ۭ����}c�F��V�d2U�f��rm��;{��o8���)���~^��Y��=/�')����.�٬V|R��w7!���d��T���s�u�� �n��ɠ�J��C^��cvv4v�$+@����EQS��,�s��V�!�V�\�'���_��СJ�+���]ϐ}����w�p?��L\����_Nm��Ә��+����ց󡬀פ���7ԧ�ꈬ��tM&���0�߯��ճb~Z �f������ǢJ�w�z����`�}�Q����	2E��;C0�g����ꒀԈV�Wvg{Ct6C�v�������6�Y�_{�y�<�T�̖�%����q��E�'���WSS/j%��jIù�R�3v��׾����,#Ҕ5�>�46{j���9��x)
[����>�T���{����|�F���i�v�j���~&]\�d���a� ���=>��/�
<�^�:��=Mм��ovm�	�z����{b��\!HT)��E��!,��k�����-O���[�t�X̰��ׯ��K۵六�1F�_6nv@oU��
�wM�>����P�M�>5��[^�,b��Z��� QW�l!q�u��c[�ɦ�ۂ���Nmv����7l��v�:sa�sQ���q��Vr������n����Xƿ9V�ϴ�;:�c�v]��1���-���eV(��^�0��|*�(�7�I�!",���i����j'�jX"d��͠Ɔ��o�f������<�ɵt��!v��c�u�2����{[�2:OыǏ	�������,X�E������uF��+[$�Ӌo�v D|����l�PkH���uT�����)���68���'�Y8�)\���~Hƣ窍�Y�'Uj�jQb����[3o��6`��X��y����m���#����c�9o�h(����ʙrC�z�m�q�3��@{mƶ��ڡ]��$6�t�����M��ƥ^�S%<�:�(끘v:�����43��C�q��P*��ߩV��6���RPA�̋3��V�DWU�t��2[)�ԟ�oġS2��*��+�R��s.�+���Vj��תy��;`��&��>�ES]/P���=}M+���o\o4��N֭q�mlP��QM��l�רϵ��@�m�E&-׭��l.;=A+Tm���A���:�?(��Y��k/*	g�)�E�Z�c��O�loRCT�~�����E�ɬ����wy%//7�7�(����-���ȇ
#�Z��X*{4{d]�~{���A��r�wB�Y@�T��!E�b�L��y�2A�����i}��ޤj�j�4�L��D��ni�$��Vb�=��]~�^���O��,����Xͱ�ݼ�T��;�sb>j2=pa"L0���T�m�cEN�O@����Amb����ͤJtǙ�f�o8���Bm�m�'Aͬ��z��"������	7�
����2�
C#e+�&ʭՙ`��W�Nvz�X��ا�s�ݴ0'u�>�tGa�º.\��#�T�6�X�I,mi"��s��	���'I<Gy�bզ�)��q�Z���8�flSY�����N-Wv�E��PRd�yl��%k*��a0�F�0��d�7d��Ğ"ՊHn�ڱ�8���wn{K�x"��{��{z��1#[n�sǞ;T���n���Wo�]ȥ��|��	�b���u�c%ۃ%��;x��}��=�%��og����u���n�:������05�Y^�m-�\�j6�;'6=p����I���ypk���֓�rp��X��q���r�:�K��7�㛙�N�^����n�
�m�9�Q�����72�g�ӹF;/oj9:y��\5q��AE�8�T�����:���v��������K��?�m;���Rf�<����> �~9کWOty����ۡ�ʓ������(y�A9N����s�t�]�O`�=9�m�|���ͳtp4і�'���9��/*7��d_Lݭ�%���*W�.x�#�w�@��D&-��x�A��J�M~:v��k�U��']�z+l���~#�����X�5�����Ib	Ir����J�Ƥ����� J�	Q�D'A����[���@�OVy�*�Vw�^��H�W}�g޳��
���������l/L�j��3ы�ׅxL4�}}���MB�- �mR):�r?t~��
l�~B�$�$2��$��&e�������F�j!�oz��X�N`�B���/+kEQ@�k>\��{��o{krY-,#}#�Nɷ����gl��=I�S�;o��>�8���u��QѷP��Tն����f,O&e�r�A����J�7�*]���f��w)�ue�$ĶZ�ns^ �ki���u�~u�P��U����{S8j�F��Xy�`�`�9m:��A�ssyn*�L��M��jѺ���a�S�x�b8��m�l�7u��+z�0m�5�[ye*���N+nX�Zͻ�w���f�>���t��ʺ��D>,U>ht�	�)����0w��ۺ����6a��s~�8���)9�dTN�+�涭�ڪ���G`߽5u�5
�	;��Sӕ�1��1>�Y���@���[��Ȝ��"���Ne�TUY�m<U^�w:H׳�ޗT-�V��U���M�l<Ӛ�'=r�O�Q=o�sz���
`���iVid�Z��7���v���sE�#�
n�g7��پ\#���K�c����%���\��J�H �u�h�0�ʿ�/άA��EAk��7k��w9�fP
��H�s��m�}��z�����6��`"1iLUa�ｵ$��S�4B'kCt�Y��{5��\�i��s�-Ȗgn�{�k��X�:��i�̯_*�qX�6+�&��!_@��5�&�ׇ�5wO����gw��ܸXS�qGDP)J��7XO�M�0WƦm��a���>�[^|h�p�M��������2s���>>�Y���6�bZ�?\�
���{����nʃۊ�v�:���,ӏmR�s~�dulqm�9T�Z��d�U���o��C�ު2|�5]���;��d�����:lS�ELASS�
�ݨw�]�=�ʁ�_C�9չ��s�
L�ge�Y Y�\�ރ�wL��u��̎]ö��{����n"ha�ۘ���f�'�|�u�>�R�kml�)�u`y5�^��Ô�e�-0B�bpt��9�Yq.����L��q1jA�d�x�FG��f���:]9���O<P�V�g����+)�)]:�O�t��vi6��h�x�$2�m(���8�E�>y��#]M���ڦ�(�!j�ӆ����]�Q�ê�#�H˔�TZڥ���Y�\���3�<��;�bWoA�Y���ϝ�&k�v�v^���n#%)�w#F�u���Lf��쮼�-�֪���n�z�b�p�Xsy]�1Z�I{2�
W�I���2�XJ��[�Ձ�t��0�L�7`[8+Dzd1� oZ[wR`�o	����;��]S�=ɚMv�૭�A��ͷu�R��}+#`��2Y�:��ow*��b�8�W��K;*)�+����»G.�O�s�;��p�VO3xt����,����,����9PV�'C�
�i��՗8�P�7�J�^�>�t¡�:�}jH�
̧��m'��*`��w����[�s:��77U�OP�*,g�Ưfgv��OR2�Wܮ��wF��6��i��׽Z'��¥[��s|E覶��ou �^c��̘���;
䓻��z4VK#�w�6�ڒY�ɰ�'I�f��f`�]A·����n=#���.fA}.�pv�j�����Į���ݲ��/����4���G��=YEI#e��2�f�G�?���V*����U)8]�_H௞檾��VEkA4}����
�!D�W�ZsO]�^�K��}=Y��艩�m���b�Ͻ���* <y�`��غ�
��V9P��T���,�wJ\���830}��&�zj4��T��w�9��)e���uKb0KmȨ�ŊXA���]����Z+�"�bD�����U/��y�oV���q����۞1f�$޲ڐF5NU�5��W�q<�Z���/7�Fn�U�Q��MYJ�����;u:�[F��X%��繞;��rn��{���ORU6MR��E�숸�Z�y�[���U��R�K��Nx��Z�J�R��ݺã8/:�-F*�⤍�f�\t����7ۉ�@(�j$f[V>���D"U���Ti��n��p�ʘR �8m���g�f�vg)�x{��%�9D�/5�;��QX���ҥ�'� ��G�U*`j�*�W�#����И�� ���7���vil������a˦)�5UFt�8�\abV.��]��/W/KXiE
���ɮ������5r�����^�WR��TJ�ڮ�["H]�:A��vc����X��f�����t�*j���b|��[}2lz�P�����.e���׮�W{5�X�I�V�n�J��g�?)����6Ғ�N�U�:_�B���n�*��h�H�t<k@}���I�Z�k���Su��szjk�x!��m�̗s���`����h^�-m��&��#�/���f5��(�!TZ�x�jqLT��K*Ė���´������g=�+���*
)۪{��\��Lvb�Q�U�z��w�#Iֺ+����s<\+���J�C!Q)#M�z��vxB��K�T�xk�ܼE�/�@�B�V`�
�<�Cl�;�pÎ�w��ֶ��݀�������a]�7_Э;BU�p�ic��:#Y�=r�q�a�Z�^���t��(�.�{�j�c�k�%DI
���ⴽ�f[��<t��xK��P�z��ԉV4������(�*�=N�UAR�II��j�4J�	��θ��"����!h�^�{���W�%"T�����VF�SIQ֗�9�֦ش�D�[�Ƣ�7���Z.���+��o0P�%�|"�[ņ�
�R6�[�43J�h��9�1�+�=�n4%�/}K�
$���Sy�V�:�U����]�3�׷�/��,W��S�|�<�,��#JV�ڭ&%�v�)Amm$�0��=x�,�(~br�&�4���{Ɩe���T��w�(�%��uZX$	1)�/e)K��a|!�8(dp��:�,������bS|�IYr��8�{|T/fs_1&i%�R"�R*��?"�}Hڮ�-�bKo@���M%DD�����\.��,�g	Y�z��ǖS�_�Do�'�z�W�����P�/y (�������L2��r�Q�q^�|�gf6��991d@�	�h�/ҝ�2���}ެW�"�r)Օ� �jT�ݬ���P9�ֻ�*ݚl��m�ZQ�F��K9N�h5�Y���.�ff������vh�[f���9Ws�n-�]yng/˦��.�P���M�qx���4E��]�7u��VǢ�`�c���ۓs��pn�7�;a�q�2�I��l���nȶ;j��Msa�Z���89�ϻT�NɃb	�;��|FA�;X���۞)MnU������1�}�g���/\;�ɧ����r�jݍ��%��\���]ħ:�]{I��t�[땇��kv�S���'Opv�g�S;���½�f��Xl�mC�{n�Y�_+��D�\tA(\�������]"�ȺB���_�x�%�k��EBJj�/O�U����篵����Ia	��̯u�����/EHD{��zH�I�1M7SKZ(���B��E��x �M7UX8��崟�:Ƒ���,,B�5�"�r�h9�bJyɈ�%�iIwى8m�8��R�+󄨊�;��0�}�>�3N���K���J�5$��N��4J����f������ ���;��``fi�����TB�+�]E��ݨ�l�%�qc�~2s�{��g�'HL�c�������dh��D�N:�X�ՉA�e鐰�ʹ��,���B�w;�*n�TJ:we���u��W�Ϯw����w���F�j���x�KG-C#D��1�V`�&G����	)&raL�MA�fx�SB�P��IDL��y��w�ę�C�ޭ����\[K
#�TF
m�)�~V�U�� EQa�-��=��c�	B�]g�\F��B�%"�#=Q������yڍ2�"M�.˕��դ�j.{���\�ep]+7ޛ�Ih��5�+�������=�3O�Ob��D�ZH[�EN�uU?b��	"���)�7nnq'gr:��/G=g���5�d�������)L���>��v�a����j$K��X��7۶\%���#�-PK�y췮�>��"��n�E�@|�T(W�XBUW�;�U��\��%$T�k��_k����G�BSI-���3&�X�I����ŋ�4�rW5��7 H�nﲮ��f�})s�ȍb/�vR|�d�y|/yN�]}����ML�3Ԫ�f�K��'������F��y��N�s<�B�֔H��J!.-w'<�+ִ�*B@�
�^�c��$���/���_�bS^f�>[k{�|��#� ~��m����(�H�!3�q.��Oץ½��(�"������B;��z�`��~���=|�%k������.�%BRx�뼘	F��߷Ŧ��U�J�z	V��Ξ�
�*:;\��KM7�6��*!��꺩۞r �U8V�|\*�KPR�B�"�������W��pX%�h#����W͞S�BK�[]n�K���p�P	*nE���SX�:�����Zڒ�-x��ث_V�9�	���iM� �,����i]sn���y�R��b��S�"*�)2$�|��ݑ�p�%Dy�SL��n,K���itQ�B���BV'��ZV(R<I��{�{�Z]�ViȬ�|��[��5�����CCK�[tj��c1q�8�u�=�$���L��b�p^V�)i�-���j�Z(L�)�%��y�.�K�ʀ�:�}a׻�S���H7�3��N-�����8�/r�K�"�k�<�3boz���_�6�rU�Z+:xP���\xf�n޻Q�̷�[���/<^�G��
�Ӆ��8�4�%��ơPĴdw޽V�.WV5j�����ľ����TG�OwO�g�!a=�R������J@S+A	%Z6����:��_�B>j��h�)�N(I���3�z*F�j�p�IӋ�-��T�Y�@���՛��K򻿢�@/� �YX�����ބ	�[����+��Y�ζv'Q;^����n�i�C�ٮ��w�m�X�*����Q]���#b���fN�Ė�%�{��҉�e	%nʱ(�X��'N?&�O�|�d��3ʽ�2�ܾ+K�k��@�R�Y(�#�P���U��\�O�D �u�b�w_��>�Q�i<i�;��.�~�]^�����q���v��tbJJU8g���
v���%r	cr�9��W �$%$&a��5鴖���.��B��~]��;W��v�]X��x0��0�&�Ĺ~��F��JJļd�nnf��ZP%�d�
ķ�+"��+5V��_γ�^�c�
���\S�쯯Aļ���p�ۭ/N�:X�X�Gr/\���anjx���H���,L&���B�yaW�'
�/���j�c3�XЁ[h��eBt�����x]��
b�B��ٵ��8(��%	P�uo���d�U3T�%�C#u�^م���<Z�X�3)�'��k���M�B<�]�6�ĉv�)2,Q}j,���b�{�29��T�ҡR�IO�u\%��s�٪��B���H�(���d��4��.]9���,��vB���]!�ē��Ms��0��D�-�"���r�A
�Ka��q��A�F^ g��x?��Gv�}Y�)Q
ĺ�1$Ԧ����j4��)��:B�Gg�&)R�g"S�9U.���4�D%&��S�^�U:�D)�ˮ�L㌾�e���P����ݍ]��52r���"���BXzd��#��/w�o�[��ч#�`f�{�j�t��N��Hؽ���fd�ي����ѐH,�@�d���w���σ�>>g}�ŚF˩*4�#�3;��!�4��i}��5ѽ��TGDW}����Ғ�ZG��"�]?'�6.sKJ�+ZT$��]�kŨ��*EX�߈�+E���kH�[S
��J����ק�C}/���]�,�v�)\۞2S�՜���j<N�[/c[��C�'v����n�]aٳQM��<&D��b%���w�=VB�D�	1������mn%d*��D��G=�W���;<�\�qE��ՑDX�����%���*)W�\NJ�I%�r�S>^kb�bƾ5���F�{��׊7<z�J*�#5���X�Y.Ͻ��g*dZE�{�+�W.&����R��������&{�Gէ'��/���j��t�V��U�Ĝ�pr�J�p�RI
M��P��y>v�-�
�X���}��-�JH�w��j��#�.	Ug�M�\�XG����b�y�"U^��%b�T�RG�j/�>��9�(�V�le�}��X�է���xG��驊��H��ngU�\9w��5�1�Y
����T%��շ��آ�ɍ�g���M����p�Pa9̻��;� �^{{7����P���?p�)�S�uUJB�9�Y�Q�j�nm�~q�5�V�h�
�C��V�6)�ܺ���J�9���﫤,<(�%Λk�r���E[��|lQJ������m����
|�	]�|�9P�\2�^g'�֏]��_�;��I�/9��=��\��P�P��ݾ�2�^���9b�n���.A��.�>6r]�w�9kg;l!�l���ѓJ�;v^2�s�a�]m�]����b��"�ݼbK��7�[��r��a���9ޥ,[��Gq�g�r�Yq̥stqgv����m�6�۞�:�ڷ]��'C�����=Z81���R/����)�#���l]nr��C�m�1���ݱ��S��r���lu��;�cj���6��Um������Q��и�h�\��NN9[��s����I�jC'v5�n�g#r�VQB�h+^��o*M*ni}�����q"L�7�]��J���dB���Z��_m�0�\������<���]BN�Tmv�\o�ڄȂ�����ƽ��K�huL�*fh�`�0v(�!{�p[��u6e�L���_�[���ip�i	N4�ЬJ�&o��h��������Q��x��d��Z^u��}��ዾ���ԅP��r�tB���R�3KT`� b@�^��Ť�:���4��_\��n.\#��W+��yr�'d������c�2��%?��(P֒�+��
��j�8ÂEYu���E��^ֶ���JZ��Zw-ƶ��U����������	�;Y��%�}���:a*��x�K�Z)8*"���"�}��8LS/S_RXsl.�[��6���pD���2$���t��Ĺ�{��NG*+]R�ыm�:*�L]� ����Yn&�k����R��%�yb�T�үR(��VC"d/{��v蕂^:%Dӄe���
�/8RBY{��������1�5T�#��TBA�<�V��G�;&:�r���	��o��eƽ��$�eR3G�,&.�H�
��}�US�\F9ʚJ���$�T�ݿ+h���+����{�?�Xϟ1[�Q7<�ߧWO
4TB�n�;��֋D��}�iz�}�ﹼވG�!c%D�f��"+.b�(R,#��|Z���'%��Ƹ�Z{a�ݺVp5�iҰE���9�/8N9���Y|8�y.���f��Z\���mv�x��b�{�@�^
��R�=���h���J����,D I2Ĥ��T)��zmO�i�m���K�Un�Z�Sy�o����˩sL�:�.�D�'�R�bS�{����]��'�r��X��̜��޻��������L}�	����ΛO�ҡ�))���o�v��ʎBb�H�E��r,SC�.A�:���F��	Ox^���z�g<xJ���j0^H��)*#�E�w�p�w�I��;�g��C����p�D"\-"ov緪���#<�x���dC�������䃒�Z������-ŏ�������tF���$x�P��{���2��!W/,�}�T,%1*�+��j$� S��/u�M���qzi�A'�����[�"0��ݩ���oeΕBW��"'��	WQ�}�Q�z�3�V`���z�ϫrK��]��n�{�G��權��s��6��<z^�8(��긧��!J"D�J���s�n�~q���~��0���
����.�=ڽX�DN��<)^q(s�IT6�*�t��v���DS2=�J��qB@�;;��|��}�v��\*�!�g8-G���0�<*�|���S�w!,o(e|�|�}���@����-w�R)�?^�_ޢmiuw,���'+���.`�X���!�(�;�-B�b�t�ԉH���s���yQd*���p�j^�T�6����(qoV6��B�7L�{$��Z;hH���Au�h��1mh�тP�GfJ2M��t�.�nW7s=
rv�.w�㸛xt�Cnd5�ē���BX%λ"�<����U�]|O}E"�eVI^/����e����Zk����P��y�� �䠄�P�&�VDs�~-pZ(R%�D�N.G�Viq���0V�e3��ji��?/$���{�_v���R���|h��J���S����Kq5��M*�����%�"zғ"�^p�'�]uSU�l�4�:ΫQp]=��+4Q����(q�8A	��A�R�ޜ�q^ih�EbR%]����sMM)���y���rMXAJ���K�r�ucu=��u�d;Wm�$7Wt��F�����X�l����V�\k�TA����z��2�5�EH�7<Zd>�9���8=����`��Ƣ��:�J��6��k��LE
*�����틆����,2W��$����
�/z�K��ٯv�'M��+"&���MgKF�g�%Y
�L@���`�i�ʀJw%/{wKFd�"1�'��3��oz����{��)��,+�����ϣNtȕ|@��o��鴬W�$T�����"$K}�kǽ�Ӗ�;��k�&�
�(�e�����U����P�bx��l0��I-�ʍ/�ϣm���7��J񊹝�ߺ�\�!]8��M71\s\H�����{4����\�99�˟]��>�[��<^og'8;Щ_ rdԨ�5��8W*���z���A���7�N;���ӏNi��d6�j�<���g��4�-S��,J}�x^B%����+%���*ѷ���h��.��~��կ��[�a�\�מ�K՜�(�(�,����"LF��=~�wXT�GF�<�Wcv=�=�i�PO�I�\A�S$�Ż���3.���4s�f�V��u�&gϭ��u�Ӎ�3���JwdP������+��� �5�T����T��Y���U��X)�zn����%��tY�R�e#+��bƘ/?�]�h��$NK	LZ駼>�q"M�=�5a�&���U�bDb�'e3�%'��]�w��Y�ԋ��f��TE�	Hԗ!ܡK�9)ܯu<�H�f3u1�*I�����/����KM�ݘdu�ջ\�!��P��\⫀�u��B��M��	rvB�S�,ZE]�!\�n����%�\m5יUt31��k�5|{"��Dc{�nSZ��m(9p�6��lKt��Ӽ|M�:���}��귘�L���E��U�k6�,�2�L�?BI$�DG�BI$�DG�	$�J"#��I$�DC��I(���I$�"?�$�IDD~ВI%�BI$�DG�I$�Q�I$�"?�$�IDD�I$����$�IDD8I$����I$�Q�$�IDD�I%��I$�DG���I(���I$�"?P�I%��I%��(+$�k$��8`�+0
 ��d��E���!R�P�R	 D�$(U�EB��	J!E�
�((�( P�V�J�AIW�(�B��B�$"PQJH�"��U$�����)E���@�@�H��R�P(A��@P%.Z��@�
I@��$��1��x��٥'z�x���ݞ�^�C���=m�P;�JT����N�{ť�������Xfwsz���c��:�\�%I��wr��������&�*    �w��A�3^{ ����*�^�=h=���{Czh�=���.�a緽����8������z����.w��w�w����7=�=��������T
 �@	ǄE��
R*EE
-�^m�{���7v�/=ݽ��gww��Ҽ;��{���wZ���{��iw�u�Z{w�a���n��\u���m�;�A,�۽�{[wn�n3v֣Mh  s��{���C�Ǖ:�u�ހ�r������W��k�<��P�)޻������8��4q�*�w�J�޻��wm�:�ؓc�oz�-���m�gn��   <�*�U)U"@R�HT�=��7�im&ǎSNV�ޔ��+�w��&�=Q�Ҧ�{��wqt�]��vX9��z�\��U���w��xw��O=�x&ڗ���S��� ��;�  x��δhhP��	  f�м�=  
�� h"���  �q @ �'@�T� @ P =�@�*�DQPT��  f��4�� w� =� P��` gp�����`Љ�i� oX �1
 
`�` �@�y     @y�r��绯mSDx ����'q��MW���=kH�������׻*�GF���T���ݖ��[swa�@
 
]�U�"�EEBTQW��(�Y��V�m��;�XK��&�����Z���^��K�y�Oh�w[c�f�=�Ͷ�Z��s�u����D��Zeiw����� � Ft =�  - @ q�)B< ��� � �`���iޱA�����Q"V�����[��u����9G�6�gyoy�j���={m�� �~�R� 0��$�H�2 `!�&�O2�T�� �'�T�SOi#FLL!	J�H ��O�����������z2;[���Rt�,�]�_a���ଃ��@(
��U[΁cq��UP���P����UT*�����U�@UU
� U
@UPϿ>H�}���F#�27a�,QNC��	�9f�S�kQv7qʲ���eG%��m% � 7q�%:�,1�&2���z��P�6)ː���n[4�42���T􊛿0?��̒=�Cݙ�+d� lgmy���y��B�L��u��s24�eaB�Pw:=�>߭om��Y�ުP�/r�N�(u������Q�=S,_Ӑ��&���0�׀ �f��2̓%�oaj[Hhgw�w�b�J֓Z-L
�/"3��BhYX2��P���eȆ�����R��8��N֌��)�{��д��P�Z[ X��n�ċf����V�3p<�4  Fs.хXq.ji!�e��ۙ5;���#��cm�R�<0�G��ay1�1��nx6�-;��q���1��c3�����{Lc����-Fv�O������ø��v���sv���f���.@F�q��|naR'i*�9��N-Eb�F��h�����V���b��S!7oChU�J�����z����C��6���k.+�#�N��n8�7���1�Ӻ�"ֻO2��3႙ڬ̐��S'��{��L6����%ެ�!�j	W��#.;��b�e,���$�u`�:7l�f�>ŋ\�/T)�ߥ��н��R؎�T�q��nAgpZ�[�'����^�R�p�7��Ln ,QÏr1�);Y����R������I��4����q���tm�:aM�[/1�f8
��jf0�]޻�e�*y�Q��ܤfm��f�S,�Ლ5fk�4q#7Ŕ�ʷ�Vfn��-���B�κ8ibB��&�L�i�MT�w$:�,��W�y���F�V=��vtKÂZ�"�P��yӂQ�_��ی�s�
Rc�D3/R9[tM=q��*ΰt[2���(����@�{z�H�ǚ�Kj+W��A��4'������;� ͦ�K+n�EL�X��rL�uJB����N�S�2
e'�6�����V[��k�:��, �-�F"@d`Ssj�)��/�V)L0�Ċ5a�f����m4��\|ds� �;�mKwɣ�hx4��M���;�7a�c�(�3&<�d�GdW���5��帐��H�8<���0�,K�"d�sFJa�;�,��.�Q�;�t(9Y��S�j6�֔�	Uux��S�$����A�v!��l���J��S)�F��Hۇ/kf,KJ��V�ۖLϚ�y�Oʲ
'v;{����&J�W�k���gch�-]�$�e�6��̘0�;XN���3�7�zb�3��Ɋǂ�x��;�kL�0ꢵ�o�Pi+��vp-�$M�Tݴb�v��"��c�,&���K��hXen��#x�r��Vw(��W���v�x� ��O��،��֜nK��͵`�ť`$��aRD&�=�x�T͵)�݆��R{�����pXʁ�o�B[����u��s�A4������b<��7B��CdZ�
�h�����W#�����5��Z�5T�xZڶ��ݱ5��̧�ճ���֡�"^�yr�cB��֜�+4���n2�%3pQ%�YF*l���Ś���Z3_f��WR۲i�wZA3;6p	�A��M=�s������Ls�
�VM�U�f+�}�,��.�mb��Ow�֪b�m����A�RL�WF]��G�%I,Q�t�����xj���k�!X�Nk�·����zo'6�#�P��mt���g0����v�Uo �x��ej��Yw��+v��M�
���Q3Rʱ
�6񱬪�w���$�6��r�����d�������ÜD�rVͧd�(-�v��ۇX "�7I:�F	���cr�p�3��cA���d:��:����"d�����(��eU�2�;bK�p���r��{��!%��-{����EY"��J�[�����ɂ�`yV��`lf��#���j\��ޜ��@��C���;9v*L���3CJ�s�n����*k^m��üj�q�u�xj-�̣�����'D�ee	HЄ�M��֭�m�;�"I�kUdc��Q܆���XD;�x�#��0���"m7��rA���9�b�8�^�J˱�R)��]��֫nK��P��iS2Gs��u��J���\47[;-�>ѹVj��PX�U���p��Y�[;h��.�,�؃$:dٖU��{��ā*,�<�b�i��13Õ�$"��3x���L�nh2� ��r�T06�� C�l8�ΫT�]�a�
bl�7t,��ӂ=�қ�I�G�Д�i��cTom�Z��sܧ0�̸g�U���j����|�R>Gju�u��4�pCɎd��G��9F�ژʚ��-�%4���l�2��R��W���/#�CP-�Q�[�H^�҅���W0<��ڂѱ�AZ�
rɖP��H{$�\<Wc6�I�b����NqE-��#�0obr)2s6R���=�Ŷ/3Zi����X[B�l��%k^�>���-�F޹�U)���M���i�����F��H�wP���d�yxV�wk
�������{̜�q�y�M�&���U��L�e[�%���2]h,f��U�N�#0��i��ҭm�3�o4&�gG''0�C�O	#��<ǖw�.U���A"��c�Y{��fL+%�a*�� ����wmm�H�U�0B����m�]G<�;�;��Hi[q��[o3Q?:W���¦��y��kF`k-�KnJkbf�P���e,(!�s-�!�u�]n�TbQ�z4Vf�Hv�B�ic�]�^.i)�6_3-j�&�Y2=m@�ő>.*�g8d�e͈2Op��4���l��gC�'p�32��e���m<ܷ��fr7K`Y�Zs��8f3�j��o�h*X�+F)4�qm,��2D4�Ne�oaX��ޕ/h쫎�"�e���Ed����F��q�	XJ�ɭ���W���T�y��/��`D���NC(�I��e��|����l=��̬	��^T͐ѭ)��{en]lV��
wQ� P��f�'e�io�x*�hG�D֌�Ȇ����Sf�P��l�ʱc (XA^�h�s7�Ѡ�e���W�7�R6��^V�º)�h� �����L�.fۥRXL�2$�%�ũ�1WK뱩�	SC�.��7j�E�u��A��1����n'��K�[����j�J��үZ�{�i��YgR�@][9�귆��لm	P��i�b�%��+�ۢ�i]�!�3t�a&���0������#Z�s�U��^�&9omm+)ʭ2�(�Y#�M]L�o][[)SX���ˌ�+��e��,`�kCQV�"�ZM�,2�to$.4�2�Ky��	W�-`:8�B��9�e7w�CqYz��h�Bv%�c0"&�xsPVod�[>4ƒ+
��W@��k1�bi��6_ӨN\�{�	�x ͱ��QS��bX�+EnaD_�����$l��|kmM��㩊m^�6�GW�0��Y?�T�Y�!��u�̖��A���XMR�k�*n� ����d�<W���e�n�@�I�:ɖ����sڎ��&�4w%�ɁY�w)�v���X�#�*��C��,,w����Y�8���g9R�p�;��FN�yl����x{�A���,�:g1�|��w��c���ޡ.:��U�8Uv�$|������}g[�#���K������]��B�Z�b[u�*�hwHU�n��&��Ǐ�Ï�Ҭ}�Sv��=Ck{4ŗ%۫\�u���T-�:mQ}`4�;ҹ7��9/I�b/��2.���=�^�'j58�X ��S�1�Gz�\�@! #A��o3w��f��8V���z[��m�Rǫm[�x�{���R�Z��[R��S,��G��2^�L����TZe�ͣF2�6h�%��ceԴvb�qj[��spf�Q��Tc���a����o@7�UdL�n�o��CZi�iK�P�y[�J�I8�]���,�q��Y�4*u	�r�[b54��4�������^$aⰋv�Ap̝k�	3�{��cy���e�ݺ�VeAN�扗 L\̨M�M�˨f���cwn�Gb[��d]l� WEj!+O&�'q���#mf�ue��o���-�q�n����0/x#�m�d��өB�r]��I#�-r�b�yl���=R[���0 ΍ƞ�,D樲�f2�E��w�+J������SX٘��t�o[�k[���n[!�ff�``5�XZ
R��k��b����3X"�`� z�;
��u�/V��E+TiҸ/2�7j]����8S���[fn��
5HK�]��؞�ik4�+t�M�
�ƫlV��{&ޔ�b��B�Cn"Q���v:U$�Z���y.��I��B�����6h��b�p�l��kPFd�P�hY�,��wm�jXT�
��;b���h:g$���T��=���LV��.^�@=LŸ�%�n^S2�й����kR*�J�c�3Y���]��fX,�m�r0�1-�6n��-i6����\��!sJTs6���I�47���u��/\�ł�Ӓ��ר���v$ӎ�3�ǆi������z*���8&=�������XB7�\��7L�{�f���.Ӊe%x�n�R٣����j+�lW�9�n�31J�$�d�)Ӧ�$e�w���]�lj��ߍ�S�k���&FɆ��6Ϋh�n�j�x�k|EFr�f9�U�F�����ȖL�m�y,;���̖�e�򒳴�,���yz�K�M�r��v� �#e�L�r2P��+ɑK������ws��a�2�Y[.� {�b;cJ��e:��w×ISP��D�ַlj%Dn�.� ٙXHѸ�&�J�@�:GKD�,�J˸FY�����D��G5�n��xiA�E�U�.l�&&�\�Dwvq�d�(�֍�P^h��{�@R����%-q�Z��hT�	�
]�X�s6��vp�j�K;vU<�##��V�0:�.V<JQٷ��#&��9Y��J֗��B3˙�;Z��������;1��.����K�[m
]3!�(�+d�����GN�kK��MV��M�al+5���-o1e���Mi����nXM!� � ��&�a���5�EW%0oX�ֲ�ѳ\*`Ĺ�!�é눗��KѢ���5XA� ���DR���S���Y���M�̎�O10%'zF�f�nj,�ˬ�2i݈a{��w���|$�n��R�! �f�E�'J��
m��5eʅŵ�v��e�Yw0�e4iR�4���Vh��K�qlWzm0��nfK��`V�pL�uw��d��u3�t�T-$�`:%�ݢ�*d,3)6r�jJ�n;:.���f��Ǜy���]� [��̥�)c2=���"L�ojemǂ��bRt]�Y�aB���E�J��i��83�� ����'��৮���X�&����,Y�Gr��˶[j�V|�h�u)\E���j�CQ�5}�McԄP�'�%�Y%��w�:�Db�Ba���ؼ��"/y�xa7�m�0^�����M�fK����8�J2�J���1������۷XB6��4��t?���Nw &��{��h�0�YVkb��V�6ⶰq�֌�8����Ø�W�f�eVYJ�:��Pd�CK�,�X������	<���9�zI�I!��I3#�l6Q�CeK�vm�ѵ*��[4�֪(iU�6�[�ݤ��2F��|��%�Y8L*��s[9â����eJ�M��.��J�^a��c��;�P\)zy}_���L��{��n	�OXs	�n�!�]��� ޖ��.H��98.�FZ25�w���	�w[�5{��S��@��	4��$�C���|�R��L7i;�����дl��>;fl	6��2�U����
��{���F��"�c�i��%�b��E�+M�x$�$9�`�<�C�v��E0�{��0/��dJ


��G�&�!�nV��$��XWa�8��\8bY�R�	�,���p�SN���bƛW+�Y3��K��W���-<쏋-a��"�CI:����c%��,�j��F'A//��d��G'.��U�

��˿���W�A>(f[�(��U�M";Y�n�J@��n�i_d��
��$�;F:4�G�t��SC��ڄ�NU������c�-
��e:xN��XT0���1t�p]棛v��R�j&�iMA\b�i?m�+��̈́�NH�<���"���B�k=;2�^J1LVl���p�c�"�QVʗ�P�6]�B`�\͙A@i�m�n�o�:_^'.�E�,'����I���A8��8M*�$X����P�͵Ch�^��vAl���Y˨]�,%Y�6�GO/�\��a-6�7��Hs�R�AM"� �Y�jҸd�ʶ��[V�op�çc3d�R��ljƮ�Ӳ�F�Ly����6`����+r����@���#/�Q%�Šhk,L�����V�h ����vmJ<e���x\Ⅱ56��s6Y�L{�jj�s++l�cP�nT�([d��C��{��q^	Cov�Y�'G ���ʶ˘���6#��B�;�N�\׸͂��1�r�x��	I�x��iW��ON�R�Ռ�Y�Yxd�P��tn�%�u���֖�Ͱ�2�2�\d�� qe���eL��T�dɰ#�c)
ʄ�f��,�N�R�*�/�۹���N�����9�st��!�价��I�`r�Xn���^���,דfZ�p�ӏvi���C-�Ad��C�,�wnLxq���,C����3SY4b��^x]�_-�����GV����e�eUL���U�j�����YUӷd��j��XՔ���
���W.Wcav�6b�
�	��N�k���۟8}����mO��{l�W'5<�����U�g����㧵�a1��:�m�@,�,<�v�݈�pm���]��#5���z�<t,|%��QE��s�+��Yϛ���,r��N!��n�n�*��	v��n90��9�Z-g���	�b���Ѿ���u�py8���)q[t�=Wm�˳M�q)�Z�la�V��\���8,��6���Aq�uk���듬/	���"�tZ��~끸�uMQ�k��-q���y���\r��JwNÁ덮KvzM�6ں�9)λx{Rr�i���ͳtA�[�u+!����gg�\�D�ti��.����	���dM���V[+,t���5rw[��ގ)�s���W�%tq)v��Z��ł#5iy��l��q��[���\%s�k۵t��{%�A��&�1�nq�֟7j��[<zxؽ�B��l�H�2�e��8��̷c`�[="O>w\���ɾ_�sI����[�vq'�`)0v:v��b�v��6��<�y�.r�!\ܴc�\ �����ƌ5�f���\�ծ��n;"�sf9�6�ysۖ}����v�\ә�[̦v�/�NR5�%3Ur��%c�ħ%vś$`�%l�}����\���!P Ÿl��n��O�[\�\� M�����Ъ��/Ca$����R�w�����&\�1ٞ��ζԡ��d�t��Kf�tEkF�X��]��}Y���G[��d���НWjB����v��F���Ҿy��˨��y��;��*ۃ4+u��� �.H���;7� mq�3���I�Uf��'/-�	A6�l.�\��M�o
���029�v�K�۶629 ���Cs��z0��1n� g]4s+f�m�[l���W�s��+�18����r�T�{���ɴ àV�\���ɈES7m���3��Av�71��e���خ�|����ɑ�m]�WAŕ4�1���撙��][FC���Hv���N���'Sǲ��Y[�qcK��^�V�w+����11q�׃����lB���˸�m67���.�t�{a�;w>{F����W���K3e)a�� L�!uq��E�<F���q�{`�vqѼ�K����oU"�\��.�+l�%G;h�C&�m�nGr�f]b��J̖�˷yN�綥h��mas�Dny��=�ǐ�0�ϸ��2��`A�]�Ô �hF0r&2YX��h8��;��E�k�̾�'��2���<[�3���e�@(�C�{b�ls����n�s`�k"f��1��l��X����ch�ō%��)�u\X�Q�u�={����ùcG����S�y�[>$�ݪ�:���c��}�q��э��-�s��2ń)��]R���i����I�����zώ�[���ku	�Z�re6z1�*�iP.E�2���RX2�YK�mr�Z�,�w.�Klm
��5��\<�.Ajf�	�B�mŭ���ZYa�s-��c��]p���Sؒ�/q��]��Q�Q�<˼zK��R�ZK���RE��k�j�	�!�{p�������Дf֢ĊL()������ԛ�5�0lO\���b�It���h�X��+����c�7�ΙS�B�+Ib��Z59.��a���\��Ƽt<��'up��1<�xܬh9^ aĭ���7]q��N���$"-k��k)4*
J����V�����8�lNtb�[��;��;�7X���,bKw.pk���'(�	�σ��[�����& +dk�4[��&�t�@�7�踥c����mIUkĨa�Q�� 6г���dm�':��x��熞���6����9ܧ��<-�C��F8/���(��9���f1�۠�؞�<[%9{/Yꎽ�h4�:�Cgj��!*��@��e����)2�j�#��q$��S�A��ǧ�'/n\��v۶E �(�"��,�)�:��'#�ub3�k�O�c�p�ɣ���h.��Y�-���g<�l�lc#���Q8�|�m���B��3�Kta�3-����#�b�e�6�4Θ8��V��9��9ۮ�<�u��ܹ���%�a-c`J�b��4dc�:s<m�(P�9����WhT8JV}�1'�Fݟ!�v�����df�G�� pkX\�E�c]ζ���I�&�)X�;N��w7<r��[1�(�(����a�yw��8����3`f�u�J��ښ9
:غ���5\�u�ݺIug�����k��x���)΋��Q���t���k|&��4`�嫅�&Z�sX�]� �T.�
r3��mepd�sۣ������Q��x��g&�Ɠj�h�mm$��Q�V�٬�F�@U�r�VV��X���4�vf0�������M�r�=���^ێ��a{;xU��r�z��g<��lq���iͳ��M5��(r�!$�#�v��D�'�g�Xp\Q���=x�uhK�xS��c�d�hC\��#�evа�rf]3Q���N)�7d�7<f1�sƲ�o}���)��]�Kٴev;kg���ջp��7Z�m�f;+��Mg�olp�wc\
$������� �k%��ϗ����kz=�C�;zܣ�Ѫ7W�\���ȵA	[2��nxq�s���l[ki6�LU�m�-���������[�MVј*ݙnF�"4�c�y��\��O,���4K����-�kPC�pX�^X5���n��;��Mt9l���k��0��$��b�*qon�I˸��m{(��L�q�F�v�D�l����ʪ�:�s�R��]n�6�\���-n|Dj������D��֭���R@�)DV&��:�۟ �R�ɮ|k�E�ɖ���%B�U�����|���J�n8w[lm�s0f����TjJ�K+T�me��q-�q��4���\�iq��k��ݻ`����;�=�Qެ�H��]��2@v�����F�D����gs�m��0C�K<aN��CWWn���`37&�qW��6�<��4��!�k#�^<�ʤ5���븍�\�K�a"B�5U�{v[sͺ�@����^[`l�x�G��㶗�v��un��R�Z��yu��6�Qǘ����������z��vs�\�������C�mƺ,;FC��>y�b�WB�;Mp����m����j��v�trEӅ����{�3�,m��[�8�5[<\b�nf�����4R[�E�RV��0�H���26$�-����cX����fe�f+���C�R�ݷ--[�B����(@�X�Ֆ��au)�wt�pqO�x��cn(�w��vɹ-0XO9k�h�,6�uތx�޸����;z��p�w�eB��:��솲�k�<֒0D��ˊ�y�%�5Θ�m�7b�*8o3��ҫ�Y�����J�X�b*��@VMl�;r�/c�el�X٦�竌�v}�$�/���v7>�4�q��B�HA����de��4MbU�(�cm�IH�m��t�a�ٖ��k�÷������<���nSk7�wh�(���A^����8��n��C�e+ؐ��/��fY�Fg�:mlq����h�����e��%&�s����iv�q\�,"�.�y�w�3/c� ���E+��{��ۺR��WE�� ,/&v���9�h�&���݋tu�^= od����P��,�&�6�ʗ�.% �:�ds�����
x:<�z�wUF���V�a�(���
�6�=����¥�hН��CHX�-f1�n"j��K��)f�qeؗt��v��f�:�5�=���#gp8�S�y���GKSf��4��^b�M�mؗm*��!���o��(�n:���:��wʫ�YR�ۛ��on�Y岓n]Ĕ�8�K#4�o	�t�%�u�c�m����]��[��5����<����l1�spVY	�o��M�D>v���C���,tz��ۥ�'vW9�!����W2Y#�gݮ��7�bۚ��r�(CC%�0�S���v����8�y����s���{vt�(�9�f,k��>Ӝ�e{%��8<]1�Ǧ���xp���j�n�]�t���ӎv6gvN$��ԝ�U�9�$r�'O:��f-���
aL9c�v�v��8�Ӯf!���b�Yff�Ep�&�k���^�ϊ���%�hw��цK�i��A��C��fel*��Wjכ,Ukk����Ic��i#�Zq����,�e�1��RA�u�ն\e�	/��&
�˰��3[�����Y;]�=�g�4(�d�eg�
:H���s�����3�9�\�Jx�t�=���
��d䝞nFS��mv8gps�a���JB��Rִ��
Rf�+tcn��x���,��Vã7}�=*� �@p/,�����36��5U��b�ZJ�]� nv�3$j.��b�a����l<��-�9�՜�M;u���vpB�ѥ�v��[G��M"���68F��������06���-,f����ySi�68�ե-�Y��;u�^nF�i�^Ϭ꼖�]����f���,y�u���%�:���v��7od�D�k�;a�Y����4,u�t-ձ�j�@��r=�܊�a.Y;N{ٵ�fLm�wi�Gl\�C�i6ݍ%�x�9Df��B��㓸�׷l��q+͟n����6�ŻL�^��b�u�Mn�ւ��M\�4-sfAGA������]�I�l�	ګ��;�I8����\[ە����|�v���l�F�Щp�aる�9 v\�H�T(l:�{"�������̝��k\kR۵\���ct��34	��3	�]l����G��e�WcF/5F$\^��K�q2l6+�NaMe��ά걚h��c�H$�lh1�]-6�bkH�k���W�qc��U���T(UUC��UUUPU��@UU
� U*Q�XVěR$̑�ۛiqm&�m���ִ������\�k��q�ĖH䣝�}��؃WXtq�g�żV�L6m*��`��͓����/n��,q6��\A���Y�e�3����W��R���奻������i
�K���.4�v�z{V���1��g6��Nք`�����B���.���Dì�e.ef��#ff�}vļ�9$�z�P��ŮRT�<�@�Q��&�Pf���)S��p'���7`݇w\w�`�gͶ���	�y�lfu���c&3
s��͓ٮ^#�r��.1c�n�Ųtu�M�ϬY��5{O`���.�7ae�`F����VY�tj��b�@!�x���E1�8Q��L�����nlea����v��M&���O ��mY.�CK�C��k�bf.���L�۝�m�Iڤ�2q���S�M,4��X;j�]]t.�K���mCäG��m���m�=b����úćn��vnn����s7I�[R�����Ç�]�0fzۭ���8'j��Xu�5���&X^͔E�a��MK0bX�&ղ�n�L.%��/���:��L(�n	no[O���60'nK$uрɘ��sƞ]�/Aͷ�Ŕ��j,#V�lPkz7B@u�l�0!y�.�ګ01ى�sR(�3k��ˌ,ko����ؕ���{h�p���Ǧ���z�e��4e��qrVi���A�@�&sk\ʹ������b�qd՜�ל�b�`��[E�k�;r
�
�VӎP�6+l3�M�pBL�p��re�����*E����{p\U
cK�d��-+��z���>�O/=���wN훨�f���zof�ρ�:����'+���1���ۅ��m�ɵv{�apd�=f�Q
��rӚ����@��y:.@�n�#�qہ�4����)e���\L�
���K\%����j뭞��yK؜6]�s3�x�ґ�T�a�f֨.�I  �#B��$T5UUTMUUP�(P� ���&�� 
��  MB�I9Np���*�]�YR�����Vu�ogB�J�aѷ"�G=d��Z�p�֓&㗬,<&1�7��k�8a��Sh�-b�pe��8�r(7Z�J(p��/B��k<��:���|�'Ú�i7u�l�����Y6��h[(�B�ieB�Z�DКM5�1�u��Mt�q���8^�Q��� �r�G�C��!�k�u M1V;0�rk�;��k� �뎣�psHtS楗���''\(�����M6h����n���pa_�k�W�;��'oHј�޽ɠ��<_L9�Y��$R~ճ���6�]ď4@d6��IL8g�;���R�Usss�K�6gFQE�!��+��y�xu�p�w�}�Aw�Z&��t��������i�MHRr+�4��wwξ�/-䝈��Ħ�s+�4+�^N��vv�>� Io�(�@��-���`^3֫�sT�5�4H�4pH �{ʘt7{v���v�=��$�p�w�-:�� \�tkO��{�{�O2�Ӯ����>%t�:���y��vb�c2���r�u1���tͲض��+�b�[���Qv�u�D�f��p��(MH���F咶S05Si:y�D�۝�J�		QB�yr��>�)鿋}��{l�$!1'�V|p�?\��6͉��FU�l�͛�@/r˒6ې&����^���V_e�7�jW�iely���.��Ȑj��8�i�{��1�ѫ_R�3o-�(!<#���4^JUk;3�_'��e��X��8D0���u��C �SI����҉�Yb���u���yW��mo�;��}̸��2�R
q�o9}����}�;@Ge�G��1g�z�co��R�tV��;��묱8��/��R���� i�`)����)N�3OQA�ܲk
��o��Ե�����kI;q�ǔ3��T�����k��/��%�Z;�#$�l�(�"-ɗ;@�_;�ӄ���z:;:��i-�/���@�l��T����Q��Y�ēw��'�����,+�kb�� U��U�\V�uvv���|�Fk�2�Bf0v�n�j	�X4 v&.K��sS�X�����/j���X� ӝ�iv�-���������nn׬(���0����n4��B[�Y�8^s���#���ކth�4�O�o��k�
|����(����v{�쿰`v�ܾ�E�^�J���'zK�u�"m�:��Ž>{�/g�\�C�ڊ�]6`அ��ճ7�G"c�p��CGNYXE��`�� �<7��6mwѭ��y�6��.�5����1_+O#�k�7�����6.�o+��!K]�{�-�����y��3�[w�}աe������B��L˱�D|,1��bސ��|ZQ��n�b�6o�ܧ�ސ.���^>�UK���έ�V..h\8]Z��y���ցs�W\7���Vg����U����bFlǻB:9NG�l���.Ѭ7���%���j:�ox,a�i:��<�7/�<IB�R�,�	�����/d@)m�αz��	�J�c1
�X\걂@���LF)���`^���gq^��"۷`��&F�b`@�n�E�k�}Y��_+K!kd�����4�d3,����;v�`�j�Õ:��:���\���Dx׆�6���B��ѥ~,�k�;��̘L�P�|�����K�&D����ު�s[��#�*I��P���\s��w�v�Z�{��w�:
C5����4�!l����ᾘ�C�rl���$F缼�>Q�R�($nZ��C�l��坵&?D���[0���ukZ!�d�[�(���|���x!�m�fΛ�b�w]�y���]�Û�yK�mU�d����Z5��b�H��uJ�k�3p������ރ9��]�}�F���ћ�Gv:RQ��Aq՝n��ח��Ӻ@�ҽ�vl}ɬ�T��f�̠Y�m������Ko.� �ޮva��⳽�-�9y��z�eXi���ZK�d�7�5��n�N�3�r�h��93c c`jHT�s��5�6���۶f��eE��{��j"���B�}��[�-]�(��n\�w��&hٓ�U+�u�1t�E��K#�`FCaF҉�+"�,�5�N豻��qZ�hi����V̓B�8W��Z�[����kB��.��{�hu��-) %)r�QĪ���akoA�/Nn���;��`�� ��j+�^+�L��(|������X�л]0��6�c(��"I�[�E)�{�Ə��o�GގVg8����:^K�nI0� ����_]wvQ�ͪ��t���Z	�DVe��^w�2�!"��;؂�G%R9�ː�%t@�u�e�e|H��2�$���=/����k�;����S�kFӉ�~���g5�MQ�}��h���,Nu�����y9����
���b]�V����ն9�����c
�Է���/��.���f��̠��E�]b�,�(�~���;�y|%��&���a80�Z�n���:?����3�����p�x�ⶖbЅ����6�K.f��gl����z�۷���l�ոEc�K��kt+��[�! ���J�1@�M���Iu��-f4&ю��S�]	�EKi�.�ǞVr{uZ��2��X�aRl�ж4�JX��$jDf�����t]=��։�e���l�$�m���4FM�uu���F��Fݡe�Ѳ�v����n����>�'V�C�4)v]E�p1;�OU�?~߼��0l4����n��Y˲rw==،4T����D��8����WW}�mY����!�1ƒ���0) ��:�o�7c����D>Ÿ�����^@��s+�6�������^�b���nV��Fxn���t۪ ���M��-�.���eX"�f&c��pD1��5�s���N�]���Vs��Eo�=I핛�Z�~��O�΃}�`ĖV����=/`ӗlH�C�ԗ�Ɍ%�͍��WIhobᖲ�q6-�����G*XL�3�e4�`�8��$啟�t���QS��.l4K!9���o6�9{�azJ��m$�%8"��%i�+��i��\�b�2��V�C5/S5�'/���S�o8��U��ݚ���wK�vݸ=�d?z�θ$�S����_eE؎�"^/+�m�e���<�nQ�Wu��7.Fa�wl#��E��h�5��n��,l��)��I��{���s6������t쭈5y��ۋ������#�6<��m�Q��Wrq퉋hH�w��c�u-����E�1s��K�ф���9�٠Ãw']��z���=��oS�����4�Jb��Cn�?]ڋ0a#CZ�\���ͺ7KF�xq]aޙ�Hc���?)2�����t��=�����
��^8r���e��j�K����)�Kq��$����n�3�횻�uf�<���r,E��P;�w!%I����R�`�K�7Sow�ڗ�2��n�)�Q�D��	��VΣv2D7����ZT!D 5�b ,�jb�VQ�=��jA�-
�hR1��4l��9��t�]�K��9���3�u�Q�e8�9&Vi�5�@�p�ܓ �����>&t9�sW�NO����r�1��mA�f���oc���T-��,�e��g7ܓ�ȡh@�a&�3�f�M��Pnf�X�;�M�l�;y˞&�!9��g�k��Ӫ����<���^y�g�Nq�
�#��LB�ڠ���Փ��9^k�`kĭ�$�ǆ�qZ��N�n1��Vx��� S��u3f�����i�a��1羹����K%<��{�!�D<o}&�Ke����`�k��%�ϷOۉ�#���^-K�S�Ⱦ%m(�,E)9$���,Ȅ�0ݪc�w��{cԽ�)�ܝ��[{%Cƈ�?F���'�sp�'Q����%bmѢ���;��G��(���[*���f����Ά��e;㕯�"��$)�T��=�+H�H�1on嬬$��;�'�痌�� F�$���8�2��`��������;:�~Y.�dU6�7�7�T��X�]����
����[�_8�Gw�iM��T�^=κ_�5��R:g;,��1t+t3���U �u��OzEN��,Y|3�����"����D$A߳e�!�>�w��͐6S�kf�n��<��gSd�
j��BM-PŃ��z����V��R�6�\+3g7L8<�% �y+�%�8B4�h��ٔ�ͺkp��xo���3���ƀ����HIV9}jXÏ�=��@+��O�!%�di�$Cm�\�nc�w�G�p��\=��Hqzy��b�j����3���	�A��!�%ig�'N�K����oև%�Ab@C��j����\��&�{2h#H����XA����~o��*R�c��7 Ʃt^_	L�H�B�}�b�5STZ�pux�d�&\M�ۃ���\��=�!o;�,Q�B�ηp�lL� `ll�u��m3���w�0�8�;h�G�{Fu,�$��v��l^\�V2�n_WZ�J:�k;�;Wu��l��� �v�`�'�Zm9C-�͝WLh=c.�ة����gW���u����	�:��ΐ�a�!#dd]�N�����SYѭYdvo`=Y�X��� \��c	==�FqC�G�w8הݍ�1��	x�L��/o�C�l�LF1�3j�6�W�K�(��Ύ��ټ�v��m��ut����('��^N�L ]��v��a����=��W|k���~B+6o5=�bL����zdb0�q)��4��D@�
�*�.�w�̝��ΐ�1�-#Vbw�񐩞�9��I�n�)t�;&uޝhsw[{�ۃ%����3."Hm'��ˑ8Ww_M��s����%�!w�9;r���ok|(���\�$T�Έ���m��`Va�EA��z��i0��!"%�/�ҧ��ݲ��CQ�潈_J�zFZ�4J�����Wܝ���ڻoJ� �',���m�%�KC�l��w%����RIe�f�Q��L�!�AF��Y������B�6��������OOz\��"��Yj��SKy�z����O�c�5ww֛��Y���\0��ݘ3ۙ>��Y�Q��_[�RA�S�^�]��y}[�[�Ν�b������Mz3k-��gRq������Gy����D6`��L�K�tr����gt�ک��pS�8Qݤ¨�X��e��Ñc��5��u��U�n�`�P��6��g��i�n �[���f[��58�/,�-���i�ȢU=�/;����'|ݠh��c!2D,*fhZ��b���₄�1ї/ �a^�cӽ�$�l��"��ah88�painc]���p\<�uڞ�;�u�W�b<�jvJ!���Σ�+�Δ�R�׍�1�;Ys]����,�<���c|���+3!b���iԇ;�]]�]XH^?!���w�,o�AGH�`]��R��W�����2��}uX�XEhe����[�v����Yε�YW���O[�웛*A�H�4;�zU�y	��j��:�f�쾙Ȳ��\�׷�=x>U���Z�H��U��ky��8�|а��4�$�^_ʯ���V*{�ٽ]Q��1��B���f�9�US�w�T�ӻ�m�����j-���ޱ���a�FL1^�0)g���K�m�p��4�[�Ax����ᗓ��\(���OY+�[y��;ܭ4���8��׿=ச�]@Fo/���z��0�������U���K9���I����In�v��J�T��h��wU������y�r������v��`Ð�=��'7�Gg�]�[��s��:ٍ�&vp�Z�dq�t�,�����k�=ɸ�@�|v�kߍ�����;F�M�y��WwL�%5P���H�dv*u�`~&�Q��InK�CZs�C�/��f��=|��1*���۬�*���WiAtN��&��ֹ@Tֶ��Y�b�B`��'.��b���2�#���v��M��n���Q�;�o�]���۾��3��B!]��Y�ZA^��͙��7z�{���}!�����$��Y�Jj��nŁ��4&v���Di���{ ٔ��i・z_V��iriW.���#S���糒ץE؃$���,�n S%0�RM�bF����b�_5\��b�n��/�;��'���$_��L۟m�B���e����]/#���I5��S}��Bc�u\k��)L��C;���w�cj
�{<Y8'xb�a��� '�|�jh�u��5C#��a!di��L��0�6�y�~��JN�pZG����w0���#�YyDμ�X���"-�M���s�Jq�!����B�0�4�9�ش�P�i�y��9�aj�D���@.N�g%�ϼ�+*�5N���c��
������NT��Tr,<�;�����7���ԨDM�T������i�3�n�A����Umr'��������ԕ�t��s�1�;ݠ��zc{{�b��. ӑ����An���T�k��ӿ�����3;�\�&�v��M��$WsX��X�÷�O�$,�sgsYۢ+̚�勝d�#��Ye��ʸ�˧o&���.��*������z�e��Gqˬ��$�������o���d�2m��/*�"���5�}�P�Őг8G��Cv�L��}fi�!��5r�k��5��6,�Cokb�ݦ�H�ʹ�R��S|Y���-�� Z̊>��՜j�@�]ٺx��}ٱ��o ��CU�C
��w!`r2�3em^hv��;��C�U��eI]�n�".�+�l;b�I .�aW��zi;0�3{��y�<��L��j��jֹg'��f�R�.����Y0e�.�ſ)�^���o+jD�*h��bt����]>�mYK'����90�*�{�T3a�����U��6�N̈́���f�E���n�������FVVe>�ȆJ�j�xZt����VR�`4��Ga]�(]�կd^���Yϙ�θ���Z�h���Ų]I{O��f��v��ƈ��}^Ws,o� k��\�qKYATp�VIUc����K4pL��А�ڲ]n��]ѻ���:�ǔ'v���Q���<��������@�Y*�싡ݣ��=���o8��JM����9t���OOq$��E���=�i���
5���[���-�53mь,�SMM�r�۳{P��.�\���OU���]��]��VXypX9R��(�)V:��� ����N�+���c{:��@��X�;����Y���n��.�5�s@�޽�&�Z��s�'0e�1�3\�潚�{Ά:�?������g=vt�!]�tS<�EII��\���gu���l��7���:�ԾqM��;�a����d=�`I�,��I��V�^�!���r	��͋�jiyK�a��
�I�c��O�CGł��݆E��ʳ����l7�r�vg��&�;�� @���g��X}c=�#y�lكH��"h�����3�7'�Af4!�P���y5�xpn�@��xe�@v�e��r���ƭ�#$m�ۄ�*)$Q$-A��Oeff+����H~w�٢>}�ԙ�|�~�g��M;�Q��6G�^f������Tm��J#E�7y�	96��/�c��jom�!n<���W�u͆v�2��"�W2��V�M�=�Y�_:fpo��@��ݷ�0Z%��ȂJIEF��B�.���#��7�!�+(�M?+�{�S��%�%٤F��;��`CA��س�M�:�G�wt{�@�%���k�ZOv���z*��|2n�Ya�����U4��PT�w}�K0`����ӑ��wN���K��_[���9a��M
8�2�G�{ .�o���y�5�啜����ۋy'�wzY�Y�Ֆ��kx4��Zf�d0y}�C�ƣE�r5W�f����9�����+7��e#�v�9J/��賚Kش�L$�x�0�i����{��|�a:�]��-An]T��K�:�kJ���ʻX�q������z�7�n���m٤�%8Ҏ��r�ʃ50�2��#�-U��7�sL4�M.���hi����#Z�n����a�u����0Ә����qٕH��]7������%�¢��qX���C5^븀��3
q>��WY�n��nv'3����p�gO5#Xy2^`��i��i�Q�QH9���Ub��*L��l�Z?!h�0lr��n��/ʏ�k�[�w�H�J�l&n�_��﷦�F�h28Gge�8s�y��.1�9�������vt�c�w�2�,4����y`��x�t��������������6#�ب���fsAnJ�;�t��Xw�=��/��i����]q�|�1���d�)f#��> ���\w�4w��!D��Z��~��ݑ{^�Oea�=�'T�\��قv����c���☨^t�^���D�[wNl�ʸd��Οv���� �ج�ٻV�o�|r\�{߄��6�iurV��]����fu��0�u��a�jP�u�t���	�.��r����1�,E֮ �r�T��dw���n'�91�m��q���bҋ��p��	�#t]m��<٣HYc���p]ណC��q��c+�s:��b��ff#v[t������.�o�rn�OW�ػ5339�k�@6,+��a�Yp�b=-!�;s��c�N�s�X��e��lR�0�.�����θ�k��\i�ݤ�\�#p�!�L�";�Ƃ_G~�������h��孞n����v!��������֐��&�Ʋ�􆥪7���hD�PE�"Q�"�� rz܉U�wλ<5	�a�����x52:�e;|�/{y�!<�ZG��������]V,���ԣ�K1rvݦ�%'%7rE[a��:���0x�i�lm��#V�4+�pVM� ��l�n(6o82ep��8FZ���������"EF��r������D����L��g��6�C�oWx6���d�j����K�J��'�=�ośCo���+K�MM�����'��aXFݗY�I����yR�̬3�o�.��a��ݾ}��7j٨6���3:� [�qSaYO5-��ǺF�G�Cx�l�(� ���eZiR< ف4��W� �7�U��v'���y��%G3Ap�=�v{Jw�:�����&56D;���u�Fj�vj�zz#z|��fv}L_>͜��9)�w��`�xߍֽ6�1r���Vͼ�`v.Tiz����	����4��C��K�>�b��YI̝�ʑ-�-SE��g��2�muM�盇4]�9Nh���VwQ�Rt�O��b�}�s��ot�}������Ѓ5m�/�O�+�zf���10g7�X���g��۽�3C�[:�A�3����#4&�\b�{h�Z##AK���Wp?)C�8��u���cZ���8��(�[L�7|�^{�=b|���D�(� (�
��Y8y9���3I��y���v�K '����:��  n{r������ܿ����uC�y*�CT��E�B$�"�ބ�̓��%�!���hR\��ʳ^><ݒO�'�He��	�Z*띠O�S��7]D$�L�\K�YD#�o/�,a��?5e�^]=�7��&���Q�61��ls�b«�n.�Y^K@�s�\%-�Vb:��\C*\;Ct*�:�o:�qAULn��e�<�3�=�((q�|�C���*x�2ݝ���c]M�K�����a#N�6�3��\��#�"���YH7k��d	i�Vsy��e\�n�1&Zu�:����n�1RU@�?�#Lj�u��M�y��䜜��z;9�C7�����L���=I@�p&��8�	�	5��y�cL�P�[��ݻ�K,+�J9����l�w;
�Efc�M@I\�PG�#Xٷ�ǇUg]��za�-���۷�O!.q Xʘe�C�b�-�ҧԺ�W8^�6�������!�7���n7L�/�T׽�*�&�dg�ypHz��߇���ȃ��C��C�F�zm��:���R��7��g6��N��\�fyz{uo�ka��
�&z��^ ɌK��j�D��S=����L���ҊS.#��Gygݻk3vg��~С��:"-�n,��L5�T�o/�&�9`��m�� ���.�,����m+Xz��#r�����]�vQ��R+]A߿s�=��zۧ�zY�m�%Z_#���0]a�d2���۷Q�-�-1�^V�=xt
�g)��1MA��8���K�H���Jm	$*��GO�~��t�L��I(��s�Cd"�z{�v���h�9�YՑ�-g��˩N
˪B�K�B�Á(��#-kس�^ ��׷T��W���t>��ik�'�#[��2�4�Ǖ���&��[��z�۶����M��Z�D��N�3�oS���/x��QY��]��å�@���TŶ8r6��qu{�.�С;k��D��+�����Yۗ�x�4���.����"��7�0k;>�ٻrA�3�m���s�n�}��ݰ�,�T�h�셉�{>*f�}cA�8�%��l'"��ȥ��=.��!�C�aߋ8�[��mVe5��e7OSY��S��sa��*�A�['j5�Zϝ��3��l2۳�6ĦZ6��,$�L�X83M1^,��BB�f��kq���,�D`ڕ��Q��{G����4�O�
�4�D(��Щ��3I����m?�N9�5��S��qϸS�J�Ք7���;�4�7��@�T�'Lȣ�_�bjd-� -j��s�W`f�_�dN7�{�i�|6D"����6I�3λ{�YWZ<+��woP����c?.e|��B�1��m�j�M�'���똫.���վ���H,z7��f�/�=WM��5;��5g�� �}L��� ���l�a��sZ�������.S�C
�80M��
X�!iO�� ͐��	K8�
E)'9�w���_pX�M�	��np��T%����n'�!���2��o����᠍r��-p��d��$J4���λ��e�0.��Ht� j��2+�]�g�������e~�i/E��bR ��a�Z�;��O�#^֭�`u�6�ʳ,�vﭷx�p�Y��E�1�{ؖn�}�⾢�m��pU"g��P����[8J�D�n�g��R�
V6m4ۚ�
��h�KU�(���%�lki�^.��c�,բZr�T�V-*<��܇<�8�z�ԃ.�\��y��<����m�m�������AocX7`�gخ�8(��t��^������r8s֔9�2��f��+b�:6�%��.���I�2�Ve�[�P�QյA�7�f�4��k��:����)n��í�����ŭ�p�R��kҲ[�ҍ�;6�'�~�뿷vw�,h�/��+8kEۥlU���#f�<*U�k=�yv����D�/޾�3s��H�'�z�Ұ� �F$�ae�T9���/춲a������T����@RT*� ݡ�*Z���|(섫+}�r�Շ co��</U���&�Zo��VhL6�eo]��<;u=��n�����T�W�锼P����;Cbsw|>7�� &�l�B�ҫ[�P�y��U���ċҜ�R)�X����O{��D�Utܳ�4�D�f�ݸ#]��!�X {���i��dbluw�U�ZP�+(��K��%������E�zʠ�J�C�g�p��2ȦB>}�����޻�O���,c��~W���^��H��!B��'��y�3f�&�i��ݨGn]�k��΢��|Nz�v5l���命WZn���j�{#q��?�wf����{<�6p��� �K[�{5�ɝ�`�`�O]��!��f�� "�I]�>�v���hCi6ڗꍷI;{s��ѧ��lQ�������%M3}����;�
��=aެc�mO��5��V�_�Ozߎf��hSK��V#k�C��w0;�&2-���9�Q�.�O�/��Ym;�ϊ|�AdY����N��{��N��.�C,��M����&%�Iio"t���`�āy ��셝�L�6G0a������sc��`i�fD����S/{r�\KA8%�̢JbUҜ��۵��䏰�f�T����cp�(���]g�3K�Xr��w�o�#( ��Hn��f-���[�izw�"j��`Q�[��!��S�b�wN<�lY�swe�P�ʂVܟa�;c�=�K>�@�GP�B1#A��!���?[�0�Q�~ߞ���Ӻ�W�e�\Iu��z��3+��a��.�֞����82�,T76	�q�]����Y�O�Ws��W��|{�5�]�#��OXܜx�!}�"u3L�;�j��!�|E0�BP�b2$�f"W��m�3�]�ko0_K_;�x^z��F�Gj��K���^]�[��f�s��>�u3�y�.t��:l�X[��j{�V�uF�<�_Ȳ!���:���ą.[w����T��vgӚSi�w*J��W����f��X���4$�3Zs�[��b�k%u9RJr��g8o�]2��d��:���[�&T��Tھy�}.]V,m��~Ԯ��媆&>�|TAD�Q������(�͐�n�#;�d��7m���P���Fp�6gp��I��бIA=gˏ�*�wu3,Z�__{N�:����~��M��&8/W�x�D�{��7ȭ4��;�K\����"	���w���;���9++,U�pn0s���c��]�4i�PU/�,� ;h���Ƽ���
U;jވ��i0����̶���c�	=��є�!����>{+o�t.��7�5��M�#�ӟK�r�;_}���¬s?+Q������,�SD��q>s��X� >/z=���yp��γG���tj;����K�5��U����#M��9{��X|k�%y�\R�G�Rk�^�u�H4'_n�yOtM�B�v��$26ㆣ��@��=����n���n�	�+��V�U�4��ލc�D�7mw7�	�I�	M�l�Gؔ�.��>�`�z���gu�3,���J�������R4���*=.5<pT�#�nF�c�&zm����C��Zoc�)�4�&`��y��e����S���N<�3�8�	����]`]3bբ�i͌^�e^-Ά����Z3l�����|��F܀�"R5̞ɐY�yk=��z��B�������zS+[lT�K0-���z�r %o���VS@3�3y��I���<��TͰ��X�9v.í��m��2�8����]���tV�L��x�G�W1ryާ��=���5�׭vzQ�y�B՝��� ��L��A�҉=5�CB��ÙE*\�*�[=f$�,�aI��0�E�!��Y��n/z|�#=qg��5L��|k.>F>�'=�}�%�st���	�rN��i�7x�u�w��Jdm����ǳ��۫ny����iUw��x�I}�֐4*!�7�;�O�*h�u������_*�c��⫷d#҇�D�E6R8�Y�X�s۸R�wox1�X��P�f[#`�j�j�ݺ6/�F!C��7�4�q�H�ѧ��˹ү��c"k�7�4.E��Ap��
A��S%�,h\i�\��O���qB�&Wt'�ɬʽ|�Z�!ל�'�u�M 㸲d�Ǽ����qv"�UV�Yڰ��z�K~�HhCw���y�.:}Fʽ���v����<���G]">��u���t�5�؊��j�,�}��BM�w3���ܭ�(ڷ��?�ս�ʾ��΁z�+^�x������cx�-�K�f���;W��ҡ�;�ãh��x�賱Bxޮ��-V[��pk��K����X�[�^�8¹Ļ)u��JMŦK��gjz�*��ٓ��ٓ���o�j5�W�U��{�.�fP㎁��hEYL��*���YK:�yP�EmmZ���J0m�պ:Y�L,���z_n����;p�]��7x�l}��jv�5�
�Wu�d�7���)7*�e��DcEq}��n�^٨~m^��C}h���G��`Pm�v6��U�|�L��=ԙ�\6������ԳT˹:�lr��I��f�A����x���,�^�N.ǐ<�]ѩ+.�:���9�=w�֝�q⼛Re���,����+��8��=o�{z@w�$�3v���Q��o:9��+�B���WF��=W�z��W4��ۊ>�,�=�LZ/w:s�v0ӌV�{<�%eqm5�Oc(�h�鏆���J?��n<.#6�3G5��Eؚd�+VT�{F�=������Y��pt�����^,����'���&�\�s{ }��F��㙕+����%�B�Y�[K`�
�:l�\;l����vv=�C�S�(cV�=����)a�qe�ٔ%���W��N���5�	5�N�y[}��K�ĭ�4Hncv�U�v�c4�B��C�]0,19,��Ζ/�wT=v��=�Y�3��Q�c�y;{���s��e=���媃�UG[��Ƣڀ�����ۆ1
BY�CL�6�l�
.�Ι�pğ��������m>����7���0�S�����1��t�8�8L�K������[<����[(��dV�n����,7	0�;W�,,X$��]���ut`��tr�ո�s"mA��GWUl��ǒ���[\�z	�n8;q�`�sC��;�i<h�J��ӻ\q��M�-���#����Y����v�^���6^��9��cN.�Tٮ���7n�'n�9ۋC������ے�*�緉�21˄�4�B،��y�n�]��El�l-K�H���c38�H�Mls���7��ݤ�7��v�s��n�e$wN�~��~�ԏ��/:�փvB�dp�Ma�ĕa�Č���\ؖ��F���d�;j�Af�tۗ���JҜ`��)Cb�0)G*̜xXu��������t���H�[l��h�[<�5�%�:=�Z5�9�q�r�^�#zGj.]�nɈ@�}���͝ݵ��)�ǳ['�u�o�c�l��rڰH.ӡ��>�[Ӊ�1��!�b�<6�ϑ(�v��w)��k��J؜P���m]N0�B�(�c �И�Mh����:�\���9�w`�i��tih]��os�g�1Y��������f�����1�-ֈi��J��-�(� /T�tl6�q�=��_|�s��y<��pe��pB�K��`˻��U[)���Y:*�����}�g��mA�nʼ5(t%�sc�@�6��z��\G�ڵ�T�cj�K�kht�k���Wi��W�5�7B[���Wgb����l���Rav�c�5�[�H�-�eN�C��@�Hm�5�.��wV�����"�%�h��*CL]Rf0���ZV$l�
�,Dx�ؗ&���vq��[�^�3����e���R�2b�vs��Ⲓ���oKp-�XJnΞyB�v�����MT\<ns���rF�ʎ�T��R�0�:[c��)&T�fJ�Ni�q��P�m���H��f���VΧ��Woj�&�������R^8���F�zw��� ���n���#���@�n���e0N��^#�Eg�A�=�\,���p��4X���Q��i�������;+غ�7fM8^�<q� �b�ˈ�mf[=��]`\�	���9�u��*�� }�7�Cv����ga��Qs,6���]U����+ϝ܃ۭW��]nxRiۢ4ݰ���c�k�:�I�l�����Q:������]lL6	v���֓9_�̆�u8�^o���+��N۞n�������N�w���]��v��H�i�Lg�Ɗ���!�v0Ύ;&�+:fR�����:3�<;U�t�S�Wd^�a`��d5�X���x���J��Eoa�:���r���wv6��Rd��iN:eo�vAx���h"��Q�P��Ok�;a�#E]�� �J��~�k��|��V��r�E�뽾%0�&�mڗQs��ה��m�	�zܶ�y>��e�/|%x�{6ř��1�D���o/;�;�w~g�%���7�P4ۂ2Á'%͆5y�a<�6j�s�,�
��x@��Vh>����������lEN���k[\Y��J�'��Ba��<�����m�Dֺ!���m،��m���X�Q��&��hf�&K��lOnQn�N���1���t��B�������@f�������5D�m�hK�m0��[�.��c��J�T��X{Y�R�T�m�G��,�������K�oN�i��t3n�1!*͘K�&�ץ�hj�j)]�OM��z�5@ԃ�Ɋ����.���R�y����=�n�-ef
�Uv5r�1�nl���MK]u�n��r�y�~u	�kl��d0��@�Ȓd��iF�Y�HȀ{�Dz�l��y�>o�6D3O�(R��S��UQ��)�o�ѭ?hX���-�t��E�y��[Ć'7�v����[�d����^@�y��2��>���x}��Π��޴��l�a��$��ӿ����u�FRw�z�#��(�y��!m�5;�̮LU8iVc�)ա{Q;��J��E��䡦>+�2a�E��_^ߟs��z�_o����5�%��Mӓs�j݊��5�1���v�uǶ4��� ,��u�K��������� �����u �l�]��"���j�!D5��k�"tH�Ɔr�D#7�r�Dh,��_QX�n�6uQ���|u>k�m���%70���M�%��Y�zt�)�S��*�x��L]�ޞ)Ӝy�p�OA���8�o���jFa�EÒE<a^1cΜ�0)i�,ӛ�ew�Vr�UK�Kz�wJ�6�S�
wҘ����U�1R�Z#��Ԝs��%n17n�D�ś2
�39Qg�ࠨ���A(��Q�xJJ�u����4�z�y:w��kO�GM�Vf�E��	�����q��3޽�7�w���|9p�
6��5�s�GWr׫�k����UXtYY�=g �xn�k�63��/S�Sm� ]Eĝi��j\p֛�u,�ƻ��ˮ5e׳C��:|���Ր''��9ƹ5n��xaݱ��^��Ԏ�����i>���=f�K>�N��"s������4����᜜6�8�m�/&�XZ�������t��X<���������EQD���وp����e��9�HM>��n�z뗫s%�3�/�aA3	Q�	97f]�AJZ����3�h�]���0��>J�{�{�xnQ%�'Cև�v+|g��2��Ǖ{X��i�5���:)�e-����]��?c���^�~��N�������3�<"wg0:H5���4s�F��h�}ܭ�/�5J��Ө0�H%����~{ww��N�����ǭ����s7��j��7�����^��[����������6��x��7wm����XY��fq�/�^�pJ��5t�*�˵���P�� bqʲ2��zLrΥ1w-fb��=1�VF糣�98�m�;�{��Vn߷GgG�?S&'J}�[y緌�F��]7�'z�H�̓�b���?,�u�ݩy�8WwӾ�c�`��4O��4�nx�vW�����������)%���6,�Q���T�~�Hzrb=��y1�/h�.��*������yU�ݢߤy�r�(��������ll��>�S툸�ٔ�W�>Y2
]O'/���$�/���6��ue�FyKEQr�y�h@e��(ڝӇ]d��_=<�$�vO��c�>G!_c7l1SU w����}�{�|?i�
S�E9�k�9��K��Y2�*��T��3�~T��<�b�}gz�`,�~=�Yo��԰�A��f��}������]�:|��l�D+�
e��ͱ�ޱp]��0��V֍ݲ�������䀼oH�{��2�n0�` �Jk&�YL��X�i����Y�Rg��t����M����V��;'���
�8aݺ�l�r\�V84����d�ٸ����[^��WF��\q�l��8��.�����5+3�֎^�'���.ҭ̘͇��h�~�;����`>�ǭ���ue��.;�4H������*�ˁ��t@Xª�T�Ut�����W9I\�+k��H:	ʸntIV6bl��t(2�6�g�J�nYV�0�#���(
��ʲ�M��VUȐ�6K4��k�pR�:���t��+�pڬ� �&�ڞ��ƫl�4���mܮ�6cC<�6c-[3Z��ms��ݳ��1�쇷"F�����\��a�Kn-�l����/]nwQ����v:0��[�Xe]��[��:��`e�Y���3*������-�����~з�S��&$W:VyX�˜}v7r�I�je��]H nj�TL����w��~ʂZ�)�q�N{�R�Vli����?W�R�J�><���z�z4:D�C�l�F5�U����7����:�
	!m#	b@[>�2�{E�����^J�����B����;�[���΍H���׀�I-{ �4�lQN��4kw+p��s�1]=�m/���M�k���n�)�؝�c�����$�E�z3|M:m�0��>i����.�U��/Uf��iyCԫ�8����k1�Ŋiw�5�ð�?[ ��3��{1Ԉ2e�������;�G��؁C8�,�Yt���Loŧ\�\����;aG���	�&a刵�w���#��k��U�� j�:�K+�9�_���y�(;��K,�^X��ԑQ˕3<y~��,]�x�$�aH�N2�p]Uĩ�p�t��:�X�ep�9/��C�0�����&���5���Y��Q����W:f��g�6#\2���*������������3&��--ŋ��{����6��?[?K��!y�Ɲ!�Hk��+�vŊ�^��s!b<!�縵�T��,
����:�]��^��a�_z���z�v�l�
ɧ���_7Hsa'��ՎW��v^1�$I���&5#���*p�/"7l+�k��B�p$�ݛu�0K���;�����*C�Z�VNz��^=%F�JWHu �i�R)�ӥ���:�����^��EEmop�x}����1�]C9���%X̵􋼌6,���r�-�K��^�ˬ{��B�j2�釛��M��s��u�p�=V��X+�[���Qf�3D�թ�N�]ƍ%=)�޸���,~�eU ��a��OD����[v}��Ԃ=�Hwޮ%�&nwQ�,�Kɓ�8���Y��M�E�q�k��x���0�Ǩk4��'���fR��͏���o�6v4f3��6j�,mgw�M�RTj�y�9lG�7��n6�zx�{b��x�S�^�YWORe���D=�w�qC%�t�����'p�Su�S�VCr��n�⾚w����p�T��ul��l+h�+^V��z,e�D@�n���.���|r�Si�E�	��m��bc��{g+�-	hJ�i�`�$S�N�X�����s�Q�#�M��x��Hv�9��I�c_q������X�Q!d@d�0��Ufs�/7(A�=�vn�B��|09�l ����}�[�*�8��^Z�\^]}����E�6�-�w奖��XE�7�+.�a`���fJ�Cr�9n��Eڰ6:Nv4k�I��v]m˭�?n}{�׬�[�~���h��yji1��(��)��Z�(�~~�Vŗռ3X���{���+���ⵥ���wU�5T��s7V�Q�R�f�;?i}�ٔ�����%(�\5�e��I��{��ds�vŔ����,�M�P��D�M�Ua�xP��3R﹮Y�KN�{nJ�Vb)����l�ݺ�Q^��M��5( @��.䆔������ �M2�M��7٬��3uؽ�7b�.�Ǫ�_W!�V�U8����YC���C�&'1��lY���Is��Lɗ�����,X8��Ӣ��چ�=��ڽ:�Ը�\g�҆�&d�U�{���8����٢�������M�����f>~����B9Vn� �a���J,��Tk=w��8��L�{n��<1�t;�	J�T�!�zU��r��$_eĹ�zw��Ϋ=QG1������G�1�
�)*���ͷ����.*�3�+m�L!��-j��������@_q�ɔd&
�]����6��t��z��W������{��^�F��Rl�
$��$�aE�E�͵P@�M4y^	Wq��i�e���(�J����T�}=��9Va��4vPu���\�GQ:x�*H��T��Em��ݞ�֋���������Ӱ�tA��i�Ue����̭��z�dV@�6��d�]4$S6�R�K�u���w9s�c���B�?(J�+��J�!���]�;x�s�3��Z��> =�Uv5��}��#d�#�J8E�|Ş׻�a^*�M�LO�?�3��4׋�@hyT�)�����cs;�jݴ���1�a�:}ӡ}��2~�Z]x��߼�/t��q��2������e3P�B�����4�ң��K��N\� ��s!�jnX��<R+:}x	Ŋ�:�"��][aA�:mM����=Z���b�J��+�o'��Ɛk�m�-�-���ψ��t-�Q���r�v�d��~�׏��M�ix�v���ŋ+D�m�.��6RFh&���v���,Ô���5Η�R[��vJä�]o@7TvM�S��J�V�S�����擧�����s���g��`{9D��6 9�3ܶ��Ѹ����0B9�i���8S]+Ŧ�ܓZ2���q�d;9�[�n(��6�cv����>�ܓ��?��}��:�̃�;lQe�+�39�3�sϕ����U��$��d����/���c1D�� [(�`�������\r�_{�B��F���,UC��4gh(8�:'a��{0����(,�-�E���c޹�>'��������N>��.��=̉w�Y\f��N.컻c���8��g��c=���e4�kOceƂ�q1ï��	�!RL2ZL������8o��A��>�*�Q�f������i(�{�e�I\�)UʻO�G�{oe����h���SR-%xyv��x8��<{'[��yW�鿒C2P�<u~�m��=��}J��Si�UX�ߣ}y�3����'b�"6#�s��ƕP��t���d�R�	�XH8rм�R�]��������ˌ8x.�wl�����j�結�j��z��G���t6�eS����u���[ta��H/xs�R1ā�Jc�]�њ�c�z�v�Eޗ�K�K+�X�Բ�G��ײzd��c����G�wayMV
�<�I����c6�nA{��:�X��3|,����W�_~�w�÷�l�Dx{'Gg=�>&�>}4��1���o3��wO�:�ۋ�u��g�.~�q�W�/	q뷓;_��e>���|��jp�$��2_�����l��^g�Krw1��D��JI�-��'7���J�׼��'��]s�ͼ���n١�����:�B
����+/k $��}�S8Dw.��9��A�IS	��x�p�L��1������k܆!�̵)y"|�����Pc��O�)�|�3/
��n���)m���"&��A�D�f�r�SBk����]E�c+%Z��p�.��ƺ4b�Y��-���z"�����E4����U��.ٶ�/|���k��w���v)�����m��
bH�%(���ׄ߭`>�/�O_�K�/���=���\���38B���y:�-�~{�g��{y����[r^�m��8�RE��D�c#�S�����>{*r�bb)�rƲ�u�N�ޖo�!Қ���.����Gj߯C�M��h�6JY^y'�����8���et�ٙ�[��e�/�Ÿz��h^����Ruu�������pJM=c��glWX���w`rޗ�&��1�ɡ|}\���Ice�r��nAa'����r,���wrՖ�N,/���d �&��坂Ƅ ��-�G٢�ԞMw)V�m��N��p�
�U��nnZ�xBÉ�X�d��Nw�# =�.\ݽ��̖�F=&8�꣖��4�����W*�ʙݼX��j����X*q�e�j�,e�&��4�1����${ֳ˾'�SJ�Y5�k1�[�u����d��q�٪L�sV'y��uY��
}�#h��C��0j�C7�-fǕeޛ��G�=�e_W��N_ Ug:��˫��%�pݼ͝!��)Q�YC�y��P�h���^q�+)�Lwӎ�z�V��̀��x2d]ʹ6h�i�vV�X9u�5w�uՉ���6+�*�Y�4v��Jt&eeq� �U�%�Rޫ�ݮ��
���4G�+b�*�(�Ŏ@]�5�w|ص���s�["��ۅ����k�xg�u�i��q���]#�N�q�����W���/�����BB�[��q͐=�9�˽p!܂���}D^�Qe���|�Cݕ�F y�T��>��*L/%>U۰�w��錼U9��Yd�h��w%�n��QD_SU�,5��J��{���)^�]F�.ݵ����DE؍�>��i��p̮�6<�v�#q�۵:��=Vӷ�^+ˠ��������޸M�˼���.��M�BK�s]4�n�w޾�W4�I��7��ʲ�>�y���(o�&;)�}\S�7�<��))JBI#�:{�ȼ�w���'Mޒ8��r���Uf��Vi}&�%��q�}ns�r;ĠV\���R��qj��9j̔�6أ�a���u���=u�j(F]i����̭�<y0FZƺ����{�:�u%����4w��Jбܢ�gT\�u�]�}-v=^5��#���(#l���M��{��D1�[��0�����:�H��z�z��c����I�K����m���}f�N+ n��-�co3�U��ut^G;׈�X%0�M�	���t)�S3y
���aܬ�s��Pb�¯���F7G=�;��)�ސ���2� g��R'�)٬륍2~1&�
@�Q}=��Ȟr�`rz/�Wuf�`�u���A�~�7K�)�+�8��gYx�%I���Ff���Y�V�r��7�u#���x��IU���P�&1��t������w���7@TChW��74�ڙ������[���圽n�l���&�i��-���6�3E�����D"�s����߳����*a�_�P]#x\��1��>�㷞eRp(�%�Q�)�;�N���e�hs� �9QuB�A�	v��Ky�9�	��;.�L�[rm������i0�V�IRT����uk�t��1��~�5L�\��?Oo^��pA��(�Ӑ5���/�UX�h��_�$��Ta1#	�""<��YC1�m�&xx�r��n����g7��o��6�a�I�k����/���<wOKW�.Ϥa�бTq c0�	�]���j�9����K���f�bЭǷ<�@=�i�m���/NR��J�N�Ҕ�w�_����ĺ�e5"����2r����+������c�)k��g�+�V�Q4_�T�'���UՖ���x̿��.�R��O������ ����i�J�m��e(^�np�}5%�4���|�w�n�?a�)�0��G��I<��o�41��C8}�o/�ͯS��yJu�ߣ�>��mi�O�[�5�,wd�õc���r�*��
�b�5҉K��h��0�(����lT=fB�s�[����#�ВU��"�1�����[�8�z��v��BU��J�JÌ��H�\��n�h�i��R��ӋS��Ļ���7��z�mʉT�</7;�dy��l�Cvr��C��l.����X���=W96Ѳ���ܒ���4y���2��k��[/�q�s�����q�2���0כbcK�hs3V0B���2v���7���A���*��cz�^���k:�l;Cv�S�*�]�i����U����6�ǡ�T�UJ�0M]F�j��}����ܻ��5V-�HHw����%:�w'��z�����{��[�/�Jv��6�;����<M�
�PFuz�y_�_r_ߓ�m>��~[�(rQ�c�	*������Vƫ�Y*���>g��z�ֶ��%?�$[f�%1מe[�g�=��7A����c��z�%W7ް�Ir�nJ��U$Gt�>�:t���ҷ������m��{���}S�wGTN�^3j�ny�g�=����������$�����N����*g�;�Ͼ���^�Q��;�R^�H��)Bb:�y%��dR�J�G��r�������6�����y�0�����������d��\6�%�/��H�F�Χ�U�n�i�ɶ�f�u����F���щ-}r�q�J��n��y����}�x����~��{'	��M3�`N�z�C����Z�v湣��.�1y]�3��JS���1!�DT��T�nc���M��o���PY�	��+�/;9���nA�{:�z#Cy��}��hf�+�|�1�m;�s.��w�q	�[-艂k�;ي�{�|��|�m�����x���.���Ob�֮���b��v�{:�>�{����*"�.N����(�WqTf$�lӄ\����A�3z`�,�������6�E�9m�6��_d~�uk��r�M��ۺ���`��K��&{�~L=��ֳ;�H`!T�Z�v�B���*�׽��aQ�s��U�&�&�.=�47�݃ϯz�����^�wm���m`�Gc��W)S��C��)-�2�7hr>ü�fY#R�\տ4���P�z��&z5+�e�K\�T�x��7|m�������]�ڋ��c3̷c��pJW6vM��ɲl��e,��A.��Aw_S�
EV�3��ط>˭�s��;�y�e�=ÖP�7ez��N|��ܡs�6���v�mM6y��
��6�!���@�{A��8ݎ�Ⱦ��9N��~�'�L�$�+�T�S�|��.��vx0|�{7}>�3/������L��4Kg}�d.�\��^�K}{�"��dtۻ�%�8{����&*�p#:�s	fi���-�ɩa�˘���yYز�+��v=4�Pt��{d/Egp��(��pJ<@�^K�5^;·9�v��=ݯ��=��&U��B�p6�J$�V%��Y�$jZ9�JW@9}�מkxǡ�vG\��tsn�\ǳ�9�k�*֞�wQ��Ӓ�k��h��;��q��FBR5$�{��Bƫ�p܈��]�/��˞;͝�.LR����`��Y�X珹��&�+z'�t��~��^�tS�Z��Zc/n��S����7Tn��HAhM�̛Cm�D�&	R���Qx~N����{������{��(��
[���Y�j�G����{�P�L�����b�H߽��%F�ICIų�j���;K��h5��U>��`���U���l��b)z�o��_���]�/����]�}QW��aq��p�"Ir��m�,���)�}W�b�o�悈:!�D%.��׃^̕���P����i-^��c0�!�$�ż�Gr�ğ{2���LםJ���	ՈH�_�{��L}��y�[�̶ϯ���}�X;;Έ&��+�����W��Q��&�*% nL"�jΪ1���zۡW���G�[�.Bhe㤷�ÚU��Ǽ+�:6ۜ���a��E�	 :�HT�ە�_�;ǽ�_@g���u-[]G,6�$�����U�~�W�֗�VH��#U��ΓW��߳�v�W�A�N�y�Ŕ+�"-�kvLD�a�G18��55.40��a��ap�S��[�*��tN[�\�e�m�U��ؖ�L�&�+<��O<2��4T�c�e��*�N`c��aIMC`� #m��[�y�83W�	���꽍Z]�\����-{Kz-��S�m�*�yU���yDU��#ًyX	j����ʌpc;��%�~�q�B�$��M��X��.p�9���u��}�Vl���SE�abu�b�j{��`��b�����l�K����P�N{ڲ��n�5�z��${���#��L�y�9��<���F�4[����J9 �A$2�y����5���CZ��u�s$��y�p����kk4ש�H�C_Ya
*��wL����86+�"��k����T����q�{`��HW"�<�+��O�)G����'b�����z�WV"�䔻Rl�c�����.��g��!y�o��#[��9Tĭ�gE�g�v=�glx��lA�s�W�N;yఎ��v ��q�뱞�-'�R�ڞ����nyo�]�%��7i�4D]�b���#uU����n
�L�����-���;*�G4�n�Br��6���-����ٗnWi��	;;AƮ��ӀL�����4Ҽ\Yl8d�e�e�-�s�=�̃6y�T��fٵx1���m��f�_ 힌nqv:��G��O	,��UB�!�Ŗn(��r�%�~�KO�=�{�h�A���(fVn����	,5�U��i��<Tͅ�Y��\�s)����g����`L��� �&m�!ñJ�Q:�^��j>�w��_����=E^n�]���z�f�u�9V;��hӤ���w��U��U4p7���iQ?n�~��=�tK�X���\����(���ٕ�]�L���H�/�����,d����J0v�r�})a�D�Z��~�lu��P��N�� ��c�+V���c��<.n�/ǭ|=7�����.]z��"(�E�Suv�ӯ�N4�7�
��0�k4� �м>�w$�^��/j��y�P�{���w0[j���c�2�k{��L��\����mӎ]��np���N��^1��o�,��`���65a �b��~�d;i��^{mfI�7��v{���_�{VR�C�J����0�]q7��xt�����#Bd�LI�
M���*����g��o��*Z:P�F��0��9*�ְ�d���.>���Nf�v�O_ay�D�;-�rP�#�Q*�].H��2����us��fP6�o�[�:�%s33M�|:d�����
=.�{��.�y[��OO�{�z�L4E�U�O{����ę���I!�!��0bS���v�J���N�����1�_+��ǅ2�{v6,^(��!n2
j ��9x���6R��)�x��r��V��þ8�'��q�W�~���w�n�#��l�w�sY��"0�L�YMi��/���q���/v��v�R��e��[gQ��W�]�����c��z�-�j���nGD&��a��z�n	,��Jq�h3��"fe����e�Ux���,��i"Sd�D��i�~����s�ŗ��6L�N�ٯG�s�swڵ����r�YU7s~)$Dٗ��[�SvՊ=�a�Ɂ6[�4�9w��7�C�"c���F�Зo�և-z�P�֙�0��3<��/H�NXQu���'	�kp�vq�ȴ.�tiȊKRH�u�*-�yn�a\<�m���1�u�ž�?;���z��oh�{*�[î�H��i.+����o��{���쫽��W7��<�ѝ��iٝ��+W�w%��=�.�+��CPV�P �)�@4A-&�Cד1�;�/�Ѭ�7�g˗ݴn�LҰ>SC٘���N���j��A�ˊ��^�������>Z}�Z]�;��ʊ*�����ni}ݞ�TU���OX�̹�J�9��W����n:L�Hc��Yjyִ�݀o�.��rAW����&��H��sA�H�Q�g�%�ez7�]���mn���ei��e*e���N�;H�Ƿ���:�c뜝ժ}��y$�3{+���*�%��
��4�����p���o�F���
���d�g����jn.��=~�Xb飁�.׽u�G����ClOb��-����4R�ǮQ
���璊���l�~�������x{ď4�iʑ��iǣH�z�0?^$�ٹ�ʼ��9��NwQ+e��+���!�4�?>��g{Bَ�����iDC��!j@��B	vצ�3-� ����m?<cC��w��s�m����.i���F���w21�J�c�Q^1�2�c[�o"<)�f�mdT�p�C��s1^�/�T�(N�C� �Jo1m�gK��������26�p�̙����׼�w-l��&�*�&�)�d��qgE{�w�o�Q�w}��czi�WkY�ׯix��1'Y�)-��^��
���ˬ�"'ƓzGa����,�4nV�摰��p����0��cWZR��Jk)d C�H�a��8ɭ|a��r���+��n��� ;um��|�[pOA����8O6��cݐ`2���_~�˨�Z��� ��:�7�\�[R��)Q�)���%�-�swB��y�ۙ���%~�F��E�~#r�8{�y���	�@�IAH�[�}����'����%(��&��ͤZJ{*X��-�T���>�6k�u���-a��KR��wvv�{�e�<>�B���p���Ֆ�!\�k��> ��1m�Ь��0?<�t���vl�RAv;�[$�:�H��Z>�"t:�w�}36b�9�m(��i�N\uv���S���՛|Fs��}Y�Zef��1��j�a.�X�-C�$q�o
��qh�M�+z��Ù�N��Yw�i�P-u�����R��3�j|�'[�wI�k�3ڮ/%]��
5����*ģ
�ƌ�eٲD7�ː��5��Jē��'�,^�>���˱;�$�h!���8���Ua�;GWXx�,�N�Nv�F����s�5�H����[o6>��J8p��{���V�!E��^SOwin�Z�l%ݨ�O���6R�6�M����mp\��◔�-��坠\:�._Iq�����]�{xGћH��ܷ*7��x���e�""k��3Z�u�4Vcs�+/wZ|.��e���f�%�Ⱥ��N��3N<=!s3�b̓i4��JP�����i�M��t?ޛ�j�3�9�w:1�0)��K�[�I�XR:yцɴ�����Q�w��C�D>��S�1���n��ʍ@�sŝ�Ko���ߺw&�u؈ӏ^��i闽��Q��t-�gЙzp�C{%�\oU�ۏ/�	4���j���M8C7���zpfq/k�U�;��ui;ݔ-��X�-��ѷL۽|ݶ+�s��;նM=*��x��W2�0��*�p-��R�jև�yr�����{���S j(oh�u`�4����d�^ع��e�c��aa}}*�����rV���]�m��XWc��ն@�S�d�Vx��h+��u�i��R|s� ����O���y$�*���5C�g�p�W1�.�*��ik]�I|�����w���p��»e�k�̓�b���Z�X��K�b��`��%���5��n:h���&Ea����7b4�-V7F*��WH�;FĆ�Q��(�	�-�c`�2CM���w���b�r���˸���r�ø����Vf���8�>v3˭ �#��܆���gg���=�C���ў]�c�;m��p�xzN��8m��Q�G-v��N. 	��h͡+<�d��e��qF7:iw�b2M���Uu�@�k�c�Z�1��f�GJ#4���Sgc���,�no\�\©�HGI��޶nw'��κ��}�C�>۲T�NۅCm�k���ºJJ�k+��s�kLRh�]�g���
�OnM�GK���˝ŋ�2�X�fk	iIc�imLq��ak\�f_\�ő��X����)5���)2�ڵ��]I���a��t�[c�='��v �njEۚ��6��	cc+Gm�b�Zˉx䑹zg��	F|�8�{{��Wd8�u�edfт���Ma�G�mZ㭓�����a��:�.����4k��F`n.���19Y4g�B��+Z�5�̹��-�q���#���&�Զ�J�ٌ`��;i���d�Dx��F���x��M�;��*�s��/��͚W���6�ɍ����h�F)�/%���XJ�W���%R�1'+0�۵���w(��^�p���L�gc<�����%�шG���f�Xt�)k�=qv��4���+�.ɮ��n�(�\��:�[�����\tT�7[�tq������n��;m�ec�O���n�Ѽ�v��(dz���l���y�N:�y��nz�6�)��Ǘu+��k��]�+R豅+s��i��fبxێ��q��q���f#@4ՊglLL���h�Q#��.z��O.��ڭ�{1��ǲ�w+"��ָñ�$x�j�".��8��U����1V�aƋk�k�t�ˋ��75��[� ��\$�:�p�	�7&����.)1c�f��KsQ3ʁ� �ѕ��Y�a�������d لC�ŰPWYv%�P�.Z�6.spp;�۷��⎻��Խ���q�nb�zj��΁x�����%���tA��TkL8KR5Z:�Ōb;],s��\�����k406gh�&H�^3Yt�� �u<Xb��c�xG�F���*��f\�a��
Q���爱�u<���ۮ���o�bf����x��m��æf�j-�q�͗+���>���buҺ�#+�vp*կ7]�2؄�~���"�\:=�ݮ�y�Y��r �)S��h ��+���B�wgЯn���3�4ROe�Xs��Fg+��ނ+��ՙZ�7���Kv���}��&�L �fHs�s���z{0�'~�������6��%u�FP�z�/m7<����K�� ���}F�i�(5H��]�W�@�U���i챻�痊��~/x���{8�a'�"��xf��~���̱[���&�A��@4�^g��.����(����E����z+ә�}��J�Lm�7�g�<�}2�S�Ƀ��÷x���D�������"(�F�vuvܸ��
�n֬<�OA�]��KƓ�"`�`��mrX�G+`�0��3�=��탸��8����^��"z����_���bV\�VQ���'I��`�Jd׳��a���O��M]�P��{I��R�Ͳh�,ʃ����V�#i�vR9�1�����w����NFpC7�tw�+�λՋ�G]��V���!/�g��;�t��v��1n���J�2V�=>�T�&�V�f�/C�wْ;'8��Qnh���8�(9��Mڛ��c,ǝ�|��N6Aͺ��b��q_r�Jϊ�ӥ�>�Wj�>[YV<GY�M2��
l^m�'S�ۗ��<%����u�>�B����w��*&9������awu�+,�/�w�˞Ƿ�\�G�o4΍�80=O}��2�	8Yr����Z���/z���"����F+}|SCϪ5{�32.�\yj�J�_N���-e�ϑ7;�|8�.���%�a��*m�(d��3�i��e���9�����
&%�i��5·�z����Գj&��j�),�ц//Y�X�jg�6��9R��o�w%Ժa���>߮��gX+��Rν�~덝]�;�'�G�P �����m:����/�$����Pb�P��2�����V��������3��B�T�a�)
-<:�}
���q���$��^��r/J�� ��b�
oZ�/qAu��5����{�e.�r��.%�Z��`�9�]攒�a��#I�\�*u�wd�1'qu�ћ:3����M�/�/	���F��	�NK/)׽b�tOm]Ũ�f�0�����'yٙ��I'�ә�[^	g��lE_s����c̑d��|g|MM2)Sa7Wa��\{����Lb�q��Tt��obye�xzy�p�# Ш��3E��{ub��EPo#��:����������`:j����(���ۇ�ӝʽ��Yn�1B�Bl띕��*�,k���lc����I�^����V���J���m{���n���o�9*Yk����%��@4�m�H�߳�q���bT�������s��[u� >@��v�X�Gx֍Է]��p}�ܕ�N&��&(&���[9�a����S0���HW�J�tLF���ٵ��-���.G|�˝���L-�pRT��M;�o|�jd�CFy�F�==te���wg^���F���,���+2w�d������zlG���S+wuV�yx�ػ\{���[��[��+�]Ռ� ڼ	<(�l�F�� ��o��R�>�s����ER
(��
�<f��kb㙞�������1X4��k5%�\w�	$��֌�f����1X)��#��W{�L�Ic,VH��(;sS�yۭ)�8L&����P]����Ű�];��P�j��7WV��s�w�nѺ)C����%��nw,�e�'�{�w׌б�Gl�}�\[��I���v������W6
��S$����e�&*w��R�;Όݤ�3ә�z�-z*^��Cq��w�U��������Ŕꖮ���H�b�0���g0�
j�8����-��L��W3�ܡ�S�,�خS���!��@J��b�T�U.W==D�m�h���X�	5	��݈�lu��{c���=�.k�'z:VP~4�)Z�ůd;�ye���p��BJ��ے{�PY-���CLoC�z���yմ��zT�+�f*�҅Fvm�8/2�K��У�}k�zm�8,��;���D2�
ɽt�����1�Hky�wuCkV��*����j��U<��|�.��ӝ<�u��)6Љ6��##��%�^�������Yl�N��ٺC#�xܻ`:x�eN�0u�V@�7S��xNԕ��/����BR(j�	cLr��fΪ�9i6e���8\�2��shI�RZV��X��ʙ*�ӳ�L�DXs�w/0�%�mȉl�n0�-��ʪg�qn���ۏpg�|�0�M66�΂40�X�11	�:�
�X�kb�cv�.��0�C7h���IH+K�R�4q���b�Ȼj�(��!9Q)IB��(�[�eM~�?\E�����U�s����XR�����ˎJ(׶4�(̆Z^þ���F��_�՜
Fi�D��\��ث�VP�U��=ɟ�h CY�~�Y�~���$�G-�_�J[٢��J:m���{udO��s!����0Zr=�D3�]�C��f�:@#0��c��}^�����^�0I��`��&]��V'�⃓����4�mY�������v7obu�����ٗ��M;�}���u�瓗|����:��t]0���@�r-x3�� �<^����#93{膛��M;�3��0�"��K�']�V�l��'�����;z������k=���0��Q�`�Rm��Yn�f8\5(C�]�յ�:�|���"��]��]�a��T�巶i5�1�/��5�g�[Pd:��_gvU�3�שw�d��~1�B �%H�	뗁`��]o.��{1�O-u�2�(�+�n�q�U�$��Y��vv�Vu�X�*�[�Z�#T�z���r�J4�m̨��J���R�}0��{�s_�GG�p�8NXk��{����}�z3:a�;�k/������礝i�b��^'>�K�9Z�ߞ)v�����*
���9���$����eUľ����><ﺮ��gr�����P��]6 ;Ǯ���}�y7��ٙ�8['7����U�uwyL�Y�{�I�0�dA"��S��g7,vd�e�N�,z]�z�]���Z��ՏJ��Ы�a`{�~�F���:���,�J�!�V���h��sR)���}gr�$�ѻ-ƓM9v�3	Q��6�N��ͻ�G	]�}��s�CFAg��m�
o_y�
�R*ޘ��;��..��n/������
e�k�f�.��)B�i=⯵�h�׫��0cK��]�f%�=4xj�a�9+̺�I�cq*�sW���Xn�i�I*e��m���ǱDN���Zy�\t�ߖ�;�E�n8tG�}�*MNd�&��z��"��u�n\�.���Ku��h�j�}�Z
���|nVz�U"Ք�!��hg0��=>�.{ts1�}���b@,@ӯ^6s�u]^�B
��/`�	ܮ3��(%�6��e��e{�=ϗ�5��\ꝇLpn�uˉe:e�Yt�M��K�^�\�n�����/v���O|�M�Pߗ�=}lOTMuOǳu�,�է���yVe.��k.Ή��<6��҉Ye��՞{�h���Y-St�����O^J{��T����t߼�������÷e7�w���3����b��:˫����l��6LZ�4�`����<����b�Z4Ǥ��a���x˱�47n��ט)ngwW���q��6�
i�r�dF�8sR�ٙ�|B�\j�oF}-PR׽M`̨��ג(�,��{1t�o�{Ĝ7F7d�"M�-z&�&\��J�QM��.ދ����|y���y�r ]�y�����笮�J18{D�-� ڕ.�S��f�����Y�{� �lV��i�R���U����� �S�Vd�U߽;���=�+����,7�8�l8\�t�Z�S�}���i�^���tɘߪD>�vi���G�P��zCo�Y��:Q�у*�R�e3f���'nu`�l��t�r�V��K�ѩ�^�v����i&��p�=ӣwV=Ͳ�ݝ�iY�<���N�o�b�\8ͩ�Q�����n��g�߽��H��,r۹����Z�=��{0z����G�%(T*��OZ�s)P�o�	|<�%̽p1'��~�s0Z��/6�mnc�c�&<f���k��[��s,��կ�]	�7��ξ�<�����9��'s�q���ZV8wG�I[LF��LD�>�8:D�y����Iq�gl�iz:���I�n��R�7��ͥ�b�F�/��g�O]�P0�m�:�CW�.yr�*�qc��'C��쨓P�"�d��~���w��3�������:��V��;��F��g^R�%���va7M!�u�.d�z{��t.�c��}��'y$[�C� jP��P������ݯ�mz��8���,ю+�#I��D�۳�-���-�:Rh�qJK`��h�,oe���v�����pB)^�Ř�`�ͳ�]jV��.��9]�C1��;rҫ����`G	V̲��U���3�n�����l�qu��␴nFzܬDݖ��lb$�qn[a�8ڵ�UX�De,H�4+66cY�J�V;2�D�X��"����`q�%5���
z���x���;lb���71��,��۝�;3�{{sp��6�E%���˿~�v���u���CE����G/b~�$�u���B�	N�á�^]E�ͳ��%���\�6��,6�m11+.�{�_�b�;�J��l5��+��ݫ����B���y�{�m�oPF�M��&��"�wO+BRӄ��Hwsg��1��� "���u�ue���r�r��&]*v�G�{��T2�z*���i���@��r,�FHOP�Zpn�&"�8Z}�*[���P�^�	y{|}r��[��La�:�dЕ1�7/''\��m,�b�6�0�	!��w������T)��-��gm��"W�[�U�(���y�ֹ�˴ƍ*۳՞{IV�8�@�	t+�Y붶�3�º��.��f�s�6P!�mkR�vP��dnV{��I�"_�·��ʏx2rT�⡮��v_�F<n�ZSb
���P���#��e���FA��7����bf����=ٽp��� �K�	�eY�݃qn�q0���:����9��5�xuݫ%��7a�����;aT��hvg>���W��a9��a�$�A��;O����]f=�.��W��sX8��I;źj�gSn;�(��(�mR�[�}�md�z�z�4t�wE(�.x,�^:*���u����a���|��ZE����l��FYSAS�^$��jY�g��|6S칧KOk�7Z������ݣ܄A;�lB^u����t��%޶����S�~�V=*韛N�I��A昬ږ��{^�7������v�
:�'ݽu|P_C�ܨ d� ��
W���}<q�åo�&m�w�]��b�'\x���\q���[�&��.gE �쫉�Æ�-WfД�~���H��{R����YB���{|;{i�����]Ը�$�ܭv^pY�pש�⌾_��@�IG �Kn>`Í�\������f����u�cIv`<u��[���چ����N��8�Y�]���8w��X7mE��ؚ[�܂��Lu�v;�����7r�w�S�P�Ϋ�ƒm����}����Սv�GD�盒��1�k_)L;�4�}����;e��63�泶B�i�,�VS+�3��-]gns�\9�ޗ]�y���1��<ۨ�{%]�/P� �;H�o':�:wzc�+{z9������\�_��,A���Bt�0���_T���YL�H�d����\�=�u��q���ܷgkVs���8k���Q��F��b��
����5�ku6�%H�I��o|�Y�j+Y�\,���a͉(���-�4ڲ��ҧ.��wt�<{���#��kt�r���1]隖�����KϲS���)�pu�S�g֊���N�wD,= ������,�oxM�C��O�Ggn���9�.R�3l�@p�=j��7���Ʒf��	ْsyW���wz+�
ź7��0���0[��,����;���'wۯsr�t]t��R��tZ�ܘ�a��-7��l���*м��vI��oY#���=WKhq��]�˞��<�[
������e'[��ouJL�j6�t��6���R��O$aJ���0E%�Q7M��+YFZ=5_jC#l�𒞪̵�ku��SP��z!�laIgv�e;uv]Z��e��}��olT=�Ё�*�*wnp����@r�좃�����]�u��d��RHM��_pß;�fN����vtb��۝N0ge�ض]����Մ����oLnX�g�u�zV�0N'���!G�{9���wKG�/Q����a�O[.�;0,����b��� ϥ�]��c����Xr?8No�ܲ�w��g�anٵ�NˌQ۫�wb�d����#�!��O�Vk!E!�'$~ޞr�'6^{7�+3n0�̹|�M�3v���!�J�{ӳ3?��x@����mWH�гY��`}����Q��ӄ\U#Q5,t �j�F��fn3K������<W)��9�y�CZ�jX����ɬ�x_z���@�?}|ᾚ��>�VT	Ǥe���t�F�hZxO�ƚ��>���^�ȼ��z�3�y'��e�Z{١�^yXH_�������B�<���L�j�At=��|>�⡦�P��݇����#���>���M��x�MF�|	?d��]L	Іޮ��Ȅa��f��5�!9�`@����U|tX�\#ƾ�9[���r��i׈=�z��"*9Q�ێ=���<D6kȅ��4}��Ŕ4�f�j��d�������5�A�����}���O��s�����5�����@���0���˔'����4л�����	�ۊ��Up�:T:hY�ߧ�<�4;����n�|y�>:B.��H�AQ�ۛj�i��P�"��>e��^��hf(!Z3�1j����m�9�K#j�;�����;��	�d޺T����QS��3.�c����)Ը��Mt�靸*�E��v��lr���ג�a�޷BZ�/R�C�'��Đ,C#*I���VhY���C�=��t8D��,���T!N�8�7�k�wyÔ/��D8G��C��>@cx����{�x@�T!���~V9�]#s2!�|�؇M{�_�q�sQ�&28��V�k���4�˒�0�mۧ9�vDź�0�,u#Ul;��t���#�,�#�D�|��E�#�w�����Єa���=Y\#���5���.���;�˗��i>E6i��R��-R"���=�����zY�k�y:���vz�T��³���۪|p�M>�5�?qg���Hcr_xl���/Gh�0��n�:yrt��3[�,І����������e�!�,гU����K���A+�;�9�;�����(�D���SP �j�y��DY�\���a���b?d`,T,�E�}���ް�CY��je��à���4]"f��dx�S�WC]�;�w<��[�����h��٭�U����= B��{��O�Ӡ}�|�~8kM@�؃"͑di���tqІ�Bҡs�0�E�Α�P���0�L�z�� |f=�V�43ْ.���y���u�?.pR0�gR{|�R{h�����'K#�0�f���[�^�{�.Ռ~�`|oʃ�����7j����U�ު��4!������e��MY�C��K�g�;>�V&��W��M;|4�5��Q��X���ceksv�4VJ[�4Wk�u�J�y:M)�n,� ʽb�C�{�|}��6��Y�Ѐ��#��Ĕ�;�Z�9��m�e2�������q��>G=\�A. ��4�z����#�QF��<7���Li3c>2�8������Qؑ�^�\�=�}�x7�v+�N��^�S��%:��%�3�k3���z콥W�ɕ�ψ�{�Y�1d�W�%bGel	E��k�j�(<�X�U9�Z�a�7]m���m�Аwd���[��m��p�̻��ڙ��;���ÊA�Ш	��%H}C����p�X�7�aG�Pޢ3����5
5��VDj�w�+��*���B��V}a#G>ޛ�R�y�5ˣ{{�tЇx��~č.k%;�拡��lz�Hi���ӋI�
�' m��1�u�i��l���}~�t0��p�Z����s�ψ�����f���,t����0��E�h}7�-��B^>G��(�����)V�~�<�x<Up�l�[h�Z�Q�DI�x��P�,��@dz=�X�h#A�G�i������P�X>������#��t����l�MyXB?qpп���f�� �A�F���j���5��#,ʒ' �dp�di�糜=�援��>&�@p�?tX:D5���:I�����+ Y��6j�,տ��u���h"�Z߸q��j�dߺ3��7eCAL} Y���dC^�>?�r@�!Ԃ�a���7�`Y�����F��j����wK.LG+ӝ���B��H�����#��|n�:zYf���vh}>���]�-P_GHٳ���Ǽ��u����Xכ�PV}p[*��º�i�F�J�]n(��9�2W������<��*���5�,Π,Րg�>6y">P�Gx����*+7�t��!����ދDa�|��Ȍ$�Ӛ�kM/������f���%��@�A��~|C��a�[0�n��]���F Ȅb#�����S����� �ኆmL:�����G(nИ�X�`)Ʃڝ���؋X/��w��G�F9v+�vOg���0���Ȯ�A���f�G��AD3�OH��ދ��ZC5�BZk��}� ���a#1���%��²�'Mc�hh�v�'w� 3A���p��*F�Ȭ�4����~� M��\�k�t�4.��"��s����CO��|v9x/��M���8�خ����q !���%Ͼx<"x|@�C�B	�\��;�>	�p��NP�;�4�M�F2��>��4�j���a�9r���k�s��I���i,�h3�j���T�����~���_[��44w��c�U�Ce��٫����n��Xcf;�g^Y<���K֝�wP@�Y���!�J�_�CdY��^�<r��$�F��3�3�vB/�z.��@Y��Pzk��-4�����n���p�k�|0��u��/Ye�jh� e!���M��]�w;��35��.����ۈ�ٴݭ��N˔:i<��{ i��`^*��Vզ�4.GB�w+���Ŕ;�A����a�O5F�獁~�;�f&�MZ�VG�s�畉iN��FR�F���|�*H�iqm��
փ���x��'�ϭ\ p��po>6�����.�"���U��G]Yׇ�b� 3|��`i�r�E�� t�g���H�w�mtF��!P�On[��n�!�FuY��+�!J"@��9C��|�#�aßy������#��VhY���M%��P���"��|>Hv�èX����$�c�e�*����fn%�RJP�.e���T� ��T��dC�`�r�)�pL�o�Ve%vspb����f�$�3tjW���,�M��@Y�,t��~;Cx�_mІ������a��$�-�} i��s��' ��c���j�a��Pеo<U՞�]�WՈ�4x�|��������G��N��{^>p�ShC��qW���pf����2`q ��S��a�}l}kH�������<�|�i����\�s	~��31�XD��_
 3A���}���A������}#MO��6�qWx�7�K��{��zk�JSj֮��fU�і��s.XBp�ƭ��U²��l��Kt�h�0�y;���'Vyu��k#
#�=�}�豥��4��oP���Y٫$�߸2�}��$���f�֨Xr�����|:'L������go8ps��'���`t���yߐ?.YL��p� �[B��`Y�!�|n��;�=�n��+M4�t����A�Þ�`⡇����}�64�����ӤB�|}�zh?M�g��^?}��q�G�{�0�AD8kVs��e�U�uo|�X�,o=����E�di�6�WCH�!���g�n���CM3W�?}�_x,в�@f?�]|y;�t�Vt�1�f������a:f��B��:A�l���Q2�iŚ|i���"��gJ'~�@'���wn���C�Ua��в6�b��C��N���j��������)�\<=5��ᘩ@���#�|s�>���{iTΘs��݋� ����� ���:r���� 8q�GvtSy7��i[w�m�ƶ<�ķ ��W\�/���\}�p����ӆ��T9���V�f9�@ۆIP��]�
4!�!��{�t0��L�zP������\^���n}'�b�:���8�4���<l3�¸���~@Y��ۂ�A�4$@t�!����Y�X�s�p$�$�L�	�F�]�u����<Z�d�m���k�,X�-u�e�f$"�����_�8���xk�!�������hm��}�߶uY#�t�f��Y}��`s���m�zht���4!k�ٖ.�a�#ݽ�0����#ob����
�BiI����|������H�`���������ڛ��{ԍG��d#G����A��@��e��i�@`�*� ��+#O@	���S�0��L�C��<�M�[4S�@�� 2	�@k��~wU�H�8�M2;���҅�4�����n9�����DF��wxlj�f� w4�>6<kMEA���C^"	�jG�D)�AqW�Ї��g����Xd!|_r�p��h]���I��x���B�3A��^X}f��\��ѿWL��*�Rw�Rɐ_���ƞ�B,��"@E|4|B�xL��QI$�k�v ��egDa�#{�����ho���Y���}��#5M��P[�'Hj�B�h��^+��|i�@��4>���5�B�T,�F�?;x���mMk��e�!�[�-6��ҷK��w�F�tr
�Y�#��J��S,�B���M^Sn�W,�͂�	m��8�f��Nq���XF��#m�l�����Z�d��1F-.kS6T�Ѭx�4z��O���`��la�����l�Z^wA�:�v�p+^���6;+�����Ύ=��q�[�Ѳ"�ݴsspd8|�vMW�'n�n� �r�v` .���AV]X�k�Ӹ���z�0�ZB�n�͸�*�n��j�sS�K��8e��E&�su�mZLTff)��U��֬�˶'\�F��;d-���Ir�s�K[f��Yb��aҴ���~#do���|o��t�Mb�����WA�ψ���hf}�h� Ờ40�_4$�jp��c��h�A5W_u�4/�c���I�E�$��ƴ�0��V@�����t0����>�m��||hCL�Gӎ�屢�{�D�k�C#���H�y�;%�,�h�d>�ϕ��Zl� �x�}-��4�i����q�H`��҄��q�x@�Y&�5�3C���.��#�hy����ý�X���5��J� dn5�,�D��Ϳ��/�@0��Yn���4��ńk��f�#���N8p]�w�;ZI�/6���NO���8k�D��-4�'τa�ca��g��=T�C4�P����gMt�ar�#������}�c;�]3]#����d3^!�g�m%q�a�P�Uf!f�9� a}�~7ZA4��A�s���2}�C�g҅��G
�uw�}�u�<jȇ����^g�|U��|oOuW��5��V{Ō4:�{�������9��pĚ0��+�����(���D�w.�q�m�����kN�)��҃t�K��o�,���Y� !�<�����n�8��E��#�T���.��dCVв>5f>}�ɮo���tf��}��:p����CﳽV,�k2�6B4����1]@�i�!� �4�f�4��w�/�W^���|p{��yYj����onovh)�֍��xe5N���i�1�l��]u�vT9��z��]'�8ޣ�c��s�m��&�Et�C!n��;5�a��p���5j�F����oU�֑5<��@�/�4�#��|/W�Â���:����hͲ[���7b��V{���ׅ���#`�c��.�{�L�Xm�8t�Y���O��f�݋�=o��7�G�,�߷��F�頌 2,��}����S oF0:p�d.�FSzn&���pԈA���9��=���ߗ��?+k��4�����}�dt��B�y�Mxk��E���Pl������y��|� x�G��k��xK�=!5�B��x�G)�-E��a�:a�����P;���GH��V|@���8kH��jǶ�[N��.��1jߘ�B����t`�Ȕ@BM��+���f���P��[�w��XIu���c���)Xͥ��	��yX��`��)���<�.4�� 8j�ь�a}�o=��w�w�� !��z�Xf��uU����Ρ��y����L�hdU�M�p�����o��w�v*?$@BM���l֚�4�|Ci����"*G#i�`Y��E����3�6/���t8G;�<�����M�A�����3�]��a���|jj���Xw��/ʰ�Y��C9�8.�0��/�}6�z-���!��g��قR-Ē0��WCM`!���dN�綮��L����Y���J5]f����W9(���O��TvX���S���)gZ�Y[��z/;sV�.�d�.���p�bsc���₣3LN��8��%�d{n_շ���g8.�qPg0q:&��$��Z�(����l����o��`�I�$��x�!f���v�z~~��� �^_������?��ߺ��w�X�!��Z|3���t������UG�}û���ִ
��[��2�?x��T�!��=��P3��dG�� �s����1�i�}����t4�f�EL�E��/�l��#>�׈��Y����aٚ��=��]#O�cp�����']i\�A��j¯���}�r�%d�X�B`�`v��u�7ɔu�U܃��-����6]����D�H �9hx����E�����pXD�<�C^#���Yib�s���D�����z��6����j�+���$�_��x�P��4���8G~\|ύ��\4TU��!I��`B$�B�6����!�d=ϵ����]�6s/����������#R��n����5��͐'�g���� �1Y��s���#H$��x�Y�������u�iM+�싺������,�ߧ�.�*��n:���\�V#ǖ8�a�7<ȱ�*��B�X����!�;�4!������f�Z��i����uȓ`���e�P�8I�@����>�{/>�������n鿈P�����<t!|�(ϵw� Þ�JI�dY�_v�S��l�9���@ȀUck�� �K����+�HW\t�@��D<&��5g&�p����@���֣+y�e�L��;#
���K"�Zw������L_�Rw�]WX�Ud�������.&�!&R�!�k�3��H��4>�J���a�49G�b<|q��̀�����A��Śf /�tX��4��m鱽*�~ |7X�Uޡ��>��Ͼ��G�ɗ�qH�'&M�:Y^#0;1\�r��ծ�s�CN9vY�ћE���Q��Y��V6{x��F�/K��C�L̕��;�]/}�.�==(���\�Gg����}�������\5�4�qf�4�oM�����3^�c�T<�Ƹ�%�Q�[�(a���:@f�}�h�l�\�����x��H��A���4dC#⏱��|p	���*l#�l׌�A?�p�w�ZF��qG�ȋ�|G���� ��G��%#EG' �h#]!�G�=��`#�C�k�4=�6P�:o���t
�{t,���ky�$R�/Y=T:hN����z��#���w���b��i��5�CCw�>Dw�ˀ��R-K��X�B���T_���2w���u�W�(�Kw��a�����a��џg�{���#ln*�l�~�y��>=4�f\ޝ��F��P���Al͊��<|Gz�Y�/�Y�����26�e�\% ��Zk�!�C��@G�~�]#�f��d{;��z����߈����0,�~ ��g� 7rh�!�@�/1�;�yPb]�a#�f�> �a��w&]�ҷ�X��-�f�b���cd�7hI��E��(�z���F��k��7nq�{r��ྻb�U�Q��c�������%�g3:�v�9�XM���;���Bu�.�̬�lb2o[+
�;�+Ü�f>���P�I;�:�o`�Z�b\W��\�6��mҺ�g�֫%u�]iC���z2��b7��7��$+��SWf�`��\vևyJ��.�� 7��;��'_#k����+AsB���6�\�݃�����6���~�qΏ��X�Br�(6�a]Y�kT��-������u��fV�X�֬u���f��Y)�W͋�,+ɚj����r����hٵ��^(��383C6�T��]n�/{1��3n�cb�]��C��os;�ѭ�M5I.n�Ѱep<�\�-Ձ4]���r;����M}Zy�b��Ϟ*e)Ի�'V��O���Y:"�r	V!�{-�]1��_FS�"����-N�س+���G���ۼ�T\�-��y�*ķz�D�ݵkD�{s"!R�C*f�ݜ+s���;+�};��U}2N��Nf#+pR�j��w���G�����$����@Vd���b����G+�7��%�]���a{Dg;�%V4�����I`Y��e������
S�n��"粯Es�x
LXZ/.-~�@ˬL�u�T�����QAu�2"������s�җu�ܔ ���3%v˩��q�ʻ���-$��v��� ڇ�K�8�s�T����#Yp�	��L-��tE1�ce�Db�R�;&�1nR<��ZJ�ު�q�X��&��l�2�Rq�v����l����֪�г�0���-�^6;v�m+�kOui,�eI�%ׄ����43ƣnB������j*2OG3���û.1�e+��'	�v�d�4`KA3,t�.&B�3G3���A�h�U�Q �@��l:�B��`���A��sx9\<�V[u����G���w9�u�^7����� �����NJ��쩻fn�y�������<�=-��8ӈ��>���O�u��7��͆lf8̘�6��vx^[r�`	W�y���fp�ncou�x�n"��,�m�ݝ�4�ti��:7W���[�8Cs� Ʀ�&�8�Q0d��b��C"�0�%�Y�����L�0c �WjU6�{+��r�\�5�$fjQ�
�� Z���S�y�c���l�zy����`�v�lCG'<�s��}����EC�Y��' ������S�ܓ(A�쏃�@E�x�][�rY�So<�b��2J�[2E�8+r��웯8�ItMn�ua�)ɟ#]�<�I���.��x�]�W���,�gc�\������E%n�,���Y��I����Z�j���-����1`� ��S-�۲q<��h2ss�s��j���ieJX7�*��
㖓/���ڲY�al��K#���2�1��Z����j��6�v�C\�T�4��lc����e�ͱ�D�ύ�Ãg�7l:=�{9k�FJ�x힞l�$��G `9��c�����;/��4���� ۲�y岹����q/��K�']q���t�P�/J1C�:������]��@�ͭ4�3tB)��ZG*jb�r���ٛ+1mUte��bԵٷI��0ۏ/��5$�î���`��Ǟ�=�ѧ��&SYpa焽pF��m����V0z[n���9���of|�mx��0�" CٲF��/.����3r��c-��N�ٰu�Z8 4�LA�U�� v�ܦzǃ5��E�cn�[��l�2;Qعnj�
�<k�\KU�70���R4���<�+,�2�jn4XBDդ�3+���>����K2N���cnܚ3js;��j��ܓ03uGGY�Ÿ]Ʌ���a�9J�.�Yf%�,��g�P��BDۅN#�J���R.��dۂ�qns�6�a�M��VXg9p��fn��cb܄�<u�<l	e�^$�L�Y;��mͲB.��k�20��o��WJ+~ϝ��A \L����t=����9�0���Q�T�>�7]'����>����\&���.�L��+�u���t�����׫���� ʆ#r�����4�^0��f�C�a^i.0�{2�i��0:Yi�������3ZC4��Y��+��ugU9����DY��>�X<0��vqϗ�{���7|�C�t��4>������&I2[�t�x�����@CC޵���B�CC�Pd?u��/�t.��@&��ծ�c�s�z8h}h�G�s�,��AY�i0�5�����|h���5�������"#��0��Vx�k�Cl�yή4�@F��w�E�dB���B���|�����B�y�h�=k����@Y�o#��� x�O{�`,Zh!h�@��3	?�a�a-ʍ�t4���$���ʡ���s��2	���9�ɥ���;]O�.�⠚�jÆ��`��h�h#�@v�cD�L��6�>��n!�ȳ@������u���WӍ��9#���x3{m�-�V�����y��㵺��6�Y�a��tٵA���v!��4��c�8h3C}C5��7^"j�h�]6hY�6�����l���~��T>;h�s�f���;��H���4H�T-���8P28o�5|�c<��4���G�r�֑�,��x8;���{��-�7�a����K$}7t���.̺[��Q4q�E�}}.��%%6Z+&Ӯ�Yg��ׇ�=`k:��6�{�2���Y�㯹|���B��Y�> ���ഁ��`@Y�_U��oM���C�;�}��Y��HF���=�����`ŔnFw�����F l@Cߍύ��0�4-�����}����.�!����[A�w�M\CH�9��i����MxY��q{��,֐�z׏ư՟�F>q�$8�e(1��,��Z�A��0G|{3�������� iP�� !�m�����_]0��hY����C~��ǒ��׿o>\fsM��@�d���u������SD[Ha�rwy�~�,�j�KMY����E�h\��l�c ����i�9�t��P�Y�!�����.D{h"4����<p�"}���,� B�R������<م��
XG8̥�3�SeӼH�3\;��V��\F�,u�K9`��ʖ:�j�A�hi�hl]"H�}�����q��γU	�JF��|���|F�3dl�����}� ���-�����GK ��479z.��XEڡOy�#����b(��(p���Y�f�!��/�ܛ�8zG}�~��/
������t!j�w׾;C��4�� {�獌#ǆ�8E��@t���k<la�4��9��q��ᝡ�]���s[�p",4S��a�!���4���Fx��}ª�uИ�R�}����V_ޚ����. nTwF�Rx�����c�kT/sPء���tҫ���qT�C�-޳V)s-sH=sY �=���\��f�7�<l�${H=B�3�f�w��b�U��Ȳ4ӊ��<>�ĮH�!�$��h#��C��g81���0��_1��9C�>�8@�T!��7��4���՚�gبY5�fi�=����5þ/���s!S�jY����7CH��*�5{�Iu��-��A`p�*_!f�=�`9��ߎP���8p��k��/����ʻ��!�H�a�"��`6k����t#Yh8k�ǧ�����IԸhCB5[}c��ǘo�IX��������H�3Fj6�HM#��k�v8w)��(�ݎC6�0��i�Ƹ*���ф�p{���T>�A�u���ϕ��H��4,� �������׈-�C���CO����o�-z_y{�p��~C�3�K�`��lx��8�@��BϏ�[�>G�-��8ɎHr�"�QP��@ϑ�٢�i����燻ꆴ��B��9ݳt9�A�����t{�p]�� �D�lύ���,���\����ƸhCC�'��X�E�-�_��{��<��Z$��_�.��3P���� w�o�_�2�0�g'rM��ˉ����>?Z��w����A�w��f��=���������B�&����!T�˂�n�5�D0��=�E��{j�f�HO>��Gy�VhO�׈�C>�p��t��x���Kۢ���A���L]�g/T'�4
>����9y��F��`�\��J�<��u*e�0Y�XyՌh��	S'nΩ�r��Ar{��a��#��x��vw_�EȠtÄ�Ӈ �����$���q��B�_��h[P֗��22�ç�@{#�^��@�΃5��Ś��n��`x�!]���P�Xhx{��oC3:`����,�g���|~�4���+�n�;[�;�q����n]J����󼧳P`�y{e��s50�8[Y�SPO�S��C4$@Y�s޷t4��h�J���r�eN�P�A���=�;~���|OO�}��<�?,���}�Ƹ|kM��g�{�y�WY@��j�1��8j��Y�gH՟���r�a�ޣҏ����8k���B����@�Z��0�gH�ϝ��<4��4!����h��V�כ����9C����x�:8��0a�rg���!ъ�9�<c��W�6}�s��#����!�]9�+��A,�u-w�9�� ��`>��gb4٠��6]4<��P�Y��h{��>�%l�KM�Ғ,���G=S3k�<3���Y���N���;�p����%!©O��`x�*�F�:E���\�'˦�ѳ���T���ݤ,����ru��U�@����#��a���Ƣo��,B`m��H4�F5ߐh)>��ihr*ߺv�H����}���|�|�wU#׌a��w�;N��	���4���i�44z�kHf��K=K3�7�i�y$�4i�:� �tUϩ�>�^�.�j#����V�s��uuѹ�fG���0.������K{��ݛ�R��F�`��5e��w�ي�Uf�pMRIr��vuT�[?��ɻ��~#16c����=/+��z��Ì�!cq�z��:M��n|�9��ZK�F�"�z�[���	m��3=ñQ�%�k����(7]T�n�1���D��.�{t;���pl..{&�;`��m�v.��.8�(�5��v��Nv�I�th���d`��Ff%Թ�Jv3�^0�0��vGc� M٬kb��@���n�S�f��fT�4�ĉ�C���Mv�1�*h"����,CXk�C�@���]#�k��n�G7��k�Y� ���Ǫ��h�}�Mx�>�����|�49��;gMi��V@�a�q�'� �H�I��C?��,�~?3���;�q]#��tNk�W9Zhw|D+��Uso�v4�E��4!��B>�勮���5�'Mw~�]��4/��#���}�W��>�K/�u@�)�ŀZ)ŔlB<l����������G5p�4,�D8���|��zA�_G��^�@|!�Ä9�K��B퀈�,���{~6;j���q���"Op���Q�!-��*Ct4���|@���E���uW��i�Q���ڧ��\fP�Y��{���;:�Y����H�������`4WMz@�@j"���n�8y�����h3A8Y�$�����E4ӈqH2�Go�Y����3����.��Lи�2s�������=hO�<���~#V��B�H�>�%�5�B��σ�������!F��v�#���{%ϐI��ㄆZ,Ʃ�/m�{7�n3`��D�۲Z;b,n��tH\��:�s�G+p�d_y>���~7^�: H�g�+��X4�H��G:8��s�t3��Ղ^"�e��-���Y�^-�����[�i�qi:a��_}r�i�Ge�>5��������3
F8��>=5��c5��_gy��gH�ٯ�=��ZϷB�M�p{e(p�U����X�F�2��q]#�0��;t�d�mh�Sb���;�؜��P�壾�hsʃ#8����t3��4�� a��,�d�1-4d@�}���t4��b�}kc��,�F����<��cn2`H�"�5l��j��d�|pt�F� 2Ȇ���It4�i�#��z��t�F��[�{;�u����lb����s�c�P�MD4�x��l�p8�Hpea�WHG~i��[���sI����+V�;��5�q�D |l�4/�}��]��4���{�t�Z��> B�_�����f��hrL�bZ�5�77#xX^O=�}�c(�b�	nW���гA@F��Ͼ����Uf�D�B���\�ܚ���v��MY�U5�4!���;G;��C\h|p�G���B��rX���^"���4Пw��ߺ;���q�ދ�c]u��,4u�"70��uJF�]ye��k�Q�eev�&4C4άWR2#-�aa��,�d{�g��'�{��лT.!�(F�ܷu�p�d!�	Ԅ��1��ʧ�����z-���#q��4;ϳ��=�\46c�xhK��~M��7$�G��U�!���@B��=�pe�����ŘF5��x��B1�S{|�>4�4��6i{�ߎg��"���w��F�p{V�y���R#ث�C�5.��x.4h�x����7-��agW��Y�U��v]����C>�P�hzo�.����B�çA���v{f�1p���5�1��t�W�ʯm�,���5�)o��kwB-9�a��G��� ߛ�n1��+ݵ��˄sæ�0�o��`#��@�g���,�Cb���cB���rBBH���5�(CC�]����Ξ�3��{>���-�@�O����"su����T��B�P���>��,��40� �w�o9��Ţ��������8���Q�F�C?'�+�a$�r&
r�id|A��:@d�%|���CP��B3�C�;��{]���� M_,�>���;���;3��ä0�PhCC��wpi�h`j�4���N��Q���r)�<I2W<��������Hڭ/-�]�|k%ht@��5���,`�T�0fnT������,YN�6�#���~7�#�<lІ�(�ҿ��t ��CBڠ�H�߶���l�j48z@g�^�M2/���5��>��7 ��U�hg3�k!��P��*(�m�B�> 2�=3�P�����__���y�F�0�Z�!\�/�U�|�pX4z١�+4/���4;���w�5i$��A�{���2D�-�d��5���a�ѫ�G�\S~�.����i�	������_i{:{þ\�o��w�;�M|A������ }寜��4$C����1f�s�5�Ĉ�P8�>5�x�WX�B���gzq-߹_�5��zqp�4=��D?[�,�����9h#V}h��d�Zjȳ�="���ϼ>�2<��>k�.K�ӓ9�1��9m3����'����k-\�W���i�!>ք���ee��/:��m�_�Iͼ�FiF�k�0h3\!����|S�HF��r��j�j� p�}��I#����#���{��ۇ����s��q������B����V���C C�di�/>���]4;��5|(B�5hn-�|ɶy��5&m����YumC�F܍q�H�dY�ʓS`�+X-�5K��At���6�pv�#�]"�4�����#�UL�,��K�拮�c�51f�=�3J��+ �s�������i� i���sy�E��z� ]�7�����;@u���+ԟ���Z��bȲ�y��b�O��u���٫�<=4<h"9�0�f�]"/��4��#�����pX���؉����66�i��&��鳽��Zp���_�)��	�
$C���gF�!k���Ff�q��#��y�����i1��D��hoe�=��,:FD< C�����`����.�t�������K�E��\��(���,�g���Mg�Y�0���f����H�f�4<��;�l��CB�9�����:�Y��9/�Ħ}��N+�!��{�c�F�ݱ(Y�,/�&������cM��N`b	ܞ��"�_.�}CM�}�t0���Y�f�#WڭoӽWڿ�:n�#�TȆ��4!����ה4�F�"��49=��XF�,��3И�ϫ�d��y�%Mg7��B�n�u��ST�sDR�̬�f���x'�}�K����V�s�W�4]�:2a�lvH�<t39�-������K��:����2��E�t��AI�����I�[]�5��2��
����[�WVA^-��!�+Wn+��[I�8�av�E���<�b�ݱ͆��8�sϑ�i(q���hʺ,��-�֦��s��7��]n5��nf�ntg��뭺�[On=�:�u��:��8Q3��bF[�gt�ݻPv:5��㵜r��]�3��q����ukr^m���͞<q�J�d��^1K].lIܼ�0�pvñ��v��]�Ȋ%$��MB���X@%����t�~!f�4����u��:�z@��8xk���;�th�p+�hp� !M�@��4�=J�k�%�`#f��~��� ����B$pe��#��i�����$ٚ���Ǆ��.V`�ΐ�H���������C�<��/%x�o�V��B@f����^߮ŋ"#ƻ��T��x��C"�D4gJ��\lW����g���!���P>�~^�c��Q�.\�ȇ�����ϸi����g����A����E���h3��,гP�뿾V!�4u\��x�h/}�$2�A1
R7��8x��d�}�o���G�gx��.����hr�G�R��h��`>6F�VG���0���@�������n�a��3H�k�r��܈�j$���juh?�����k��x.��hv!�x�}�d�'��-7���m��5g� Y����XOCMP�G��k�+M�o��<u��#�xvP�W��<����,Y��j��Lƽyd�Ʋ$mq���$�^PK�X�Me��W���1����;��`��gܞw����g�݀2&������������dwC��A�:a�P����܈����oY���^0�9��{���V��vi�f�����x.6�MD�c�hp��XDp՞ZF!�{~��;���կ�?V�M�.:8r���*
Ňw���ß�J{�8�{�m�Ǭ֗Wʄ%�7����:��g��<�Z�"�﨔@���U;�Ǎgl��#B�}��`ˆ�44'����O�풽�w�z�(a�4	��o���6�fR��a�P�*���C8D _�Ͼ�O�Uf�6@e�G_�h�o�J�A�P����Z!���_^j��q�B�YDx�C3���֚EA��l1f��vƷ	1`��RK����}j��7���}�+�t@����\5�ZF��47uЇ���+O,��F�48��v^zj�3f�S^�ܾ|s��xW�^�A��-W�CP�j����.T%0��A`3���h\Tֽ�ۆ�i�UCCَ�"�F�����|��ݓ�����B"B�4!�t*�s��X����j�(�����|pLCǆ�����XӝUί�ŭ��==��o ��P��)�����u���u!��n7C!�����6^,g�L��(2Q�(�$�$���G_i5dY���l���ɂ�G�y��p���2<hϺ�.��C~�\"�= {~�6��%%����o��@��P@��gH��s�5����qW�BO~���Er@���)9P�!�:a��dr��}��}�����/����5�!z��!��3���<T��١g������:zx@����
�d�]���yP�����������!��IC�������5�-:{� p󧙪�5�KVA42��4����4���kkޙ��lGՖz�Z��J
Y#q��V�c�z�!÷�vݵ�M,b<�gw�2����+*m�o+�df�ٮ'���bt���d��k%F��t�j��.�W��]G�����<�"��}�e�MvXo�6�]��#芣p_cC._s��6L&�����ak�s{DJ󒾼���VIǕct�=��/�b��J+Tכ�yD79+%7{��V�����Gt��wBi��}h����q�
��T�m�7���;e�٭cͩn����eb�.sq��_��XOn^�.�����wV"R�;�;��oTy}2�Z��S��#L��ŗ���$�;����m�G����{7ne�ֹ�m�.�%^v�Vε2{N�(֛�xK��WjN����VaWn𶑾�`"^Нd�i�]�1�,�X.�H�^����������@�9��o�&��˨+5�'"�m㳽ak�&�Sέ����.�Tr��ő��ɩ��Y�N8�>ȡ� ��������s�Y�9*���>6�6�f8���v���̾���1���{�/�!ɽ�5���������e�+����{�,Q!��KT��;7%K�3���y�W7n�Q���b�G�o���U�KHhp����ۼ/�K��Yۻ��\y��<��%�Vw��Wk:ɗ{Ď��r�wz�u�nݔ�"���ع�gR��J�;�rẕ}W�b	�@����-qHou-�F��P�=&�+*m(�2w���m�Zіr�Ǣ���=�Zl�$��>���C�GbM�]�a5��y�O��	&���!�Oğ�B��x�w��s46A?q��YC�#d#C:mЄd����>9Cz�i��O�	�͗CO�@;�!}���dw>ɗ�h,��ƫH���,���T���:c�r2�rH��Y�gH�ms����~u�����0�%\��r�������>@3
0� Cf�ύ�`��7�6{����ϟj�ȫM	eO��0�#ة��������Uؾja! $I�`;���]M��L]l]�u�3HiV j4K�v4�#h�E�p��d���@�����m��#p��C��_eE��ύ��Uhu�����`y����gH�����4��C���X�5���-�k;�8hz�|�і�$R2E�4֐���#�}���_j����-{��e��Oʰ��vB�P��q\ w�:�Y_�E���{'ܙg��2����||�pμ��$�%�L�ܐ�Ng���g���Q�c�����xj�ܔ�^喏�ա^�U2�	��ɒ97�}v�<�e@�MT�	X��w\<���^l�xJ�s�g}�ŋ��
;�>e�x����1�����ݺ�9Π��}V�7E�ۇ�c��F���P��������H�<9�:�n��eM[��Y�v��X_� 0�3��˜q-/g�Q�#
��:moo1j��1pz�W��N;�a������2�q�q��`���=�Z)�D�{_�O}ߺ.�8g���P��VfF�ז3K�"���B�6�x�윿��}���b��MB�#ˍ�����gG7x��ќ�k�<���i�v-�2�@WwWI��f�|?4O��:K�F�M���e�ҟ���	��K~}�E2��pׂ�0�^��X�����h̙|Go��QZ�I(L�p{_-o���{:�wK���|�:m�����;Cu��`�%�O<�bo�~��׋ӢZ���H��h��l�:siW7��+���~��jԄ)�=�u~=�TYjP�����ou�k��i'�qw�i���
�z�0�%P(�m����0�{�{՗t��R7:�+/�]+�$��`�ºZ��.��Z���z�t���cP|v�(Zٹ����4K^���Z�)��V�Mk��+�V!��\�^���S�b�4/�l1��:�'��bH���vu�xo�|o'�Z�����Cg���3&��Pev�bM4f�q2����YLGM�H4��NZ�aK���(D�[��ɭ9b�$�h�7:U���m)	f�If6]u8,e ��2l^B.������_ktr;-礬�]����.��zw�k?v*jSGp�;ilO0{q�I�<�7��k-��[����B78Cl��oZu����nq�v�,le���-�ܲ��kA��>�� BK0�{cst]Od]2�4�*8 RA��XY��68�6�3٫O��_�����6��_@���q�]�^z|���TIݧ`�ͭILp���`<\��oF�Ʃ���n<��e��Z��]��f�������w:�y�e:x,X�Wu�ci*i'V8�ų��j���o;+_y���1�E�Swu2��~B�so��W���<��ǁ�W�a��.���}�u6�m��r�^S�un{}�����3-� D�+7oF� �fp$�v���g��S��OP�lH:`��-:���B�;���yi��O����s��o-g{\X����N{cŃ�y'	�9ʍ'�YV-�a�[ew6��&�[6��q��,0�9�&T���rٸ��������?N����q>�>K݂s�� szi��w�o/O%��<V\0�밟�!�]n_;0��b���pd��~ٙ}����K��Ѩ���8'/P�b�-��m���&�������+C�����vAO��D��J����\	��E9���Mv�K�GL�R��-J�e�%�����5ɚ=�*o=�^�a����'�o5>�8R2��)8��%��nV.[��}�A�w�s�pC�k ���uӳ�]���!؞{����t��L"�O<{3ď���;�~�իK]�����m>w��u�4���q��g���0�3���p����f2�r@�l��lA�<ݻ��ίkW}�.?`�S������gq<���q�v���b�ӄ�D�po�']5oN��֟��!�a*�+���8�XCJB�t���ˍ`�2�̫�2@�
��V:��F�
}�}�׮Ծ�y�P��Yj],vy�j�\�N��OWAǽ�u�Ŗ1k̥���-��J8�b&wӸ��)}0΃���G7����V��a�
�/ڽ����֍!�3ۨ������kb-�	M��I������,�H/q������H=AX`�o�,�s�1�����(F�i6	��0�\��`yͺ�ivk��ά�.;s��N�M�U`R�K��7qV��R�VQت�����V��=Y��(�S�S�BI�r<�?,���k�@���'��S>Ӝ�n6���)�ב�������I��]ŏ&��7�u>)��������ӆ&ILfhH篮��8366+�І�����Ӡ����f�-Ֆ垼̷~�j�s��!����]g	.@ɑ�-N
�=�3��vy5��6�<����y�����n��]H�F%Gb /�����;��߾����Ӭ�ĢN�q{ǉ��Z����4�w��!���݆.-*4U:-���Hk������tV7ks�/�6P,�:���V�c��>��)�k�����:��Q�}�?w�߾�]cr۸��۴��Ӣ��צ�[��-��tb���a�~U���瑿�X�4t	���F��g��1x#�wd�m����� �X��
�-����eԫ�`+p#w�`!�Nǻ��JZ:�Y&����u�D��y��*��ﮅ"�����(��M��_fJ�Q�{��[�%�m��E�S���N�H.�l�M��Q7Xs���W��3[ \o�Y|�z9~����-�]�s��ߖJ^�ޞ�@�"TH0B0W�WGeҰ\F���-��j���c:����@���-r�?=�Ρ�u{��t�,�On�;=z9^�}L�\㗣�h��#�D �2h ��Q�)v���m������[� 𘝦�{ފչ���iR�Rσ�~�]�{�RA.��s�=E6�
(2M�1��=w�sϼ��q	��Y��1o�	W���v9_1�33f�\z�$RF�	�$�}��h�<���ɮ�ka
������μO0��n��][�}맅���S� ���c���E##!A�\��;��6����%x�V��_�g�!3��>=o�Y��X �5�WGb��Ohf���wS���^E�+��r��2�&�����wx�o0�>���'_Yg[�������wu�V�&���v�%K���.��f.%96�I)�����d�nI���f���I�dj��ݙ�{c!�h�^,f3���;s�<oX3���]lU]��漹_����s��Z�!�顛kaL��,cJ�-�Sk��WCz9s۔<b`�n��l��m"�d�!���-ymeҵ�6���Ry��er���۷Vx���v0������ga� ��Q�W[��nԳ�l8R-�����W�y��� �峲WQgp8���3ͮ7R��d{�8>�=�8D}�=W���K�w�ɜ��c��[�]xƯ3��5��/*Z��{�y�?~׫�C@�J�|���*���мѝ1i�@F����9��5\�#4z�q�Y+��y7���$�o�D�;9೘yVrH�M��tܓƇ'�><���W��b�&l̙�bM� ���y�2�Ș>Q��M ��
RKϞ�}��5�s0X=8י��7�4�oc�ӕw��1=���=I�eC���К���4X�1��1m��E��6�t���|��]h���k�%N��Sq&�O}�q������7��v�Yn���XF���XD�E�Z�BbT�]-q�+4�6���vIX�.��	�y�U^�̹gz��[�NNe䫯�����b�eL�/���⼿?5����H2�e�I�m��M��w�ڏ?Z���="���rp��5}`��`&8��n��t�Y������QY��oFE�&�$:����j
�V�{{b����W]*���}��{Ov��+m���eҾrc��=���j�%�S���׮����Z�˻�x��!y�ެ�eCw}9K�\�����{^�^��|_��r���yg���_%��(H���?W�ڳw9Ϋ�H_t�-j�S��{H��\:yP�d�q{\�<�zs|��R-���A|Zl��i��HD�-~���^�7���P�6H�z����c���ǆ�7w%CϗZY��.���]{s��^�G�66��;]��/��v�c�iw�6� l�Aث����˹am��Ƚ��.�~���k��+�Q̃�R>[��ֻ�-�V�]�b{㞈�se�1��6�Ӣ�a\D�ǣf�ʼ�ټ2\����jy?crnM�S>����������ߵ^� Y�	��Y���U�����
��f��'�ϕ�d��_��'Y�KU���Ը�T�r�3:l�|���W�S�Õ��stU�: Wv.�gvw�u��� ��:\��9������:�Cuڙ(����2��)X�uz��d����T���M4�,�o��o���ν�s��^�����rY��xx�7�:b�ߧ�A�
6����]�7[}\CO晠��-�����f�G��~�گ �^Z���\W� H�u�]�^D��][�k<�Z:줚W}C7�Ȳ�i����\�M��kr[kk�с)j�anyR�j�#SP%e��`V~��������{8m��V3�C:V�Y���g���wq���\~�f�t�s��]�\���z�NANA޽��{E��xB�3��]�~5�X�j1�=�Z�O9w�R��WO������K'A����r�E�c��ˍJf)`��������Vtx�ix�zT��)�]ۨվ�#S5,�\���ٳج��+������&b!�X�Y��;��珨.�=W�O�i>TE�Pa��ӻ��-vs=�m囩c�B{D����\
�/���!x�Yu�Ğ�g�8	גV�Ю����r�52�T�À��b ͇�ˬ^�to��Z���� ͓;��y���]��\$�p�����{��/�`OZw��Ur��w��stOw�N�h�u��ؙ���T��>��"=�S����̑�QYfFUcm�4՚�J6��[�n�f�1�9I��)70nf)nT� �4�)���Ӟ�Yu�էo�S;}�;��LE�x����	�����O�ۜ�	��o�3���bF�^�6�Q��x�c�w��ջn%��͞����7���j��.�ŧ�����G��.L���*T7MSE6Sh|��yYm��[����=�=y�Я����i�SR޼sk�!9+��ߺ�W��ۇ[,̱(�����p R����幂<��k_Y�`X��v]Y7�h�z��]{Y�W5bbf��Q7�-	��ԃE$�MP)��i��gs�Ӡ�b��'K���%�бǽ�G�o$k����R睊<{GB�	�=)%��BY.yG̥��ދ4�� 3��@�Ȩ⭻�&��/����"2Lj3�������⦡\�������0�M겣�b[Ya߶Zǝr�����ݳu����kv��1:p�Ә��Qj�j�;�.���o����=PH����VEM�3d�tP�&.�l	r�fv���~-��I�����o�np�q�ҵ���Z����:F���/6�ok����b�qz��k,�KSE�m�c�����"��[Sb�e3�J]��"P��������x�f4�^�l�w;���|,k���\�)7�4 39�JGa���K;��ͬ�Y -����ƞ��P�x8gԱ��-�|L��wV�l��p`{*�Seuݡ�.�J�2_fo[��U-��v#��&��.�vZ�^�52VNY!C����Uit��fRo%l$][ޗXwgI�)�*B�
���0�����KM��;���mfȃԷ��o-�()���1; �Ta:&�22[,����}�vdt{�am��|Z�K}�zۭ���ƁaKVa����[�����r>��$M�>�5�M����1O�_]�NS��t�l�hk/#Ԯ��j�]@���f=���4t/��[�m�굻Y���z�mI�O\�hV�F�+��o����|�v�ƣ�l4���Ǽ��[Vi�b�LL@�ӷo^�u�W��ܺ��jW�f�"�����5B@}��-��s{w��ޣ"I���$J.!˵f�4]mĺ
�l�
6gn�I�Ӻ�޹n@P��1l� �q�.YV�����O+]�R�	�tru4��輴�W�n��ܫ�f�eM�a��+��Od�ۮ;�eݙ�#��Z.1�<C�����!,hm����عg�`g	׶��	I	�:�.���K��\=ȴǁ��n����C��- heR�8����*U�Xr���i/l�����=	Ӷ�.�us8!*�й%�<.]N�͊�f��F�.���c<�؍����Sc�s����pԈ�H)NV�E�%�U��W!a�n�>ى3���<Z�hAș��Ή��u��p5˸&��&uܱF�!x�C�:�]�J�m��}=	�� �xb��q0T	�1uvU8{)�k�p<:�86�qעǣ����0����7
7���<[�Ѡ�Û=��h]�lƊ9 :�D�66cAu�n���f��q	M�p���.h�n��b�vM�������(
�����G:km[W6En[X˲F�.9r��[�I^�2��F\�.�C��^��&Ȗ۞_�}�޷�\��>�ԿkY�&�WZ1"<v�s���JH�P-�MCL�Zh�����7M<�康grG�W'h�pp�"&�;�%/]���m�!�s�
s�:�"ërG<�E��-c�˟z�\���r�c����mZ�^]H�f����%���c���(D�)�m��������]���2Gg�����g&�#��L[�a�����Yb��#c�%G'GU�iv���f`�>�`4un���7/ܾC��N8�MW�v�0�]]�k�j��;OX�hK3XJY6���&F2�# �`��k	]͊��P�%4��pz�� �1Z�_YY��q`�\��U�W9���;pqѕ����\.6 m�ۊNy�cC��N�!�4��O1s��^���9�����г�6��ѻ3�u<�/k��.cϧng�l;ur�v@'���m�#P�2v�+��.�s�f�i])+�3d)�Ӹ��`���/+�gg�"���s�ݶ��e7ؒ�xC��+	��f�Oc�0��c-�SV5=X^��G�"�v-��<�c;ڰ�.�ݗ��w*��p7m���#l��]���1���ں�Y�0G[��I��������G���������;Zv���u���.�v<�֜m��*�;��5R��-�ݕՎE�U�q�Į�v�K�u��e�Y��)R5%-�fa\FL���������U��z�Z��V܇.�_g+C��z���������3�u�oz<���a��I �=���e�m&Os�d��di<��՛k�r��NEًzW�7��y�[�o��÷�JC2{���c-��[~��C0�J�t�����ŸC�ν�)oz�G�:��:��uu�=Ad>�b������Y�N�T�t]4�n=��[�.�'.��r�Q=����̽�7��}oj�'�iUc{sly�J���ܻ��e$�T�tU6��ɏ�b�cZ��9�Xy�u��d�y���gqr��-�N罚��u���N���zŎ�y���)S���k��u?1��b�\完K;ɗ��s�sYW�g�ρؘ�vlE�s��õ�c��$$�o:�#��OeOy]&�.�Yy�ĦЩϬ��'M���.�P,�T��xi9ۭ���$�H��d�ά]�[�C��w�Z��)M�Q6��fa�b��b�K�n4���	�,���٣%�]��TN1��ۋ�z�'> ���Z�����@v5�˥�z� �E����]��q�N�ܬ��;;�����K�+�
�1e�.����6�sn����&1�@�1�rΣ��R�����}�)�ە�;RWv���h �h�y�7�i�9�����%$
b#$Vl�m-�==Ϭ��Y�r���ιB�74?.�>]�=��o���XY*�z�n���AI���?wp�}�i�0�	@�n;MI�ܽ[�hF�jE!Mt�zg]���K�i�7;���\e� ��Y[�#qga�$�!�QQa�Z.�"m��v�0G9;n�8��3����@2�"�D�W�s$�i:�$��=��b�`��)R��v��>ւ�*��%��JZ.��7��fv���%��IZVst��O�b���k����9��n�ί$�ƻ
6��8DT�u�=�gI��M�+��g���Y�$���gS����5*�N����z崥a잻�Ǧ@-��@bK����[Vփ$+�����{j�L�$������8)xtv̖�+h-��E�����FƗsev7yY�e�m�9)wfX\�g�F^�]�{���ǻ�|�U�wu�tl�#7��q##,i��X�cv���>M��,�T���>w5��]�Hkn��Zi&�v��ⳔҎ�-Hz�fK�<7��{g=��꽁��A!	RK�2f�{����Pڝ�C���`ֻ/m��x�nr/󇯲�YU��&pu/2cO�,�uK���%��C`�j�7n�m<j��G6WWb�3��x�aG�,�M�����Ac�;�\J�|w�x{���Y캺Y�)G��?j}ŗ��vJ����-m܈(��|�E.�[�M�K��i�^���O
�N���"�Z*5���nf={3����7	��m�(h��4P�*U�������:��\#�+�Ӭ��C�|�U���*g/�Yӆ��s�㫹�Ѯ���.�z;�^BIHaA�$���{ںޭ���"���W��Zr����\�	��)��������s�U��w�Ɋ�t��m[\:�_t�z��4�	\�r�Brc���BR�a�n�[6Gl8��z��w��ɕ��.��VƸ<���D�Dӑf�ۖQ��\'/1�7s�W��%{Lj���#=�U�=�"���T��͙��]��Q㕏ߛ�xG�k:�5�sP	X9D.a�����n�P�j��6���U��V:k�V�1��m��i22�X8�r}��� �7h�|׭[���+�����ۚ}F�d�l�k��*d������ە	pJm:��y�lŻ|;ަ9jFϭ���#5���j/v�~7ǩ/=�	�ϑ�;��j��\�����E~��RN�i�L^]$�e�>qo9f��Wࡘ_'9�NNr䮟ofV*��>sǘߖ1��P�E&��ގ�6���HX�G=����p���ǳ#��&�{]4��[� ҧ�|��AQmM��� ��&	���k�vN���F�%��h�ꇷ:m���?�X�D��w8Z�5sމ`-��Nf��g���2^=+E%���W �z��M;�I���W�As��\�í���vWJ��J�Wk�i<�����e5g�o��]��iF�n̢�P�qq�s�����΍����Z�\䗑��鍬�������G5�^�znAٺ�҇4\m��%�c�V9�ǝ�
�j���m�[�8�]���Y�,�Dn�,<�����Z��Û<ı3��z�s�'.�ZC����-�Wp+�F�.��
4.�)YGtkrm8���Ќ�s���N6\�
�n��v���7���\�"�u��v5�.�.��i�Um��V�,�ڸ���?�Ӷ��T#n4�a5"��o?6����g��l�ws�JzY;����*�Wψ���y8����nǼ�L!M�ʒA����o�8��͎�;/I��Ē;0�i���>��L@KH�mY���Ǳ F��!
	0
%���#̍���;"�k��"�>���J�E^�N��6���o�=�상|�Mg�l��"B3W��P��CZ���~ĺ���(a��՜'��*w�g���Z5>��[n��x��<�<=�s�:�H=$0 Z0X�j��OW]w���M^����Eu���u�Q�[|"�a4����=�ן^2#�9`��IH�0��B�݃�sT��\/T���@.��&�kv�ܐ4&#Aa�5e�>�ݷ~�I��X��7��^�O,,�1#Rſx$nϘ��KX�r�ٻ���a'�������cj�p�X�3{�,��&��qf�X�Z˷~�79f�8o�6�Nz]��P+p�Zy�gZ�oj��v�B���������3q5-N����V�#zdY~���Z�,X���Q{_R��U��U�`���T��m�_�����&_l��{�_BETb"L!���<��g�ֵ�$D����P<��7�=������}�7R�*�ԟ��ɷb{zJ�-ZڗUj���P���(��A�����#���9>u�kc�:���@�A-�S��&�(|��ܾ�u��lq珙�~U�������LU�����.�&�$���{�{ʘ[&���_1��$4mm�3�	��������ם�%��?#E�_�]����G��-�2S$��ۨRJ�A*���3�Įƌ\�Z�Q��; b;�rZ�r�DD2�&�D�l�X����?`���6���N��׻�yy�FN�����]oD�$�.A�n��W�/�T�/�֚�2����=�}�c���Y0�>�W\�+�m�^�j��ܬ�|!uW�ю��;5{�|��:��7خ���~����:�kl�W�n�V��=%#�1'j���n�f���+2T~�ia[I/b*�>����>l��u��$��I݃�c��f޽�5%��T���m�318D���N�;�a ���t��EFߟ
����"跼���sL:F���&�-�-��J�M^Y�^fr��r�y�*4:��+b���az_0��:v�϶`K~{=���|��r����d"����	�(\a�̉�c2؇o���p�RWox��!�-��'g�J��O7Ϗ�����ڽ��~Vפ�S,��i��u�����f]���;�k��+q]�s��sTK[�v��N�[��Ŭ؀�)�$�Ҥʵ���q���^L��0\�����5�ox���4�m­�7B~���#��d_��W�J���� �24�1�~����)�5w����c�c;s,D��Y�.��.T�����n}'�`��`�1:�-�貺!$�Y�9��{�;��˙�i/l���y��]=����]�guS���j��[g%���&B�m�(����hg\��oK}�/OTr��׹�X�y�=Jf��鼊OJ�R�gme�u��S/]L�	w���Y�J弔Z�/eI,g��z�)f�y�>���z�pMH@�N��K;�+���A�=h%�΀�7)�o^�K�?eL9��Tt��z�&Je2ӑ��؝�#����d<r�Ӻ��z�	w���/87=ܐ���3kp�m�7kĿ`4��g	�kOF��똻e�&� �ъ+H.֜K1U�0Vf`����<����*�E&�
��M��͂����{��vt�2�0^X%8u*�W�o�$�Wg��<G��x;�����RzqS��k��9ݍr�jQ{���=�ґ�������<�]���ã6eYp��.=B7%��+t��G��>v�&�cWO\'+L���#^Ip���������2T��n�T�����u�J�&v�w)3��ųk�r4J�=/�z��-������n���x6�=��'�È8�G	�
jX�ƃo{��l�w�(t[�j_T_?DE.�3���n�w�q��_����6M�i|7Fs��~��ӷa���@�+�C�A)#m�xt��7k���^��@�~�!���ޤ�yv�7�0�R���غ[ԥ��R�8˳#�P[7=�y��;U'�]g"#`�
x��:��D�V�^C#Q�C�=�9�1x���VW\�ߝ<缏���Ɨ];���}m�{��lD�vL���֛���w5p��ݥ��t�X�# ��`.N�#av���
k%fɒ��&�x �8L���ە��z�td�s��fhě�܁v�zq�p�V�=e��wnyu�uj�=]]��7/c�<�iL��o6�Wm,7SCK�6T�&��v=v<r�<qË=.N���/5��F�!���v:+a�`n՜4]�F]��)�ej8	]^	�W3Ԏ���՝kè��΋,�\��:�76^p�펮�bLfb�Ȝ}����ӿ/�����wq+�����(�e�J^����8Y�}=R���w��so��'}����D�/v�����m�"�b�M.���/2�ѡ��:[tNJG��ǆ&�r�w����J
j���ʈ���af�`��4�����{{��:�Mli4\p��=��,γ�x��I��ڻ��e5��y��l�`�>�jX"]m�K��;q�ӏ��S�%���Sh4��QD$ܿsUj��
��2f�ͺ�QӼ�ybN�ѬC-q;�l�^���:M6�����&/��od{l9�&iC��:$�r'�D I�֖�yq�^��rℵE��;�EYFT �����S���Ms�X��Kʩ�L����+ق�_]Y /!;��k�`i�F^�������)��8Ý��l����8��Ô��d�3mf[-�s
��y|��l��*[�m.�f�ʻ۝]P$1O�|����k��k���d?S��2Z��N�7�nŤy�cl��)�`�6�W�ZF�j�y��f��Gg-ߩ_�K#�k&�:�.p�+;m�'vTf
̆�kT1φ�w;K��+�9YŢw,۫w�N�������
���,�ݻ��*�mRƯ�|g��j�|T�s�:�ܿK��S����XB��w�lY�}����"qb���VH�" Y�=��jv���_��s�������ek�~�`g�r soW5A���h;�;L�P��/����֑�i�5�g����$�yCHi��}^/ÁH�]�WU�L@B*ǅ��W�o�z����4n��uS��e��T�ڪ�^��c�s{���m�h�Es9���\�44���cu��E�1@6e�r.�����D�� af�H/ڮ�m6�� ggi�`B×~v�\Syu�H�j� =/�v+9�Bb��ShWsۢ�����H14�5B������~�<|�_!��Cb��tM���N\]v@x��72��71�XF;��b�.��L�T����F��4+"%����LﻳMi�Et��u5��K�l�6]̙��7����Wp���z5]�C�CA�*�6Ef\�u���ڠK5�*�۾7H�d(�@�%�@i��d� �(��zt]Vj�y�~ׄ��D�5�e
�TM7]��T"D!��� *�ߕ׮��w "�GH�hB!��.��4��������f�v�>��XH �c��a�H���Oe�T��`V8j�#���d
�
����S#�\8ha @�y��	���ۿ G�Q[�x-��2�{�x�#4*��M�ҝy X����9������������j�g��Y��X��\i�����B�G��4������ų=f����]��7.�Ѻ�w�R;���Z���콊R�U�BH��;�{P�׺)^�Y�t���h����a!.���Yy�	dΉ���Y�s$`l�Oy.���1t�b!u�]�R���T)�r5��Gf���y�ݹun�p�l+�g��3z.jUrN�u�����F��s/7+����]W��l�5��Z�ů�[t�o�����&[3�Z�����_P+�I����v���@��#��\�T\��ܫ�Y�Y֪�;ذt�:�'��=�<�%cB�I�Z��Ej�3�.<Ԣ��3���߯�Pm���o�����o61S9���+�s�Wig=���4vgY��3�����y�xj�[�5B�y�e�yF��y��dz5Qղ�S�g)�\����k���&em��� 9�d��Jh������+��r��N�p'Y��jS"��فd��ԪXY�պ�|U)���5�]E��]�YJXg-뱛���8��{��w1r��\ϛ:�� R�Ɣ":�A�#aO�
{/����0�؆��}�;�mb� լ����b�ȡ�a�!�y�^��lZ�����5V�Om$O$��j���hY����&��/.���M2eu��8���� �U�Ҧ��{�;�w�\T�m�i����fV�j�3�����2TC�wl�Q��3|�j�W��O&z�e � "�F�}PҵÞ@i�}�`t�4�ӭ䅞��r����W;.02�}j��:@�H��7��\��=�M��@�EU篊���@�hY�X@�HBE\��X�1xi�Uf�w���"��B�_|���P�CMW�@x�x@^�� �{=�^�M
[��<�Ut�htІ�@j�	�y�ao
	
)�MȰ
D Y3���(��H�>�z]��s��YP�R"���Xz6����t+�� ȩ�� @�y(�|�"��\45�(d@Y�"��ߍ�]�n��@��\� d vj�;����A�t�8�(#7�Ų5^i�c���]h��Jث�FX�i��ۗK��2�n4�$�䞠<k���vUaU�
���H�ڬB(i�P@�"��3T�K�v �#M :j*�f�C�  ��V nՌ��w @���j�Y��#MP��l�VEVTH��� T��6Ӡ#�ȓ�ֆae�ZnE�(aS�hP�@hCB�@�zy�A��3�*�î?o(�Uz*�"���h��,
 i j��Vk��D�� �y邐4H��4�P�Ud
�:�<�U�C�S���:�ސ�:@$ z��J��(�h��nQMH�F�ʪ i 3UA�ZES P��^�P�H4+X �MY�+��"���K  U��t�"�5U���凖0T a��=���ngM��PY�4B*�hCB������P�vE3@YA�[���ߌ2$��!28�Z:j�"�*�n�s�5��C�P s^yتhT"���������+<@[| hhB(YU���F��}w,Y���T8hP�	�UT��]}U�l*;�eFh}ԩ��Ӈ�_�֣�':�*��(L�G��|KVG�] 9�6�i��;��ulBooqsh��e�lbN�r�K� �٪�<t ӆ�4 E�RA���C�W��#50�� )��'��p� S5z�
^B��r͊�Zh�TAqR"� j�'7<�|<�H3FwpX�� 
F�R48j�"�]����p��T�ܴꀲ*�Ea�4$�뺪��t���5TH��@�c�og���glt��C稅&`5n ז�eG.���4(�
�S`	D�s	c�a�t���Y�N:�l7�r?i'�$jEP���� j�\����t� t��@E;==��"��,�En�h��=z�EU�� H��*��_=�t*s�=�1�}�@CB�j�dh S5T�7�� �5���U2 �*��y
����6=��L��D4cM�t(i����U��5\5檀� @��tء�T8@�~d�>�Up�&�iH�4� N!B��%�j���@�P�E
FŪ�9�WUV� f��  H����y�rz���L��ͫ�p�Y��@�;��N�:��~o��*��g]��$- 4�$�� � ;UT!��⡋����� p� 3P��T#��A��8@ԍ4+q��R5Vxj���z����xi T�UW~޻��b�� |F�45U
�Ϋ�B��C���!��P�@CB���ΒC@��0"ar=�C��h@��咰�(x�DU^ {�CM�@	"�m !xF�T��wUD�qtС �!!�  ���b��T ���XhYG{�3����=�EP�{��zt��@� �T5LB
"�>����B�16�ʨkMP8�T"�f��4�}b��U�s�r�顦�@� p���"���w��k,�LS�����uX�=Gƨ@��U"}��PS��uT:@��UL�Cް"��5@?s4�Dhh0��(#U���j���5�,n���w%}^0�d:}�^}���kf�J^2/V�Ӥ.�-뫗z2�+�J�oe�q���7)��9��X$�Zx��;��� v^V���������6���E��Y�I��Rg[p	��l˽���N��D�RT��L����v9��Tv�X�n�l��-�8�\[puҒ^��5]bul�&"S6v�;����b������ǌ�v4�Mů.��,#W`�ebV�,��ːy�rn���<r'&����<�<�q�v^�[���L�	��p��g���6�'g���nۦ�l�G,,�:G�f�b3����ά�f.bp\B芎�p5��I��E�����_�P�a�B��Q�0>�>�@�4� @dCTT9�@fv��a�UP��5U�! �;�49�<���;�G�WH0�dBH�������~�b��i@������$ƫ ���C�(��4!P��wH����zWCHf��� nzqء��#���y��� ��І�*E�z����z>� �CH�"��c�H���wT8F��p�$hV��X@}��;�Ui�^}ޑ�fwE4q�d ��{��Cj'�RG�\"�4��@� j��ϬW,�8n�\"�B� BM���UȑK��NU�E@���_;�H�b�j�Ɏ�V�DwP@�Us��u�+�T,��O�9��r���#
r�s�۠0�k��4*���zIo�Zj��t'}8.�5�:kM5�+{{ �H���� �	,�Y�U���j����s��M[B��#B���I�������uX� WmP�5�a�W�y��1[	p�kW"�в(LB�"����2��@�!PՑH�4Mt��*�sj���\�9�o��ǤP�S f�J�H�81��Z��X���4��{��t<�)�
f�1�Y��{��w�1���\��AD-4"�5VlA�F�v��IlX́��X�Im���d���ͫIf����n�9>���UYj���ȳ^�o��<#�B,�]�ad"c���Zj�4EQ3B�=�|/;���Y��?#Fxk�44օ�s�� ��V,�@�(3C���i�<A��!&A�������f�"����.�p�ʀu�^1Yyt~���v-�j��l�����W+ V#��Ҏ�l��$�\����ڷ��s�<׼k�7�d�ݜ����|T�����ۜ�U�Vhz*� ��wH�0�I�i��U��a��;�ȭ:Grd}#�������-T<D�U��� {M�!m6�0��R+�0� ;XD"��(j���w<lV28�p�F�L�:�n=�qjȨB4-������=�/���=�03�����;d pЄM�YF��(9�;��i���U���"�E��o�!R2�(�P4�ڮ��=T�X�w�o��X�$�U�.�e�4�,5x�t֑B���yء��8j��#0�P������p�=���U��>��z:"�7�"����B!�"}�r�������/rs�9MhT#sΫM����e�@C�Qh �f������L뜮�e�M�4�F��6B5onP����R08j�����}�zX
���~uP�^UP�����z��m�Y�l���.�U��ͦ��:�ƶk�Ղm���EyC�c@�B���,�
���bp�Q��] x��uP�B����7@#[j�44<G���UqP3��t�5f���@]�0��w��ӜZ��]��o=}�4<l��4,�%�3�0��C�#�Ȩk�3H�y_8M¡�2c�9S#MS ?)޻ �G�м�-�5�������&�e��"�󥓘�t���b�a�7��`�i�0��ha�*�f�y�x؄Z�  omc��[z�`�f�H~�̲15"�$��+��<�Ȩ{jV�����{]i�@h#H�P�������5K��3J]��¯5^�KS�k��AO��B�RO�R��.�Z��s��yr�t�+��:C�24͓��$f��2�ݪ������,�|�V��[��!�j���f��������t�5�誹h2MU�h;��T�)RN A5��۫4�Α�����O3�{���$\사� E=C�3��SB�a�q�W�+�����B,�"�wy�������mڵXhpZ���b��ZJ@��H���,8 BH�ʭ5��D!]��7P�N����5wP�߽��v���C��/PDY�~!G�;u��9�C5�E����`MS"�T��"Z <����k���!�	}6�R]v9n��w���:L�=�u�B�6�Z͛�\�&�q��!g&�Y���}�6O�"8��Wn��t$ل#[�%a c]+��јA1�	w�\�i@&�[ �a�Bp�x�vl��0� �F���VF�J��I�� p�T4!-T Bl�=,2��|;��ܺ�g� �6���M\�
���ǵ��VA����@z!{n͜Cf{U�#�H�:��^��嗰�������y����W5b�s��yy�/�2��&�}���!��D�M�����az8F�����P�ն���8p#�2�a1�S��}���6���`��Yy�/$S�%��p]i�6���Z��b���O�����B��p�⎄h3P�h�9��4���YGF͘i��|�t�ʴwN�[]~�m�R����ˮytz˙]����s
�ې��}Gs"�cx����n�	�\&�����}V:��͙�`}�v�doF�`���kna�uS�϶�9���H�L���w�^d_UL\�j�4/p�a0�]��qy��{��P�=���)�+ơ��?!\>�x�J����dS<��vŚ�לD5�C���e��m9���i&��ukj�ԛi\�GJ%�!��:�[��t67�Uڎ��*ٲ�d��xw�xV�Q<�z;�u�
$�q��|e.nټ5�Y�4��{����%���VE"ט.�WTu��U�s��"�-�y�#�!a�7DI?S���ٛ�=��}���E��{��#F��޽5��8/�� �L�@���9�8��w9�;�0�lY���U�
',"�v:�3#aMb��~�l���!�Qi�y�rŎ���s��T9���"��Lv1��D|�l�]��ݣV�av��#1�"�G�����O��Z��t����3e����@�"��u��:kP7[t�ϷEq��R�ʽrF3����-GH0�ab�v@��\B9{y�wBQ� �A�$���Q�C�PE7���~CQ��m�.�����ϻ��R��U>�/{)
��`�\,p�!���:U�g�.%�V��z��0n�$o]�[�=Ռ��Y����"r���@��zކ�}�%�&�v:KD㎙90B�p,{Yλ��R,vU�ε�D��.�&̏i����Gj�p��WAG��D���L�d�ڌeu+�ntҶ�-VP���N���8�n�(X��FK�GZȴ��V�[�"�t=o�����Q�2���F�����Y�O;���<�0�B�8�Bʖ�,&K�i+u�71�E��V���r��11�h����xɯi�\m�.��m��xD�1�'n�Nq;��W<�B���1��9Ҵv��rҢL�sf\�˦`6bZˢM���ŀB������S5� �$h�t��Q�9��Y������~��sw<cFs����W�ea��uY��5we]_�gW��o��ۚ�\O�"g+7�2m�Fn?@� �N��Y��*�0�Y�d���y}����]�����ݝ������W��Afo����(�>i,�S�͖l��{�x�݂m�x�4,90��f�m帢*Cn�1�����s=b?L�p�sfi\Y�Y��_��4���\b��w@_��������R�寝n�,)t��}?K���c�U���v)�}��uX�	2��t���T��j���˫����-Ђ����G�Ge]e�4;��뫾��A�'�Ա}��A�B5���^��	��k�T��'J�ֻ��p�5YS|�ֳ��g�]�|�)�vP��,p��Ⱥ D�s�sV�o
ˤ����?�޿zw�7V���#]���K��\����4 0�.`�CP�$mҚ�K��:�ĳ�&�&D�q�x��}�f}k;Č�4rN�ߎsx� ��28�=/G�Sq��y�<nx�5����uɻw�{�:3��L.8-��_-8>}-��X���+=I��?r��0O ��74��"��L!e�ҸY<N`��݅7cR�8�v�u�n��i��VtE�Ofv�+��wΆ'�Jb{.�B���:�x��]4�*o�?���ݞ�V�z�$>;�U�-^���'�8�>�o���t$RP�I���r.s����������Z�-U��+�x��ny���v��s�ar�����yݺ��騽�����`�i/ACnS��I��"�M������sT6��w-o+�o�Ƀ��.U��pgj}|��~��iJ�=��S��/���Qh�b�{F�����_��&I�)fd���M��B�|�x�e:H���k�NǬʝ�R�$K��/b��Rȸ�1uja������-y/[��uu�s.�^90�v"��y�5�{���k��M6�ٙ���-���#Y�%�auY�޽����w��b�u�yH/����n��{��[@��G�9v��U���w�^w%�r����a��R~��ZE��H#=���\zF)���Yh2����
y�sYYx�c.��K�ȱ�ջS("�f]`���w��y�mҧ�pS�^�&��Y��E����1Ǡ�;�z7oУ���C,�l�4��`zTYvzS�[�6��$�^󓺌y�+���v�2����ٹ��H���,f�����n*Z�r�[���YK'-��"Gtۮ��i�bԪ�^�t�o���R�*��x$	��Be��#���zU�W��3�ڎ�Z����h"�.�ݜ2��Y����1��.����,E��PJ]�e�e0:/{9tW��eQ�7yc��pߢ
�PdH�"�'���/�}}����a���s�D�N[�ޣ{����).�;�9�~#��c��=?</�����|CB���0���Ů��ݹ�kG8e���7�nE�l�eL;�6�5W.9A�ϩ��6�����?dIo�
7oyE���3e��Y�j+�5��t��.�]X�����Fy��T��,�b�����F`EIH�
�'����;�>e���`�%�:Y؄���[�.bct���e��v��2�v��ǫ;�1�o;��~b��9ؕ{����I��-"��ޝw�s��ˣfW����yMe��w�s�J�De����K玻M��>I�;�|n�{e�A���(�l��+�PT��]��fI\{���Yu�Q	-cy�꘣S��={���S�{�v
�8�kuqf��(ʲ�m���2�R�S���L7�(��1��1&�ӂoV��[�G\�5+j�W2ʒ�[R=��F���B�~��ިQa"�i�E!��`#��������y3��2����}��wRs~P6��.�*b��Wɿ8���~��X�u)a��/�}���@�QF�Dv��1��:6��;���z��`�K.c�!m�\�1�%knmo���Z��F\��Y��1Q�8�"�.�Ip����r��/7�P�b�v�x�i��^�I='+�A-��P���S�+S����v=���ǯJ�$cvP^>Я���vƓ���Y���X~d�/��Q�!�"�:0H�0[��$���/�c��cCd�i�T�R{�y����X.�Sڸ��r3N{CӖ�m����M�1� I(�����&�X���Mfզq��R�F
�$ҪZ|��6��峳(%
��;�ʙ�a��[�M̼���L��c�%�t�}޻խ�m� �8^Դ��"X�d��/���\�|��g#h���*��U�UP����(
��U_�UT*�@UU
����*��U��UT*����*��U@PUB����UT*�� �*��U�UP���
��UW�PUB��UP���(
��U_�UP���
��UW�UT*�����U�@UU
��@�*��UhUP���1AY&SY��-���Y�pP��3'� b9{����P��@����
 � $P
(    P ��  U @�
( 5���*D�������D@��Ѫ�QJ 	PP��QQQ$*-��R��EQ"$(��TUT(($
�L�Q�U**��E��*������{��=[N����l�^�U�0�3q����@�ïkm��v�zu��������z��K��7!Uv1���5�w��E;���3s�)@@ S�{���Ǎ��L�[�RC���wYŐ���^���0�a�޷^�S�ouB��P�-�{:�$����BI^vz{cV�����
$kR ��@(�
T��R�<��W=���6�u^��l��n�T��w=P{j�zR��R]`�����r�*m�=�Qr�Z��B�JE��z[E� (--���eJ
���U)�R��:����A)I�d�(\���)w�䊥C:T����/mn�z�^�-�綊�j������۪��UH	 
��P�P����)��������M5^��s�����N��+����vbޠ[����Z��̭��c��*���z�$�.w9J/mF��{�lR��n�����]Ҕ��(���s��BM�r��o
�y��m����3MK{�<����m�����tѣ7������)ݹ�P�+�Ji���(���{ء��@Tw��J()H��$����q�Ov�^��I";���U�2*%{�� �����G�SY�;���l�{t����`���R�"�t�Vh;֣�s�$��XA@P /[���U\cN6�$(�;ʂUޤ(H���D��J�\�q!ջ5lՖ$J�9d/,J�IIA�ǈR{© "S��I�2$J�{�/&AH���
���ds��@�)�( R�瞚�TR%T�P�Х *�m�
UUn��z�BC��Sg9�����J�x�U�S�Д�oz�Ug�*�IIqj��UE��/)E�:"��P�8إ**�
^]�J^tR���&U=e
{`(x��x�@  �C��
 U�j<�{0�T���ǕIN�I.�:^f�RK��x�f�[��R���m�E%O.�T�Y�(�j/y�^Z�F����ykCq��-�c�{�zڀOL��*   "�`�J��@ �L�j  ��D�J�4#@OĩRd(   i�P$�&�@��l��V)M�j(�� �'(���qD���D �99{��k�賫U�k��3�ř�I����ĳ1feŘ�%����f%��3?�31,�Y��Y��fb��b�X�f-����?�O裷�+�n�:�q:4����7�)⡃�ku�GwS��J`QcA��n�GFmś*Kk�q����,�u����>Ʌb�e��Fe4���mꦬ7eg��X�u�"��R�h��]���.��Ʉ�ɴ�ӡa�,�*�s0$�aLcY@�^YՊ��J;F�V��f��FJBؼ]�6��!��s�^13e����$ �-�К�=l̓UY*�2��N��w��z�r�4�2�n�jq
ۇ.�B��cuR�~��,n��̵M�%2LZ`�Ԏ��X��������!P��82�0�L���SY�DQV8�m
d%@Ɇ��B	x���W9,)����y�eő��['!����
ܤ]0�֬�V�.�;s&�w���Ԅ��*`/Ru��Ԉ�Mc`˖�݀�+�e*Uē�+(�C�Scna����FP�����y�6e��(=�H�^�22�sL����x �c3eM��4���&�U�hŘ)�cd����
g� ���,�t�9�4JJ���m�%1ݠ�F�{-�U�*��ٷ�-�w%:��d"�Sc�	�G �Fa��1+�t��{0X�񶡬w��MM`��նƛ.^ɪYiؠ(��E�T�Ò�c���/ڛm;���V��j/1�dUJde�3��HPBb��R����;R�R�m:�p���ݹl�qx��h۫˫�4m��ӓq��奏K�腻t�e�eeǲ��Z� LͲ�K4�[�,���h�iZ7v-��1�.Aiڣ7≋
vn�N���5�ȕ��S�*�d82���#�яq����j�Z�����wD�¶���`�^%!P]ha��q�̻17��["��y{�w1�r�����q������%wq����N4s&1^m�{���g	���v��x-��I3�i-ז����E�8�)�U٫��xbg�F����8�b�A�ø&�ₒݘ�f���1 2��v�{�Jp$d
��Ad9nh\�V��#"���l����^��mj�{*Ev�Q&�=J�4{}�O��l}�T���]k��d��GLݍ���w�����f��X�<�B��[�v���o�[b0�ಌଛ��D%�I���Ro"�3rb�pmm�jf�7Z��)]۬6^��  W���r:��򶋌f�{�O�Qd��P'J�V)S2Ḽ����./om�Zy4���{�/k�$JY��aGpЂ��V�:U�T�&�ͨZkr�Zv�h;����9��r�^��[��3D^�ݰnP�·I�gUk94sp7�Uϴ�z������ܙ5b%5*[�k�(�ܛ�T�.�m��3�����lV+5'AL��֒�1���ȝÅ�2dsC��&�1\�Z����óu����pIn� א7V�<׀�=��76�X�4Mn���{��Y,����m.^�I$�C$+��16���2tC��r�saݽ���Ai��DM3*����eF0VT$�D�D�ɚ��!�otP�-�&���Ŷ7%9���I�Xg6�nL�¯lڽt�폄Ƥ�B�[���ۨ����)R"�1ް�익�w-d" �rT�~���8��l8~�F��)����i[��	���D	������8�-�[y�A7k�k+w�tT�����y��y�5�Q݀iS�s1�)e��JAn���㼗I��W ���̲�q��A��ʵgA7��{���\n��j���N�]��nl��9���@Q�KE'��ʸA�Z�f^��3I̢r1�f���ѶF���BqnjM-%��u�F7[dA����r�7��ӎޘ��K��;f��&��X��2��86^���V���xmI�-�V����n��{�E�f����xȑX��c�Jn���B�ۻ�li1j׺��0�n��{N�kok.����R4�v�1��)�U�H��#o�UR���M��%km�Pphm�Hl �͓J��k{���v�NY3��7�1�3o/0t@�nk�t�B�J���n���m�4�����m�0�ء��]�k|}��[b�N���J�4D�`�4��^�ܙ.���4�@c��HSA�^�,�R��H�7gh^�����-e�ݖMM[�Da��\3.�3Lޕ)T����4�ۮ�1�Ŭ�X�C�-D�5��d\��ǭ!�hTԝj{corؔ^�Y>$�;wB��` FE�B�V�Mܣ-F
B��Lj�.$
�肋v�
�F:�7�"i�D�N������I#̻�;2��u�HRoE1W���sB˻��Ӂ`�M+��hX���-��n�^c���q�M��յ�N��>m��>��hM�dږ3�h
B���6B6��V��:�S��	�6����l�7E���gk%�>����MV�e݁�7������]	I�AH!{p�[Xqِ�L����ͽ��hQ��Xa�YsM��ؖ`�Wr��$��k�JSt�囍L�	�P	�hR+a�r�����l�4�S�u	ycr�쥛>9�R��
�c6�f�r��d�dU�^����{�����R��wSi^"�J�ʙyX��/l���m�kc'(�v�f�y�ͺ�0���<]!��'w�y��&&�%�}�#����0@[t"N���QW*m�å�.�O������%I
�9�WQ��r�k��v-v�����
��6�̱M��UwW�6n�;��ہ5�I�t�Ii��5m�ѻ�zP̂����;Q�*ؾ.�T�,�b\��˙s^�N�J�¢˕�����p�u�͵��j���v�m��g�ar��D&��+��&D#qHͼ��52�����T�c�m��V��۬�Y7.�Y�e�f�®	����\�n���"ZV)��s]@����;�Y���2��r�2�.u�3i�L��,j�&�"���ʃFj.�]mX�c^��,�o���eYX�X�pT�T��q��7�f�[�5C�N�,+��*c��l��pl��3\ِП\���sj�;�%^)���f�-_,�t�l����+sj%LDb�ॷQ� �W�� �\�f�&HٵJ�0�QtgTC���%V��P���62�ۼ#)�1�s[�֖�w�3q�^�jok3r�J-�A���<80��U��8~{ DQ�c`8����!��B��R��ũ��'�16 ���̥Gk0�i�c]�P1��E:g^�!B��bb+�3z��l�4����ܚ�酽	���&��ۖN(��c6v��:�С�y`��=Ǧ��p�43�F�N*5n�@�+n�fKG9wY�M���Z��x�1y�1[�7)l�B��PnQ�g77U�DTp�;1�6T�͹�3;��7��TP�a���20^kR�nVh��N$�9`���Km�o���Ki$um�#Usa�T�����vdY�Na�ǎ�0Z9Q�4D^[3�c&U�����kow-ݽ��B���/oF`�3+f��ܺZݚ#0�y����cQ�`B�P܀n��K%����Pư�ŚH��!R�I�C�sh�у�/^�vb:��^�j���+�ɗ��k+@7�p�f�6�)����:^L��� ���Y+%P���ct�k ʻa�7����U�dz��,u��׏C�������4��v�b݋+/tIКK�TcfD��63mU�(��75��ٶ�������
u��r7{ be]m�d�L7��9Wm���i.����s����r�]�CD{
VocF�S0�Z�����5���ৡ�����0�,��3s+/&�GKrȺ@�F6����e��j�n��ƙ��n�Z4jP��e��̛�w����Ʉ6��SEk6S�
�'V�\ʴ�>�6�ukG5�كE�h�q"q��/b�h�@��Pp��Q�%��M9-�XJh��]�y/fF�U�esf5kkn,٤"鷓lfƝ��-(s�.Q�q��7w*��1�I��n���`�)k"�0nc�
x	st�[�B�F�蹵���c��Gץ]�e��K�4f��aM�ǘm��X��E}�Bъ]�_?�Ь澓>M�2�>9g�<��u�c���6^ΐ��xa�AW~.��3��i�r�S��J�$��X�; �*ؚh�2������f:жfӻ�%��vv<	V�!*Ͻ`�a��Օ%,��۲��3kt4Iy����%��.��{cqVg�@$��.oY�n����A�ʴ�sJ�ek�m�qj7�`cv�����&�5�ޫwF�3a)`4͑���;ǗF�D�m䇆.�	8j�0E�r��-
]�*��(�S�p�!�i"�LL^%VA��S:)^��������:M��w�V��^�����F� G��Ӣ���g1�b�^C�@�<-1�u�U�.�g�L.�X!��[M�zֵ%Hp����R�#��ޅ��a��^n�h��˕7C{���U)�ЈÆV���^f���r�#�hfB���,�NY_h��r�itidj��G�W��҆�M��(��ypZ�`���B�f�2�͡�
��nS{R��6�G]I䳋Md��EL3U��%&.�7��>��#K뚕-ܥ�6�/f�j��F�v����#:�^[I���u��s1 Y����V��z��BDΜ�(��V��%o�Ͷ�Yyx�h�0�a3[	���ɣ(VJhݬ��el�G�da�Ʉ�QNN�����(��,a�oU8�&
5�y���M��jd���)6�$��j���p�J�󘖹,];��s0�F2�3@�����h��*�

6;4)��d���G�ٚm��.�
Ȫ��;6�ܬj�+��	�����9�@��
�xVn�N,�Mն��²�J6RWB'l,����ȕv�(�/"r���!7���e+�wv&��U�M���	������r��uo(-�4��G用�Vk34�nͽ��R��,̬ۋ�Jژ*CB�b�-��so�Pm];Y���Iʘ���5�Pܲ �),ӗ%��L)�
�E�Vc;Wz����i

L��t�ar#R��[[(�@�$�M��İ]�9I\��Sl�j+֬��3Wzi;��~�BYi������NԼ2�+�A�Z��əDSvJK0;�1�Q�Kv���9.���tc�U���GF�:���2j����"��Ue�Sj�ݺ؆S�n��[�A�&��ޜ"�;G2�*tvPͱ�t�"���
�#�1tK���D[�ˠ��V�͹�A���)��F�!�y�3��l�����M�D2�V��hQŊe4�U`�46M�sj崪]ܷ�vF"��t*&�KF&n5��X34��׋N�eȍ�r��Uu f�U(�e���iښ��;�����Ӡ�wq�&#*s���!�p-������"ё5SAe���@�a
�6V���ج�S� �a5-�"��I��F9n�����	�%ՕGam�xE���W�ixV�Nm���K��Ƞ�n�n�rZ�4I�V���Q��+*��T�H�m-�77e�k`7��R�ź�H�2�܂�R`6^��cҴ��[}�泙�^^�eg�A1b��OU�I�5�(�6�PGd{��k4R�k&��%k/o6�4ٛ�VԱ2)�B"�,�FKL�trܡ��'p��	�&����Gs�ig�.�Z��wE���2�	 �������g2�$jdLKr�X��
|Po 	̚A������y8Y�R�������SdX��Y$R˽v�	S��y*CJ�76�Gj��"���O���f;��L���&;�uy�
�06\IY>pQ�hY����i�^��q�ۂi�G
���&�C�'2h�W���vmE��n���� K$�oDh�'tb��w�䵦�'�7��U,˄���Ux��q����eAoRkC�ˬ?�I[�d��%��D9j���Z0����`�d��N�JvVf�Æ�wi�{i�M%W��p*�b$і& -^���ٌJ2\ ���Q&,_�kj��&L����0�V7�T����(lb�"I��\C/u���j�aŭ�c1*�)X�enYzSrh+@:�R�6�㫬*��6��̧*ej���=�od��E�d�� �n�ܫS�(@I�c>�J�`YFl�M�;�BϮ��n�ږ����6nO��-���k^S���h	S h�f�b]�{/(E�W݊��`SN�L�� "�+�%�pP�K/�eL�Aa�96���4��}��4!�6�'�h�\�U4V^%v�9j���8+�m�kAB�Za��gkEP�٘�-�V�`�4e{u7]�X�qf:R��5�������(�J���%j�Z_�Y�ܢL���g2$�JL*�Z*�2�9.��6ɹ�l�q-$�����D�v٭l��
�ⷲ�ݝW��r���R���{�t��<D�
pX(Iw3u�z�kF���$bزV�7�y9��PYFa�46��7��f�+	I%Y�e:��&�t�)�U�6�X6SG-�F%z5G^d�E��ۣ��+w��RאC�b�*n��ʻ�k{ �����A�z5�V�)T�v]����'��j�V�ܽ�v�5���b��'A��0Tc
T�ɤZB��[6����i��Ui�0�`�::�����&���զ�B���Vr�,��'Fh�ؤ����s/>��-M�xn:k���J�l=��ۦ���c�9-�zb�"A&Im�um=�Vp���單��b�
���AX�cڱZΪ��z��7Ϊ^rw%բ�ήkxR�Ю����؛�XH�j�]1މH�q�n	�g.��	���ڃ��2EH �q\լ7J)fL�Xr�pn�ٻ6�������(��YA�Z���q�e�n`r�Ӹwa���p��;���9tekD���x팕y����ZۯWV���MAIT�(�vURr�ckp�v7��(l�6�K3[Mm�%�I�9���z�;I���N2����rݢ��p��U�[��vێ:3�k���Y��o�Elp�����lt�yl�5q��\vIfpGFF4
��:�f�tҋ	r��k��[Z�s-��g��S�i�O��哭�\q���C�/̴ՃetZK�\`���z�$[y��ˋ��2+�t��
��HXD�
����o9껵��t�vk^z�2ܻ��kX�������K,�%E[��&{^�x8j{��{ƞ��n�mێ�.N�w5��2�(�{;j(cΝ�n0L������dlՎ2m��6��u��^7Y��<@����۳g�dΝpSLQ8a@lk/��5Fh�9:�)BY�r����+�r�%!��xtS�P�Z][��c+��fu�
$��-v��]l��4t٪5����@%%�s�[.Q��kG9���]�b���`nL*�eu���u���b����O;�'����Y3���ʇ\C�p�z�Kg4�E�iX��y��u0�/f%�`���9�����u�/+��s��#X�K�6���:���=x<�3[nކ���vxct�8�����֞@����i��;n�2U5�Av�!;�a���)u�]6N��������Tۓ�Z6Ĳ����#pi-�HF�b5�N)}��9��g�&��K�#�;��6B+>��=)�^��8���چ� ô���:�8,�۴��]��<w;���N���%��\����JB+6�����$vis'k���W��vkV�]WT�9����u9婱�Qs(g�س�78�ǳ��(��.���\�����?8w�)���2��<�\N᫺�b0lǐ;z��v��X��MӲGm���X"�D?c�f�D����q,�3�_#�����AƱ��/�,�qX�c3۵$Ȝ���vNg�N��v��hM\����l���*�D,1(��KnR�ҵ�iYS%"�-[bְ�5l�M-kqc"Y�7s]��1���ֻ
���;�^4u0q�.�y���>����oo8B��i;y�pmy&�I�1�c\c����6cso#��bWc���hm�9�GM�c�.玆:�=��p�<�܅�������쮸a�8%�W���V�N#4b^������wV��:��8��q��aC�3��n4���� 1�P�U�8Iw3 ]�oR�ʹ�:h���m��H׋�l\g��v#�dX�'>KL����+Q��F�5wS���v,#���]@[J�n{궼�:���:Q�J��i�h�:�Lc��Rڛ�<�db�'8�{y��z{\l��l�K<�gy�U����Z�6;V��jI���&��QPX�"!h�Z���&a&�l(��ff�Zܐ4L[ST�0K��2�T�es-2�i.��dѺ��b�[t��cu�K�5��Q��Z�X1�VЗ\/;�G��Ä��Y7\�H��� ���j���;F�_GQv83�nI:� ��< �����t`��O���S�s��A�9)'�1&��4�toXZ�%��"3���C�v��GS��k�H�mɠ� �Sf�Up"䵎�m�tԛK�;m�����C��� W��9 yU=��M��/A�K���v]Rd/h�4k��LX;,S�.ˎ���+�$|z[J9��B����s������!���)c:�v�+Q{�3�W����<�T���izx���{P]nݮ���]�n�1p��ƹsڴ�<ɹ����;�L6�w��Ge���M��{c��.�S1���ێ�X��8��lmAr��ܣ���V�v�N�(.�n�&�lq��%��\�	/W���'�D��by��1����!��^M��q�OU^l�v0mp����+������z;/�g�-���V�a�2��8`:漤R�Q �֥�]�ue��7n����{w4\�9v�R���1Sa䵌��؂G-�8yɭ�J�+���&�����8�8�n^RN�yå�A��v���u��0�ӷR{��c�m��|3!�dy;\.S��p�XLGd끷���rF&�cR�Vfm���""��A�b�s׎�\�[�#�ٽ�L��<����0vLq�ݷp�mPnj\��y��n����x��)�MIE\�vҍZ��6ƼE% 靽`�����ۮ-���&�:�u۳髗�-`�r��$ɸ�8͵���z��1��9���t�������]K�i]�Ȝ�]i�G	&��Rm���=g��Nwd��8��۰��;`-n�]%�4U�F�L�ѵlt��Gs[���`�㫓g����)�$4�%"�ܷ�4U�,�+��*6Î��FM��/���29�㭩�7ku\�h�̛��;����c�.:��QwX0�&�,ɬ� %5�:̳+�l�h�4ȥ���u���G0Q)�u\�b�iM�v���$��9�YN8'��r�O'n�U^��TM�iP:6
�!4�v�s�V�Xa͙����햁�P9{=�(���$����kc*�ѹ�,D�d��BZ��GX�U�i��Hf�p�#H��js`��l=1��҆9s�g�ۺ�=����.\ƺin��۵��$"�6�<mf��Q�'�%e���k� �p��g��K5h�3՗���Z��F(`�Y�K�:�E�;�m����-�Y���2o ��ٮ���q�u�,s�<ًc�
��w8:L�k4�M��B���l��!�O<Ѻ:�0�k5�\��f��:YL�A��\ɐ�`\RMc�\�0� ����;t��Y�a�j�@�ѩlъ6�*[kZ�3\kl�q�7a,t���S���ϋֈc�l��nW�e<n��:4�μI�We��ǯ���.�JV;J���ԭX���v8�)S�/�iT�x�F�P�i7+��ù�E� a=��>��fc����v�'�����˹��N4<oe�$޻g�'k���U��b������,�e�	WZ��s�9��h{BmZ�\ø�0��8/Y��ӭtODen�LӰ�v� �yU�q��nn�����`�[����hX+I�*�g8ܯ��5����''Q`Yt �ٺ�5v4��ΫTf�*��_X7��$���#m,�����\��w��>i5�=mI�!����5&���^�"�,O��c�
�n@@��X�#�g:]��4kb*��sv�2l��ZZ��f��s��*P�*�y�x�\���吨�9�tfX�Y{�ֲ��­�dřI��XpFZf��гe^�x۴�v�v��]�^1�ݵ�''�IsRá�����=#v�k@���c����O��#p\�6݄�Q�D:Zxɺ�c�	�V��iJk4�e�"�&4�k��� ԷlLHh��e���km��q����z8�u����݈�;�7�Q�
�9ª:;�g�	�҅ט+�l0��[
g��	[թ\ʅ��m5� ��)��e|�̠[n���%i����<B�ǋ/.s�9�.G��ynަ���z�(ɶ��&-��z]�W���S��X�z�aJ�X�J�6Z!6kuV�&�^i��#@�Q7:ڎۆ�]:�m�^���e9�E됍���G3��z��G)!zs�h3�ۘ��Z�1�-���t�]��!�k{Vh@%ͻ�,n��4�m2�n�{x�3^σ]io=c��J/Vu�>�ϵ��L���N�N�Abm��6��[��f"�s�n���.�[�0/m�3g��W�9�^����7*]���Y����XE��u�O����J�K��WJ�:�0�/�v܏�-�:�E�6��Ofe�����Q5�L�G3iq*)�6��C��wb�}\zSj0Kv,�	gb;!�7d"�t'u�/��W8��f�,����8��0��/0a�nk]�ҚL��p��m^Ggi� kӴ��Ud���O ���$�ą���\��ܬ��m�lɮvq�\�^SǶ�u�<���A�2��������[2\�&4ի��p9jD�	�]t�2i\�����j��� �%�g��P���wpwj9�ٕ�����\�Z9֍lsj��l�3�ՊI�ك�/e*�n�&[L�o�s`�H�G�e����SXgp{���;o)��=��O3���Wv��:z���{���䡌6rm���p��s��4��^̶�:��ԝ��3�9�uìM���3V꽊J��mi�z�I��]�n&m:�8�/(ny.�刧�'�����jy��E�R���Ѵ�&�n#{!�v���;ѻN��y�>@��QN�-���S8Bm�Զ�J�]dC)ó�L\�y��E-HlG��A�C�ӄ���ܲ=[k�4Z�]t�խP�)lV�j��[[ �!�q�ܛ�)�U�8˷4�n�9�:�]tm�C�&�C�5'v�k��>�8<!��Ҡ���cHs�ۗ��L����k�s�ϕ�1l���{v�9إ��, ۤ ��^ޏX^I��e��օwg�5����g]��d�g]s��K��٠�Ƥuf��]�I����U.}�1�Ó���*]���]�=�nmܲKvlmO�� ������0Gp��=���S�g.r�ŋ� h����N� ���R<�CBEѢ\̇X�i�K	�Tsm΋U�{�q��ӷ��	�q͸9�}��h��cH�a��GB������:m�X���єq'��v>Ŏ.Ri{n$ݭ�K�)���渮�â��`y��>��Y��W]stsTҲ�l.g%��U+��P�m��Q��1��fj��i�y���Qq�-�-��-���eS\�ؙ��w8�r�dU�8ܭ�{i��g#�փںU�s��s5�����ݻ�S&{s'c��ٚ}aM�5
�O���Z�s� ޹��E��)�=���M���kx8�n��ܜ��.�;�q׷=(��l�S`�l��(��	«,����K3f�Y��f,����k3?	f$�f�fbY��0X�f%����܃qRX�`� ں�Km����7`�<b��Q��w���\�s9���u�� DnZ5�]��ӡխ��Q..�0-G�K��M�t�t�!p��w@6�l�*���y�i�+��5Z�4�E҉X8L@#{]g�nG�.}�a�wX'q{.�r��L��8���&Z���h�n�Ù�6u���Eei5$m���s�آ�I�׎�cnQ4��/.
w:�m㳚��+��g���i���qb�&@�2�#K�-ͫ�WM���.�j�^
���%e�m�a"������v)ڰ�PY�3�Ŷ��ˠ2�����&#Gc�<�s��r4I�1�\:S3v�<�]���=�����X1ۄ3�ո�z7�6�gt���Dlx֠�騥 �2��6Je0+�^)�.��Е �$�Ѹv�L:�&�W�*nNpp��,{wF��p�r�����6GD�8ʎ�2�����In1{u��Rs33-i�"�7d��6I�V2�mq͊�q����#b��43���bG��;��v�4�P����%"
�����v���IjIM1��]Xs��.�e�l�����3H�2�mɥ."& X̱�Fݘ��؝��b�v�e�|�^��F˰6�������
7dI�l3I��7<F5���-j�aX��,���Uz�m9��"<�5�&�iy�����6w��磮�}����N�z�v^-�ѭ�����k[��,�6����"s���碽�[���n�O����9�mֵ�^N�4�����\�<�X�t����u+F91�oS������!�W�m�r�c���h���p=�u�aU���.�6����8lk�`�c���K����ؒ�v��#�+Z�c�9�F$�s�g�:pv�ȯ���N�y�/<�%笓f��.��Zi6!5�˖ˢ9.�����3K����Ԣ��#-�h®�lЦ!OU����U��ܝ7gG	\zX�33_�Ė`b�İ1f$�1b�A�bH1b��X��X�b��ř�bă,�K3A���f$�,�ĳ$�%��3Y�	fb̋B�ݖ��@��p�^���6F��[MY�֤��L�P��a��Dζ��%����d�m[�Q`�0��O��0N.\R�WS�;z�Ņ��p���S����l�mj;�y��ax�L#�IHݪ�6&1�Ԯ^���i����s5Bz�ᰀ��e1���d��a������+�n�T���eclŷD
����\>����=�-rt�tOu�<��$�O
��pq8���j'�Kl��ٟ�qR�OO���"�$9��f�Qe�����ȼ�f4��������qqL�(C�	8!&`,rJ{�hb����5�1�{u�ox�-K^,�ao�P�Hw�n,���-:��I�ywB�����HA��-��j� �1Qq��]���UK藗廏\;�0Ъ��jؐDZG��z�}Xğ��}��
�͚������H�5�,z�v�W�J�屺�� ��
Շ;��� ��o��L�Pj͉�Ӫ�
D�l#0YA6ڒ���c��^@�W�SINY��)ץ��
��<N߻�~(��s�Or��5�����qh��h�Q��9��A�}�ΐ�6�;q'$����Bv;�A��iS�Ã��K�,-��?��o�7|���|�#�ϻ4e��O���J�T���E�e�u�Q� �A��k�b��Rf|�!1�bS�-M�8�:���V ���o�:2�7)e>:�nna��β�n\�E�*]���耈Ƭ���ߣ���5�6�C���Z���L��b�&�V'"a��JhR�t!�D�wtQ�75�L\(�F�8�o:���)}�r�F%n:�Y�15y.o�z*%g��r�@кzӦ���n�kjc���@q��M�B��]}�}*v�����7��Y�$߯��b�������hp}�!z݊�*lq!P�:h%	�m�0�� ��Ϳ��d>-�q�CK��<�2		d����&����ݥ�tbf�ڷ�m�IG�lE�t�=�F�v	p�B�G�	\ݴ�&fb�K�0��F�*İ�.z�d&A�D4�k*7Z��{χ������ M+ۗ�f�Ŋ|Ld��i1il�y2<�Γ�D
��F��	A�Cg�dWv��Ok���&ȁC�Z�̠�TN�H�ڐVPg�����M�a�[0�S�����D�A���-��Rϲ���L�"�m��y Ջ<[�<����<*�l9�7�]�50x��7oW1�K��yM>�"W]q��"���.��:��HA�5��y��>H7h���;7%�ĳ�����T�94���Nͽ��Q;\q;.:��]>dw_NV�Y6㧌ې-�d�PrJ�ƴ�� �i�Ub{.�`6rQɇTj3t	�*jc��ͧ%n:�+2;V��GY+�O\ir��Y'�n�"�*ά#��-����/_)[�� 5��c���o3}��ش��eclDĆ4�j\*h�r9�^�6m�mƽ#k�$�.,��F�i�w|�HKHQ*��j�`�roVש�!&�ޞ�P�]�2��r�:��*F���(�t���-0�M���M�����Uz^�����5�����3T�M�ϟe؈+w!�b[8=�y��7�+�v_oK�iBh�!e��Dq���Ƀ���ԑv�Q�8i�J��smS>������O�ϑ�2�M3a2R�ⶎ�i��Kg:������ovE��Sv�}ى����p���#�;v�폺�(�;�x��V�uj�!wsbW�ea=C��$k���N������ |�^�Zz��o��Gm恴���X�$�sP�,ݤ&bۏ����DS�i�M�X�:w�KRa̪���>ɚ����ϙ�b��2o��&�v/Yk���s�[�Da��/�s�5�d��e�5Y�i�������yy�K�kxۧ�
q���a}���1�m&�
��i��)A}��˲5ó��`�=����0�B��e�0!���]と�ʬ���e�n�o�ܪ;P-� R޵����_�Ȧ���W�Zt�a����ܫ�c�ۙwl��c%Zڛu;u�d�`"��E`e���P�*�����o�'�G��ٮ��*7.���al!t��^��ƢK��ϟ5����L�s�.���֞�����v��v��z��k�/�wی�L��v1(���p�3e��d����u�TL��z��8� � W%\#������ퟍ﯏xm@7܎+�H:�I�J��O:�toE�,`�N_l�|���
��\hv�yj�v���n�(%��g����0��i��$.�O���0�鑙�.�*����hn�5�Pr���3fqN�ZsI�njv�;f*�K ���
�EplMmJ�T�B�,��c��`:,c��7������5��݅�B���]a,���Όl�j=�M���L�۫mK
&F4{���b�L�ݯ��L_�Al-�"���G����%��)Woe���n�sٯl�q��y��L1����*K�S�W�ò�3gӛ���+"�;��W�c������k��wk���6.P'�.��y�C�d$��n��kC+=�iz:q���j�vI.]Fr�Ff�ͦ��>�����@ ����-��ݕ����[�$��/edL��U$�R�}�e����d�a8,�RbZh3���݅�H�75z�:̑Xv�J���+�z��D ��ߌ�Y�W��8��kX/-��n5cl��fNT������>q'G�$�n�ƹz^
v�]ec��Y�(��a��M�o�ͯuU��ƙ�y2Ƣv�9� Uȃ�5���yR���to���9)?A�ʝP�  h��e,u��T�=lζ�۫�~[+Dq�l�KV��c��Q�P�X�3Ժ��EKZ^I���.6��B���`əR$B�|����y�k���l;�oj�RLt@un9��vv�^qs�l�hؚ$��m[�v�
�'aɎVY#mڣ��ވ.'޿m溜��^m�x0���{O/?O�U�*�p&�\�R(�۔����ɶ۪��4h}h���}99�湠���*8\d��AR���y���A���9n�X�*�nS ��u��#Y��v�+�T1|0euV;�dj8�	˭¸[����"�bVͩ$�Ʀ���F�d�ى"o���Ͽ�)w��7���"�!�<�C��N��B)B0㶺Ń#k��á9�T4�Pz'��7��9��,.�[B[�x�Bz�9
Tܫ���u��1De��Q�3[��㩵+��v,��"'ʇO�p`���ϱ.���붧�jf���ۭ��*#*t,�j6���{	�Z�n��1�aU�Y���"p�M&�b��*�q�8���Vު
�|rPӞx(�B"��u�6Х0����
Xx�4��l�NQ,�+홅,;6��s-� n��)���`�����ԗG# ���h���U�pX�����z�C�֪�����}FP������s��y�ub��Fj��k5��ֱQ��H�T��ⲵ>��r<R+���B1D���[m�\i�c��e&&�
L�׆`�s^wWL]J���i��u�(�j��9a�����n����0��U��Zw]�/vlx����ݚ��h��0�|��9��������J�l5���+2X��GuUP��� �t�"�&�$�)3�&�e@)U�d�2�����	�ܕ����/k�q5 ��H�{�7��b���Qw��1�xU�6�m�%޴�"sվ!V+l]z�s����U�^�"1����O���ws@��^Oy�$Lȇ&o�kZ��p!�Uy׿^����j�HHΣ�������X�y��:S�p�\��w�7�]e�O6٣��\lb�?O�!l��>D�z�?�Cvz�i��%2!��d���+�7Jy��TI�T�ޤMH�YO&�TKK��l͆6�'����䞳�Zf�m�	�5�(q:P�4�re�8�����1���'�h�g�/���ܧ��o/쾸���,'�6��Õ4�u3�3�� ��ǔ�ʒ���[�'p^�$lh�Z��t�,���O����}��}�g�L ���~�����Fs3��sy8:t�����٧�VN@~������:Av��AbΑ8*��#kE^�ـLP��N�[��a�,,�}�Z84���N�jξ	���`���MYNe�o'-o:���C5laUĕy���
�E	��T-�o|o�C���w꩚9���1��`��3��qhs���s��x�*���Q�U\�զ���IM�������X�П��k3�[f��/m+T*��b�.��jGT�P�.܁�t���)��M�t�J.4�5��F�>N7e ��Y�,�b�r�	�$�+�S`��]���0x��7t^�V����h�0˅m�̊m5k{"&�驕/Y�2��&Vޭ�!FKS,��duE��[�3��"����l��PBeJ�",ϟ�A�4R`��BUUȮ�ܫ�hc�9�~��$T�Uي�l��0xvEP&�����J\fړ�YAX&� 	�l�Ö	�+�F�9a�E�`a�W�p�H�,2'gn$ç�}�2��Evؕg/M�:���g9u�?����ߑJC:���1�����X��0��(O��t�4�g;�%n�2�X�;��Gj����Y�S�O���ȀGU�Un$�Z��[���������� YV\�{��B��r��_+�얪�}}�`8�-���!A,��+F�]�𙹜�T���t���%e�����%�`�i^Hm�[�<#s;����l�U"�J�O s�C����I��v�e�N˓�l�;"�I"���G)�۱�d�KP� 8BD�.���p4_��;�4�F�L�bT�4ɣ���:ْ��gEG�zض1�%]���z�{k�Y�`�^�w!�]��4Ά����Qa�wR;���͘e]3f��:m������ �+,M,�vf�.n�&sp:6,�����&�n1Ӓ[��m��-��$GeRL�"�-����kLi���=7�L��=7��.NJbi�_W�C��EKڙ�{��ř���:T�y��*p�5#ރ	�6RL�˳v�XTd��)p桂�ałH�j_t��þ��̿��s����;�u��B�]#�A�ac�l� �>`A�m��� ��|�֥�@3}�km�������cƟ�Rf15�p�	��˭��w���p�c�n���(���S�_���'�W�Ul�FnA�gOk���@DPCφ73<�+�m�"딫�<[t�!�Ÿl$��h����pB��L^MÇ/���<�2�Rk�N��r�
�]���U�ǝL�6�(��}����JF��j�9���}���z������
��P�$�+���4uwk	��%�-J���Olsh�a+���-D&WEl3�,J�;|���]0.8��8��WPٗ�Ϯ�i�رY�hWn��!����ee���06���S:PB�B!F�Rb�a�I��1�l�/�~V�����7�]56�<�M�Fݐ�D횻0�Y-d	#<�X'[�˕�y����E����X�</^)��x�PK9���K�([BfHZV�d�Lg���Z���9s�s%)m��aCi�Cm�.$��tun���޿����Ҳ6�*���y��C�m剹Y�4`�H�ݱ�ެ|��6��������Ha�]����;)Ƞ-���,�{��s���:�'Kj��
J�
�w#�|�<�9�4��[��L&	���IE�擈m<�t���"nyTc�
�6�$w��*V���W��\{.���e��@����j˹��v.8ۓ�J��(%����~�C�\��I�1Je�v#�5��c)qg��́��|���ڷ2x]����M]�ɘ m�h�x�P��X��Ӥܷs&"+s�݅ke>
���*�=�=��?&��.B9]��ߤ�b����c/�2�2"���۪&�$���5ܥP�#��l�[.��U3�q?^'��q��U��܁-u�����bۃZӀ�7���3Ah%�����}v�*5�A���;vY,��a���k�Wu�����0����<8tH>��e�2��'8��2�TkGv�-s�Tj�Pp�����r�͚��1��̮�k��Uk������ı�d�EFj5��f�b��{�^��%��Ս�V�����q>��������Ft�,��X�㬹N,�޽s`nP�~�b���Ś��$!1KU�����8�r����2�cT�=l�38�K����։�M�Ȳ��9ՙ[A0������/k��ê��0�GR�*�A��0������"�l���4���͓s*U��J���}[2�&��W]�\����>��8a�r��3�]�B��
�n����=�붩�0L�&Z6����]{�fs:���� �oo�C��pW��h�{kL��Mn��R�M���1��"�b���DkPB�{�1n2����p����N,�BۚW)���ޱ��3%��nV��p>tȜ腐�If�r���K��ݽse�Vf�L��>���c;�R���5a�QΫ�n��1x8Tc�+�c�nl: ����ﭼo��wW-�Ǚ�sFvT�s׭\]����V���l]hQC����K��,�V���T�Ŷ-.����Y{��oi���%��(���t���p��u������+Mؐ��OZ��-�2�^�c�e��܍�z��8�g�'}8m��-o0_U�K�y��U�Ń��u�Olh��'uh�N�����\E8�n��NP}z�R��F�y�t�S����sm��M��C�'M��<�9��uY�W�u�/�r��"�a�XE��c1#��5�XJ����Z�6����4�1U�Z�5�ɯ|�e�{�V�A��粛��������a���&P ���)E��v`�;u��L++��L�W��[�jS���6�+���x�Wy��e�g��,�����v�ݡ��taGy�Q��2�0H�IF�:�vT�8{n����&lN�"3����X���:e<�z,]�ok��(��[�wۺ���m�1��3�c)�OX��3G��[2�iDm���t�+6B�L.STݗZלg�H*L� ��ȗ��s{Y&�G���;=�)����ư)l���T���0�-����p*�{���N�]*�o�۝YHq;6��5j��F��k~�֍46��:�i3<JF�b����0D�uB7�5�B����P������9��CQ�C����;���o�x���`�����A���y���T1 5��aA�m2�A�F:'(<�n�@Z�s��lU�x�v�r�&�WSOCy��B��|6_T����!�T1Cm�v����7���Z%Z�0��E���W-LFawqz"j�/،2P1�fש*c�*��~Ͻ�=�;;۫�5Р��Ս����Z�1R�RYY8H�!�����YaP(�a ֳ	�o"�;�Ç<�d�bM���9���,s"�O��u}L�z��q�;m��:ݰ��:"�pE�:����[U8��;�"#'	�m�j��w�f� �<��6�`��*̅Q���>�j1`��bd4Gaw�v�c�i�?��zY��fM)+��],;��X
��S[���BmCq�ڭ=T�dWE�T�]��8,� E��I6&a���oK�o��foZ�$q�5<�wi�C�����^F��u�Y+eģP�N
�s���V�AM���b_�x�)g&�j ��Z��r@��R!%�~>�EJ$�s��_�k(e�K�T����m���[h�S
m��Z��,)i���B65nN����O�ʻw{�4������|61���s�j�(bl��g��M�*%Y[-҂Ѹ2�����y��%*��ЏS������~w�^Ӣv��6�ZQ
K
��,R����Ytr�[�Цj�k�f����>�cb2!qM�JgE�&�1���.{�z;g�=�qi��n�ۢ�7J��['$=��4܅�etQa	Y�ל�Xk�Iv�4`�z���*u�:̈́�޲qt*e6��s��9l�j❠��w������S�e���6�p�|��s�I�q(h2�-�ؽ�.>?15�5�:�h�is
y7�n6�%P�S����Y6)��x.Z���x�J�>J�[:f]�cU�p��Zs}�*�CQ���;�G���h�HD;{.���F������Yu��$vf�X:�P,��%m�ڻ�>5��'�����2z�:\6�{V�f�7�d��Y�,�ӱ��4N_u�����lg��{�J�Wq�C�<s3*�$e�`j(��)r�j�����������=m{�E�.��4�D_vlC#Ne��-#��M{o�*�%�m���r�b�A�	]�#�Lɬh�eC��E���Wj�h33r��nu�Y&[��SǼU]�ƚƯ��4LXDV��oe�>��<t+.���74��3u�C+�F᪒ˁ^�+%%[��Q�̻�j�V��\ݤ�P���-�xd���wcr�X�}Մ޻r���!*�Yfh�蚦�o�g�n	��Ը؀q5��*bl9t�(lW���{���.(�E�����G�a��(^�:�w1]��1۸��og0)<Er�{��K~��sV���St93B�1uZ�+��j��>i�@�Vc����Na�c`�S�7��A�vh��1B�n;Tq���k�v����l�pN��V���3�B)����������t��'�Gu�Lu���ֺ�1���-�Ӌ��%�r�d��ߑ9��j��Mp�P�"�i�ډ���r�DѮ����Hf1C�K�!�$�H��]*�2a5���F���]��r}�&�"u]�1��m��0�D@�G�{��2\�9����0�����n��Bm��4ѕ��e瀥�gf�b��Fj�-L.�-�4[���h(�j�"j$襼Q�v�\��g�	�J[��V/m��q���4i����FT�S.�[GQ���E�nY�GB�D�F
��5V���e	]B�2u�QS�X0�f���2�-�Z��qY��i�g����<{U�
���M�-�8��\�д��]�=����[��j�t�+��;��zy�c-�����U{�2�-��hl�����ڽ�$�������A��G�3��ڹ*�h�͏>�ַq۶�������w�ñ��p���. �k2��g	א�F�ׄ9���ז��u�6����Uj�����!�̦2Bf�NV�X�1����E?&ۨ�n��6��ђ���9[��a�bz)��Յ�[Ȟ�W��m��))�k{=��YnB��1�2-ȱ+a���͚d��5Ca�`��nZ,��K��X�nikT��9��F�2Y���S��ffufr�U�4�3�8��~���:u�Ƨ�g�W�~�K�[؞^Z�G�p�g�3Y�2�8r�4%$�2y�f%����Y��uR[=��o"���
&#�&�x�6�!4���z}N�S<�S� �<}.LÈF&�
0D\�ȉ��$3�Qs܇M�[��&Lrqw�E���-*l���]�FU���?�a��?�я$6ZF5y�%`O-^�ܭS�S��	�}�]�Ԟ�mzhj�<�Sr�k&�<̭�O��X�1�'���ۗ��j����׍b��:nQT$h#+S��z/'�UQ�ń�]6��E�v0,�N��ؙ;���:{��{	��H�� �(�R"!8��	�'�jTW^T�2g��u�L���n�xn��Xw]
�
�5���TG�
����=3���o|���?����� ٗR��	��Y�63�a��_v>x$;�GMR�X̦�f`��nFa�b�r���l���ńb�uv���h�c�o�w�=���7��.���]��0�	��A=<cS�KM��ݯ\�3�U���ߘѢ��H��$\*�fN��C�U�S茷�j�a�ם*��s�8����{���XE�ܟd�b('m��i9t�i�L�g�tv=�]����0����l�Y|Ǌ���1V���&}�s3%����y�eEq��#�ٽŧ������3z!冦zv�Q�	+�ڷf��q��eԾ}���OWA�sN�^��>~k��1t`���y=����^����Xk33q]?S������c�MQ�����}b��'D�Xm�DSKqi�C�̲3��t�/�f� �ȠK�ٕ*i-����������c���+s$�.�6,�+V_��T��z��0Cw)�Z�ጡRd:R�wtл�r��KZ2�9tM��씑�����Fm�C�d.KJR��ͮZi�h��,��lܠ�C7��۳`��uI��.
��i����,cg�����׵���"i-��\��t<u��c��f۠W���k�[=x6��)�i9ظ�m�g�^X�6����M�&my�v�й�QP�葎�:��Ǡ�7����O!�M\��N	큍�(��.��>'<u+s��˝�u��Xs���pu@3���de6M,H퍆�f�e,�3��|�@���ϯ�U�y߿o��]��U�m��K��fvme%�y��|g.Ӫ	%��D�o��n!��l�N��%�̇�y8T�lQ$i�*��u�iV'�
�fsr��#4q�0�R�5�٫bntP�l��6Lm��Q�3wg&w��uM����F�(ȓ]u�p@�8�Nqz#;������5�7�|��kܓڰ\�l�µ=��dq����%-ӓ#&��{��0ei�ҟcvn���6�=����8���}>n�.�#�fy՝k��.oV��������bvQ��q� �%B�o��y@�˩f�F��{�A^��	,o��S.��̮^8�,�_����'�y�I���U�J輿�����j� ��l5������+�8���Ogk�J�H�je���b:��Ahң���<>=��N�l�%FZ��%�`�?kIf���a�����Ɯ@�C�e.��0�' ��(	�d��h��Ϥ��[����������s�G�EcY9K��"+���?u(ʃr��h)r�=�[�󝵳v��̘��^#[��S�
Wb����#Sv�w��ZY��p���Zw��s�i!t�e����Ǚ(�kȁ�*c�1�yg�ٙ�0�
<qKv�w�ϿHrP�Eaj㎥�UekHA9DrקU��zP������������@�sr��چ�;�P� Dm�BnS<��<���)����^7v�:Kl�dD��P�xj!�yǪ��a�4���P�F��x�z��c��5��#���YOr����N@5)n�7����6<����+iH��,QS�n{f�#\�(H��2a�\AԿE�7�,7�e�<�v�ݮNzKRmQ[[��\�7���Qu����d���]>O�f�#&��U���D-n(��T,�;�[Z۽�'����J��?Wϧ���I�>ﶆ��-¸�F��_�����S�,��ǫ`:���$w|&��^�	b���[B�":0�<vh�"N7-�%��l�;�j�X��P������ƦzeN�Y��� n�VmeFo�G<�F��,�Ei�ʼ5�s���2���!Ŏ��cPeڊ(aN]5WAt�"�M��B��x�\��eY&��w[�Z�Õb�d#" ��a�[;���+mu�9ԌZ%�p�-���\t�r�3!Tk��T~�>;�����L��w�5�ʌ{�n+���=H�h<�2���̴�W�(B�9��Q�[0��N,e${� ����8�3	1���{��2Q���YgBҕE,)[�����!�£Mt�(0�
��.�sp��r=tn\cr*�v�]���]�`*-{E�ź[2�@Wj���۟�O'�v&�.��`6���F[,���~ӽ4�R���'R��m ����V�;�o�RS�������ܳ�ކD3�a�!OQJ�G�ac��+6n�rvr�������Fk�e���ԮV��r�'_Gy��[d	��B�A����^���͝.��0LA�Ǧ-����!wɢ�ER�l3m�J.�TL���0�z�CF!0�)�6�j!�t=��c�|ۺъ� _.@hڵ2��{1z���2��{϶��]lG�n���R�X�gx�M��s��u�In��d7B{��(9��P�Q����2S���Znh�¶��-���!ܲ]\!B"L�wOK6fnYR����>Q /�>fԟG*��p�L�W��[L�T���'��E6�`�E+�����x��eV��#�K�>�M�vp=��(d���O���8��JDu-��IE�T#���V�O}J���k�����ڙ�t�Ip�u-;1�&oFz�S#��}�+7��A>zO�}��X����d��F3�k�/Z�w���2%����#��a�fw&b=�x�<]��4�w'Y��E�xk&�=$���ơB:5E����yS��T���az�S �3�����j{ �˻\m9�]m�p/�dj��껎U���P��4�K��Ja8�y�l�-�E��#fO
��U���d��T����=b�*`��)�Sѥx�=N�t��x�Pl���f
L��j�����p��!�?^}Y����^�k9�ـZ�=�M�hȗ�PN����.�k�,j�Uq���ޝw��[��|�� ΰo��H��c���n���&�w��r���l�8��P��K�4�W�s^mof���mԬ��Ivx8.�Y�ز3a�N�U
�
�'�k1�W�]j+Y!����*��{vH\�K]r��f�g^�w]]x�.����n,=E0bF�/~��]z�OR������F�#61�ەF��RJS���	�3�3sz 8��cpnS�	�&�۱uu�5��n��cUv�;FIR�na	>�2��f?��D���o�fI�]��ô�#%�>a�#��Fl=���E;�v`�@��o��{Ӧ��}����V�𾇄{[��'��7���0����	�[T�f/�7N�]`�Z[r+��+�t�=�A%X�{CN�b�@ƫ�S�P���{�v"���+Ȑ��S&�x�N���b�=md�ºv(���i�E����<�[�ffgt>&}��p���;�rRރ�Ws������jE�mA���y8Vt��F5o�6m��s���y 0�1�R��k�Ȥ��+d{�J��jAK���yC���K'-��q���J�8}3+�����:���?=z���)w-��₻&�c�β���fXv��Lۄ\�n�gc�m�NK+�!z���L���nA�A���ҽ��4�
���õ�ĺ�N��Kx�����U̳:&N��)��5!Y�{��qu��%����2�;���w#���le����t3aVZ΋U�2�j��+F���V4d�	hi��TLF1�%ZW��7f�
ۤ��3jKtJ��X35	����#��m���� 0]���n���N�V�-�k�^ю-���4�+6!X隂��ΰu�.4�k31�rZ��uup�3�љA����a��?s}�C������3ga�E�QװA�;v:����V���j>ޒE5���a�kY��\h�wp[�va���u�ڎ�8�V�=yMk��Z{=�I���'s՚ѻzk�m�������.�!��M���\dKr���3��0g<n2����d�͞�j[d�7�kL�L�����i��렭���/����m�fa����k����n�Dh��۳�,���ݫ�Ǝ�^$x��a�SĜ�rr����g���t�έ��2�1uٸ��l�)M�\�>�q���n:��u�g6>�\N˥�d��z�tvpv��ۭ\�p[�&�܇lmT����b����4�[�z�e�57g$�Q!�ڟݩ�v灭��֣t��qԦ��K��ִ�#Κ�Ŏ��&݃n��̽n8#wf�6N�Ɋ�WT�-*�4!Uju�Ml�s^!n�� ���r/-��D�[�Ds�O$mԇEĤsS�͍��;m=�����sZN�6���CN�t�粼Gn��Cc�ݞ��d�d�is+���{�v�]���)،��c���\,�Y:Fr�unى��J�&�e�LkaH9����M�rh\�n�yx�V������z���P���ˍP����;]cvo���0��MH�\����o�I�V�Ǵ�.x� ���ug�:����=g�:*��n83����k��tݨN����ٰZ���ݹ�u��-�y`������i���9kiKqm��m�L���bD�>�af���SZc���Jn�nK$����]�7�3�
�E�؆6٨�hQ6[��d$]㞗]�9*�Ց����rYm�U,)��D;n5�m����i�酦��u�w`wD��K�)h��Mi	j;"Bde��E�q��6��54�X�f휼�q��ݸ�c`�ܫ�#L�����&��f�^�=�p)d��8:I�܆7VP�UQD8G�Z�jZ�k\LEQ&��H���[N��v�6�f���#���r��f&6Uֆ���M��N��|`�p����C�ꌋ9�]EĻ:�N�Վ�jC0����]4mL3BM�X�!k��*q�[��Dڍ��8�i�}����	�K�~���EEBZ�"v+�4�8�2�]�.�[�S=��� �,����ڛ��UM�
�8���hL�0Zji���-�[�t�*�uF�Ɩԕ���kph�p���~�5�IcV|?�a�gBҳ�u�>�_��l�0T8p�0�^讬7qWKV�ɮ���S�m�R>��~�x���#����ι���*���^�՝ۏ�|���?��O"V�A���dp������ۻޓB�V�*���U����zrǢ�{	�#ND�:]ڵ��l3�<���p��(A�qrN����
&�:�a�CW͵y���P�Pyx�0�xv��� =e��U�T&Қ�^M�J!A��K���ݬM�8��	�k��q+u`H���Ŝ�=<nƃ����ٴ�b]�7�g�<����B"����Ym8oq��ywz��H�VK�zZ�^�G`dUIΚ�}]{�S�W�]~�j�!��'�
M���wHfF�]������c��̖���������T��ʎܣ� %�u�τ·.�� �x윯Fc�nt�pŘ�R���ٝ���K���sU�(Հ��0�՗r����_y�St�]5���a�wRfo��Q�r����d��X�R�Ie��#�Q��������41e���{p&h�j��"O8��th@<K)^P�;���Ma���I	��$
e4л��7��w��Td�ڹ�̗�2m��=Q{S��lc���eH-�H�_<�O�9ՑD��4���}���V��3Y�����efm��Xݼ� <���de�k,�{Ċ89��DS/P��f��y�^;�l�tS��y�L�ё�j�AF҅��V�
��f�#M, *��w.|m���n�[ �8	��)3t�5wr�^�X�)��C�	]�J��S�BE���*n��dK��q�r�ג����o��!C�X%ڻ��ۘݮRN����M�yo3r������6�P���� ʄ"��m!w��s�؎����<�h�C╦Ԗ
G-�wZ�H��`T��]S�>r�\�.�t�UQn9��C~����hg>m_s��q��Q0G�Į��9���봧�+f!:��݅���QV���;D��M��n�sv�
���w�7z�L�^>���݇yȫ\��}�r�8}c�������5=F�z�mY�S9v_-Y�y�|��r�V,Pt5%��kL$ ��3�&2d�SsEɵd&o������QKS����9je�]���ٸ�\�!ݕ������&'1�U�5RU��gMX���9s��"� g^�"��˻�Y�fW�tt4H3<5D�^�ט�����A��cZ�;V�7�ۑd9֚��SF��s����+��j*�F�+�%�nM�*���"�)�4[�����~�b�jW�O~ϷoCib�Gl��e�fr}n�Lks[�T]z�&zu�3��ɃI���*�
W{E9A>\��鷦j2��'�ƍ�K��P�I4�C	���o�����uA����Ba.�S���t�F>��]�6����z�W4�b�U���f�D"�f�"'����@>L�D��$�ڕ�M#�h.��{�*���c��q��Ty�o��D��u t,N��}�����]y7�d�ə��
Y����Ԇ�f:���&����(��o�z�6�fu�����n�� ٘��m�=.���d�i]f�cs)�<��婾�a���LB Ge�j�yw�,����+g���������'y�}uoWn�@9��	�٧����}��7-v��Ԋ7q�Rh�&����[��d�DbXcB\�EH$X�h�D��P�ƲN���ss��+bD��u�-b5eO#�̪�F�G�q���h���(L�5��(aE�YM��Ե=S]5UWQ&�3o���ua7�y�,��Le���]�u�}����Gz*�`��%#���a$���ʬ�:mH^뵏qL���Hr]/C�[�V�=;�K�WRN�v���1���P^��i��!Ck/(NՉ��4�r^7f{V�qk�y�sr;4�{�W����ŏ�c��V<�s��$8���̩��5�
�i��F�p&�O]����W��=E��׌qG���'�3��׏��逌Ƨl>��]W@�P"�f2y�P��Ȥ|��0TЮ!�(.`���w}*�(�8W�����q,Æ�^ә�7�������ީW�U'�e=��ߔam�W\�\���(CHSs7h�W8�8����DnWt.��;=Kmz�E(9�s��Mny�与^��b��Ǽ�_F�1�Lu��S�9[��Rn6���d��ņu��d3�
�.���R;<�tfX�:=���ηr4���l�%���
�H�p��n����u�����u���X�rm��8�������vv�Vϧ�]�>/1���jlaR�":��xI����l�t��ɍ����z��h�Zp!������y	Վ���y���u(���pW�]5���Ŵ ��:������cRd��u;ݔ�d��O�qI�J��s��]��8��#_J��^��2��j�c�)�״�e��zǼ73T+z��f�Yq��v��Z��IP�*
)��uB�[0&�i�HH%
��Sn-@~F.��hvF��8;T�>�:2�!ރ07��0�����<w�M�|,��_���$�x�;2�jHB�3a�o�c��i���R�x���`ѪT"��.f��R�5�4S�W���x@H�aBje�fhZS����@�\�D���]��1�E�$r���i�8�T���fCy3j=��"i�ո��>J A4���u�1�Ά��ɶ[s+�=�Â���@���cb�[-���7n�s�͛}�x�^�AL�t|�@��Ꚁ��u/=�(|mxھF��t�:��<�T,��i��ڂCp��"����]<�'��tf+9-�P�r���e|c��E��!��ł��U#����v��c�Y,Z�`Q��NS�z�t��ߦ��m~��"۷�ַ°_2���zÝg��1��e��&5j�t:�B_Y�B�'��?�Us70	E�&{k��P�j�bA���GU�wi��Ey���kAv��uoy� �����6fɖĉ���$��PP��C�N*o�4}�ì�t��m�܉yL����j�~g�# �Z_��,*
��Qa�ӹ�b��Rc��x��ea�.Ol��A5&����6��k	�YǇغx��I��l�EX�@���fgW�`��v�&D�soE���:����ee4�7�QTۜ��Z(�{G��ugr�\����{����;�g>bs��h�-"r�N�׽����.������.U	^�S�B/�n)�-Z�ِ�da�˖h<h*�p���~Λ�$N��a#���p �� �fT��o&&��ʳ=��.�;\��`1�y�뜹�Wd.0�����7x�x����.�=O'j���ҳ��!H�n-��]�ȡx��O0x�_��#�12�u7vV��OyR�H�m�Ξ�G[K;(^-�\��52.H���ݷm.�.�]X�ۏ��W3J@�����n��cZ��勬���Ivg�a��d���Gw]���9NJc"A�"���P��p�j����v�Y+,cO�5���5�#��w)n�%�m����W�AGY���¹�;]T��#pB=ѧ�����9��m�A��%�p�������ׂ�#m\*��Vn�u�
�El3��P��	�� ���l�� ���kGv�u=����4���'�8���f{#�C-���V�н X��'dS���&���Y%9G�Jck���Flh+���Ͽ=���F��nV��ǯ�)�Kє�f���_���]I0	o�����a8c�i�I�d�}�{�����Àᵣw�Q��*qS&L{9�NLʘ}��������U�M@�n�N����oi�֦$˸\I��Njmt�2�zv�	�l��I�;.�����y�Aq�j��t�c��M�C�"g�{3���^F�b䏴�s�E�K����RL2�C,@l���b0÷8D��ٽJ��i�	�W<X��z�K��W$
eg)� �u�h����]�|�u�2���� <�|��/��%K�뚗�W˺�	����w&�8�j����5�b	��4\V��Q���
;%\�}��B�Y��Q%�VU�E�������p˜�scyۃdD�`7!wv��,��GK��;}�8�{$�)~�$���n+�S�{�[cFT��Ĩ�fM���"�g�\;o4Ӈ����瞊�BNc3�[<n��&��0�I�\$��uYu+`�=U��+������PX�Z��XT�ZDi���0��Q�꫽;�;L����%�=Ac	d6�l���bY�r�{��n�FGLdRU��q��$�1O���խ�n���b������̖[���������䜝C�"GDDn��J"�I6��*87/�5Jj�*9m6�;F����"zh��҈ȧ~y7�hp�o1�90�˹���%���S��i�����!��Q�A�$����Y++�}am�xs��o&v)�<��8�[��^��V!*;8��Q���ȵ��ˣRߚ*����:�Y�
.L�b�ѽa�=Rغ�j�M�5�TA�{�{�W��{�(�Tz��[�_B:d5�ru`ʼC-�
����~�{*ᒛ��94���4�H��-u����e�<�o$�ֹ�̫5|�E��(
w�[��>�cQ�w++e��<�H��neևd�cnEm�_�ܒ��Yd�;�z����˰�.� *@��Y���Ȅn��K�p-��zM�<8|k`�!�Hq�k���qq=�zd9���v��l��r�GuX�'n��UJ�a7>۶��%m���Z�s��j7V�F��4v�拃g7b0!�d�=lQ,V4oZ�.�4&�
i�Ȯ%�[f�)�AYC-�cs�Aٹs�l MǎΙt͸�y�۲�̱y�x��k:9�#��]��z�!�9۞Ղ���w7dʇ9u��M��M����hڨ���J�4��(Q��|�wdS|������t;m��Q7\#��'j3���ds{8�'ePLxI@$�oЖrc�,,��w�����K���[H_y?h�ڀ�=d�K���c#�#53�m�ǡ+��P=U�b�ev���0$�D3���Zm�b��Q�!�i����e�c�O�e.�P�����'�(��M2��+��p��.�]��(��!y����j
MY��f�w�߯�L���Ї�S^�g@��Z�,��+�6�=�z@vx����M`��uG�̹Q��@�6�W[�K3L��s��H<�)JY���6cr�ҷz�O
BHo��Urv��m�-x�XA�o��Jѯ���)��hh2���[�ݩ�JF�)��=5϶@�tq�n���|�m��蛁&r;���Zs��c����9��QMx�	,K˚�tv#�����ܦ�����U�bU�[�[EGS(@mB���ū��T��	��[��_�'����:0�5��ز+qS�S4�w��3t��#*����ie��n�Դv��1�/_a\�H�3���r�)Zo�d���ŜN��4��'���b~RJ#a�{����֎��%)�Y�r�J����4���/���v�o廾�m��J�w��r�*�f��u��1�ȱ��sfe.Dڸ�GX{��6-�}5�o�p�UXԒ�be��f������C:].����4��SkУz�],6�Y�\�l�ۛa��v蛇p�o�n��ٮ�d˩UFb=�K��B,��p�)5�%k;�9(c��o3���Cv��9��]*n:u��j:�˓:��K�+����v�Jb�E�t��� ]h\q�Ibm�$n��;9f�)Ɨu�;4U]f���B8*ʤHGe2L6��A0u�Wb��%��Ջ/w.D��U�?+@Б65�̧�t�TM-��2�cC��H�F=��CQ�M���6AP���U�'$��HE�0֯ܖ1ٳ�e��ɽ������
��[�"�Ξ���j��c�mÆ8m&͈��͙a�*�7v���0 +��E�����H�7�\+,f�1.b`�z��[]Rn�$��;:���;\�s�ۮ�������Ķ�p��U8�]۫�����s�t��յ6�z$�G��ۺj*q\�\��E�xp�\E^3��R����OEv�.�w:�V:闕��N]k4Po�30��q��뮝���(ۏ�D�&eA�Tɯ���b_�w|�j����l�OJږЊH�ّ%J�5�x�^RB㌗2 8���[��޾�u2[+�3��Ck��w"y�KEPP�r�ͥ[��ml��j��L	�V�zF��Q�����R������<�G�u�g�������UG�V�6N�ꡉ!���+.��}�,���ӛ�m�ת���[Jp�ʆ,�E����@��s���Sm)Kǳ��cN�B�R��
�F���{ʆ�f�D�q����Sv�I���ӻ]Sj�j�E�����e����?��[�%�Pe+}�w�FF�^@EG�oi�)f�d4v���T��Vݦ��;q�ݓ&S-ާ����dI�|���-�V�͢��va���-,�DH־�)��k^Y݅m���N�8�����2�⬉�\kIeou﴾�i��k)��Ig]i��Y/v�O��-H���D�"�Y�u�9�AΚ6��f��\,�<��W"�6ͼ�":i�����N��tv.V��H�0v�hQ�U��i�^ŵ�߂�C%�+��yZ:���Sݻǥ��].|z=�G+�-(��.��	��P��w�0P�v�.��C�b���~����C,�F==TbH�U,֨�ǋ�m����[c'���t��2|2���	��U�v����} ��X4�����(B�&�H����Xs6�k���ޚ�b�k��~���s���ȥҮױV�I������.@�dM��`�A�Ү�3��Jr7ز��{י׸rb'�(u�ɛ5�2(p]�X����_i�6���
�$UH
'm!A�$X�	��hX,�z�\Bf[kb0Xk���p����q��v��'[7"$%+�t����ٙηF�K�M��a�ݯ��3�u֙�����G�*�&=��m�P&�GTu�����?w�xx��e��|kg�����P�����)�ܒ��C�޺
��oe2�.i>��&�ĵ����{�
<Z-Ca��@'f��c�ݵ$FBe
� �^��:Ȋ�ײg��%ʀVU��U{(�Ɉ&�g���|�r.�QU�q/z�B@���F5��pIZ�"�4w�p7���Rc��""hB��ý���]]	����[@�È"�xa����n��hJ�U�o#i2���F�i�a��Xz�";r�m�$|�Xsv������6�dۡP�;-;�n0_)�h*hy�Xx����j��S��f^\�Ɇ�fg��PD�=(H35\��Y)Y�W�3���!�Go/��,����dM}V��GX�b�"�p��j��6��8R�ZE;��eu�/���wL#���m��[�L�����l^c[C�c2��=�6˫����������8}Ň\�[66�����7Ѓ�ƈP$ʲ�D�q5�͔�7�݆:όltB(��x#u�h���E3ȝ�Xt������
�}Q�|�#�WN�\�M��>׻�`��21dBUp\��u�Q�� p�D4�L\����N��K#�&�4�LC};܎������:�X�ý/G�ˍ.�'<vT���oB<�q�f
p�co2�ܷ����z���a;���H����:SȘ}֤݄36�޴�gb�#,����w/:��oJy��v˓�5�e�B
-��jWw:f���e1�)���6�xl�9��P�!hEґ6p�˷�je���b��{r���Y��!��+�8CG�N�E4g(�%|톳�:Y�4C��ʝk���vQ��U8U��-.�3�U�mXv�{�M2|�ʇ͒ƺ�¦ck-�3.����a���dF�XFkge݂]>�p���1�v��gU����9I��k��e���]1��FiP���q����8��痴�ؾ����nQx�\e���{crԷd-��q)��-U9t !���<���=�� ��`Q^��Z�O-����u��]gmp�;������=�P��p��+y���[��X˭����	�KD�[������湚��,4�8%��"=�3>v��ݮ2F �Aa�n��
���=�W�B�H����zf�#�Z��c�w9$MT1�p�\d��)�J���]/(�NC����}Ҝ@'��CA��_t��7�O���V�G�F���r����'����_<�|({7I�{ӝ"cXp�f� ��hӍ�FP�w�6i%�Z���!�F�:���[4+[�3��V>^�j�T�ɢ�8��U�U]�;���-p�p����W3o�9F�y�* �C�;�'&�EF����.�%��:7ӝ��M�069�A�aCM���R+�4�L�gu�q|�f�0�`ۅ
{��3��O	1��H��>� �7��Y�:{X�n�h�8���ܜ��HХH���e�����<��A��u�����*��m��a���6��s�Ƅ��s��o���m��LgfX��i*Ľ&{�P#-���tK�����3Q�ƌ���H��C~оj˓��3A�١M�c­�b�	�0�ch�h�Ffn��3F��4f��N@f�����m ��np4.��#;��t1ZZ7`x�(�@
Q��iԶ�>�����n]���9�W��>Y��wb[�)0{ADq� ���8سpBZ���
[������:+#4�a�e�BJ��M�쀄m6GMV���c<��0�DJ�ִ�0�D鄶�םM͍�BP/�h�뛣�"�ʜڗ��XpYM0b4�o23��As�T���u"u@�劎H���$C����s�ެi\1S�7Z��PEJ�yMmc��G��r]E��M��AÄZjX����2����N���5��ވǴ��I�F��>���t��P�B�{��irC�oUv���JYP1�k�Z�X�
��q�0��n��c0T�M4q�T�#L���n�\������O�͑k��k7P#�)�<�n�%{t7Hy��kl�W���]�`�^�X^��'
��&��:f �-�/'
WuI2�`���ʚ(Q�B�\�t�B&t��/u��%�w��c��U���L_H5g�_���,[*^g����5D
L��k�f�u�\y51m)PǊF���Cb�C,��ά��1����۪��@ӎ)ư����I=ۧy��b^�5s����:C)�]�(�iՠ�n�[���CV�C��˺s�5�$H:FѸ
4�LC�Sd�p��+!�܍)�!-R.o����on�/sV��<|�4W���I��$h��R&��N� Ī������7�i�e��U�vMD�\&ZlQ��Ȗ�>�>��0Am���wd�b{��Z�O��.��e�����@�X�Um�en�oU�߹ٗ����
ޚ���.�g��笞n�N7������M���#�)��xk�~���9����|ާ씘S�Y�rȨT������$��ts�Ϧ��,g�W`�:�Kj㷁CP�������6F��ʩ�v��q�8St���?�k��H�"�W��}��7j�~�K�O���y-ڱ����Ϟ�g�U��K%��C��;�m�I�o]������dy�+}�:�{`n{y]�S�. ֫����c���,�q'�o�S�e�S7
Gs��3�C#6�Z'0�n��Q�U�N�3K�i�)��liy�QD��lK��T�[Ifej��&qћC1�^��[+��Վ`�k5���[˚��-`����8�w��Z��{�/3z�E������]��6�$�9�^�b��zW��Q�i2�(a���:�[ �y,-�	��s'ݸ'%���F����*�`��{i��5�V}���	tG���f��U�o^��7��P1���U�m�9%��a�^����Ev�f��O\�E��bU���nSr�L�����!�G�*.�x�����*�џb��Kb���d.�;�:��I��y���.R�L��Epl&Hp��"K���Q���w��鄫j��)BsQ����P�X���9~kt������=�NH�bգ5�&
V�0�!C%�j6�Y�R�v���[3P!@��9yֹ4+"��3�QU]�]gR�" k�f��:y��f������4<3|,�L�i�چѣ�X��U�槈C�ԗ�����odYQ���,^�Fp�T\�������y�(���Ԫ���f�5�b�yBȄ���5��;7��߲#����o+��x��x��L��e�!��������1����<��g�r=v4�t9�'?z�����(sMn�C8��xWS����v���u�b#�䕔k"fnT�+2����M
� M�MEӹ��#|����v*͖�Pvt�D�U�u@y��2�%�ֹ�����N��i�I�f	�)���Bkm!5���uc2۱;hCBdW1�zÌ;�V7mbs���M-�F,�7�bF��ƷE���]>��� X�����,c��q�	b��4��BV�Ƒ���j���K5��x�/���#4�4%���	���B��Vm�p�%�jF`�g�̆��3��7���Fmv�o=u���(0rg�j��Mb�]r��������������ڲ�H��3c6z��df�l��LU���N�0���?``�U� f� �ׇo���[/���*J�AC,��?���c�O	���K�:q�v��.��/N��Г�.��p]�N��iw��t�9�uF�>q�B�rӐ�p�&!�Z@b�+ޓ!%�W�Ä�(�5�hEك�Oc�g���h]A�q-������j1AF3�EYh�$ϘN!7SG��m�e�T8&�_��mb�\����l2DB�t\��n� �VG�uQl�8�/ɞ����7����Zd.���ߵ�'��j�������S,qL����oc�������&gyh�9�<y=��OB��&������Ҍ�8�[#�;/�{�7��[��66�m��ګ�h�+R�k�x�hʹ(��u��<1j{��6��VN��p�&�lw2D�ٷ[p*�g�".I����QϼdУ�2�b��ow���Lj�ސ�o6F��9��v��߿�����UP��~|�:�E/>$�v�BWVe�%��pvVL��F���__P�����ܵ4X�@�kP�ywF�^NW�'q��@�b/v�݄Z{� �Q��=*n��38��n��D��)��yF�f{�(.ꛇ=�,��h�����`�M�C�,���'<�"��mb�A�y�J彴�c��|P�]�C�w>���y�Gm�un�܂���S�	c�th�:��[;����}ϷǱz)&�����#��<��Ŋ�|]����w@�k)6���S���'�N�^�N6����k�FS�҆�D$�ק��b� 7j�~!���%�b���f�G����բ�����O͘KL�o��niaWn�3�{�����z���*��o�"���;ͷ6ݮ�툭��m�u�v3��$��s�gg�M��q[ͧ�[�@i��pa8P�"��˒���*{q�}�W��(�HA>�x.��Y���Jۃw���T���ࠏ�7�:��>�[��?:!�5���B}�ȳE�R�<�,�Eu����ۙ�B��U���X2��g�Y���-Q�D]��ԕU>��3HEc Aj���4�o�&��P�"!��i�&�/���Eو�p,��q����������.W��dɱ�ǫc�m=��[FQF��.��%�۴�N���Z�A14J6�ĉc2���ݡp	f�5�4fII}��\D�L�C7u���癩Jf������@�{M��a�=�o7���w0����U �څ].�u�>ȟY`�2�c�����><=�hV@|j�cb�;��͈�%[���
�	�A(���������Z���ꙷH��U��ۨ9����m�L�A����́�F���9��,�o<��l^�;�f~:y����̛|,�ׂr�*�i1�S�3�wS/Mp`Vي��˘�`Ż��L���6�p�/��̼�5W�w7{���V��r	�8���Aeٳ�0�>�s��3�MJ��m�D�p�,@fa(l"a�W2�q����tz4�x`��|'r"���<��0y6�)��W5�d�s��Xn/�8�0��*Emh�ê+=�(\�fnF!3;�[N��C����9�3�����.�	9�ua�=���6��5�LW^*��~.�j�U���ꇧ�b���텖W�&�̭��	m�b;x_yWvꬫw2�������V���o��98��Z���E+7�F���o*�䋻r˝}Yk�ΧaVP�
��e�%T*m����E�m��j�gTc��Ӣ���kXƋ���=��̩�[��Mz��{S�_
|���`�%2�m���Z�̛,�s�|��P��LU��Og�u��o&��v�4q,�qr��C	���ا{�����A(B.�e�<�Վ������Z�S@{c4t�Olf.�V�ґa�cgdQ1����I���6v�.=����TqN5�E[��]]���GG%��Zt*��h[�.U�+&\;e]p7!G6L"���	�5�Ǘ��e?.�8kؕv�6�q��s��G�ޚ��t��kHs�Y�茬�*���bp��^�@'�$ֵ��Y��'v��u����[^�؁�&	[��Gp�2�}7n�lB@L�9߲��eg|`��ͧ0_
��S�u}��2�N�����a��2�e@H%K��aF^�/k�.�+1��6	ʁ��p�����'�.x�sv^��}�Ϲ��3��X������s�<� �'	�e6ɆұY��^�7�ǌ�˦��m3w=k����&$@Z���S�d��!-/�*�")%��"ZD�Vr50
`�e��	lͼKw2uq[���}�j������N^%l�&`�˳(�ӊ}ұ��o!�0���}r���X� ��6T�R�X�H��Z��3�e�l^���V<�\�A�9�
xx��ת�fp�b��p�~͇)CY��5y�{1�\ʡ|���0�R�ìc�����K��ډܯe�H�T�3fA�ƅ�5Vy1B5��ˁ�H�������f���K1a��]�V���-����X�՜W[[ɛO�� wua��72a�pN���<��x:R-]�����#�;0�ӣ��>O,�i�÷�u�g�2*p��*eM�e�IŢ�%k���o^�
��4�����]��tn�[��Ƹ닻1؃!n��ʤ{ë*����1����2�q#�ޱDڽ�r�i�H����r��9�!��B�Z�f�a����uҬ"�cA]��Z(S0��0*#���}zo��2�#M���YB�9�F�W�\/��[�ʫ����UFE�:�$]�]�2"[�f�ը푌!����f��d���ݨ2��[6>�8c̝�(us�ٝt��ʄv���C1�9Go�� P���VXSkv���ˀc�b��v���Ws��qgfR$#ݷ �%��U@�fУ.��|��N�vpͼh\y�3F�0�*n*;�On� {cNڼu+n`�[�;.��f�g��ݧ�Wu��q�X�,�;�֬�4P]��ͨ�S��*��&^7�_J��9��7 2�o\��ٶ�GX6E)S�ި7Ww�eD1
 �,����E���фG0��K�.+��4�>�uvxܢ=Rd�������.��t�� j�\�"�PK����;����f��S��eغ�K�=q��Cԉ=s��5j2�le�t��WE���aɸ�p�ҽ��b�̺�������Q9�F��m�z�h�Z������L����1�6+yƉk.�#D5�1�l�.Kc(��.3�
�E�v��X�m��'�f�Sl�z�\�uۊ�^\n����Hq�{Ws>^�N��d9]��,��6ٞS�:��^�o/�E�/ Bk�$����W6 m\˕�K�1�#�]4��Y\��-ђ�3�����v�M�F�uy�!�bT�k2Z�e5�\d�4�,��+e�m+.WlK�t���Ўv�(��x(ٌƗXوLr�c12�11�,���F��u�r��5Ή-�J�6f5�)\��r������m���H��k�
�<��۩ø�`c�v�J��,<����x緈�:{j�1�A�7�f�w�6�Y\�G�G�/9V�-�;q��+�Dby���ۍN�rb��)ރ�#k>yk�[nR�a�\�0��vm�㵵��1��;B�Xƪ�A�ٔ����vo\��{k�cҚ����yisrNt槷�&��d���va紉��1��v6T�銢�n�T��sZ�[w\�t�W��;Ff�\����9�u�%͞��:��ԣ��@�ݫ����5�����ϥ�Ib�MXJb8,�� 3Ɏ]բ�L�v��U�+�b��8FZ����K��pѬ3ac�]���"�wup�݆�0��r��CO>��8�\]���F`�����̷Me��N%,�R���q�3P�f�L͐�ˑM���m��x� ��έ.k�V����r���o��1�y1�u�bi�ٙ��n�\F-8Q�u=e6����=l����^��-k��m��J��#us�A�)�"݈]���K��! �"�g3g7C�[4c�So%�������W��^C�nW(gf�kۭ�9���'k�����n��ɀf�6ˣEJFk�[�b����u�t��F����g�n�x�x);�C�qo]���P�R����9Py�Mf��[&��UI��Lv��X��V6˩�k�Q�$ZFv��v��%�؃������7Hs�l6�*��`��@�U��A��_ ��N�vvĬ�ЗB�9�T�-�h�f�e�lM��#�X�*t�]�n͗ee�Fm�շ���kM��-������/ǅ�e���g�^�Уҭ�2��܋_�g��v��Y8�m��Q.1B��Q��6�Cf��b
Pbz7�e�ek�����Jݬ��W���
�����B��L{8����B���e��C֌�H�lB �li��[�\�D`�ʵw�ԸdDT�k�C%����\��.�s�t�{ʰ�m,��vyM�"�&Nq�_ݮZG+Q��%zup�m0��w����k�Kq�+������2��Ko�Y�������&�}Z{�l*��n�ˆĩ���b��.`����M1]�fd�4#����L��eX�z�"c�U����|I�&�����R-�X�D�F0v��z;bc��1�jO�߱_�<:�mN�J��x�PnsDm0��K#P8�_��M,�[M4[\�]v�b����}�+��S	75���a��6�S��*>�]^��N��C�|��f�o'�T�yE���X�û+�p/(�Y7v�Cݬ �W{'�\�V��,x��+���Y�b``~=�;w�����7qc.��҈g�v����m�\��u�c�k#c.�[[�ƈ�
��Y|��dm
�7�>0���#FfZ�)r
��Y��t�=Q22�]�t2e?��~�}�ɑb�1�]�������(��O�]�`��w5�7�������D����yx�U��\�ى��zIՖ��C�I�_:��c0�PI0ث&G0��y�7��"�%�>�֖�m@�ϼ�S>��*��Z �k��'�L�pC�nr����8����S{�(_��alm֋i%zǙV�^;�˻�`$Y<���li��iy�/%��B�{��)�N�u�<��,��QXwnLvPy���l�7$������a��p܏R����� M3�.H���.�i����9}b!��w�]��bs����S���^,�j�lq��[��>���S�g
D'�O�#��Yz{!�]W����,K6�V;%��1VV���>�M��z{��ۏ݂���㧮�;ԗm�桸=/�VH��Q��_^LA� ��DD�M�2yJԫf��) c ���i���lM�U_�=�u���Oo*���ú(4�*ð�D����kQ��ᒅmc p���R;�;Y��f,���:�f�Z!T̳��#l&�l�e]���φm���*FМ<&!t+¨B��.�����$�AP ��r��vq6�ޞ��z��;
8�y1�k�_�����:q��.��"rb��m��e�	t���[CFl6�@w�'�_�����/����~}t<IH�,o�.�A��Y�e�iB��:�y���}]=��䄐g���^U��� ��P�5��g9��nێwr�n�Ųumڤ�.Ws�J��`��2�f$a��nD@�Yi�3b;yX��areN�Su6��[�8+a��~���/n��L\�=V�=����ϊ,��n���(2�ޤĊ���!P����aQ���ΐ	�.Խ{��.P��.�k����d�M:�7�۾��|-=���b���Q�7��	�;�K���h2�߽�"�=��'��?&*������f���'<ܬ~�ȼN�J������ѳ�I#}��X��V�^u%\����u��;��.�b7D7�"Յ&�]G^�o;ν���Y���s��mc�u 捦�����W)�L�+52�*F�j� ��U�W�zc_�{4 h����(9���G�d]R�I���ݾ���
P�b=��݄Y8qp3�<{�^E�ɘ-ɿx�Y��Oz%Z{T����/K£*K{�d��eF!�8F�H��s���R�� ,�y"�w�y��m�i�b�S�L�٭�\��F2ᔕm�O�oٸ�x�N��.�2#�yޭ�$R��.��.��P�N
E�\%�QĚ��z�m����������\�BX�dvU9�"a8W"d��G�y���b���<؃Y�F�$Wʮ��=�{���l��y1^e:nX�c"z�'�m�t�BO�BM���q}ʡ��$h�����wR%tGgٙJ�.�8]e7<��t�3���j�q$,=�j�!�3�%(yFG'ܛ�@��Y���/�}�R�Ǖ�n�����5D&jD�r1-�Y�E��jQ��)c��w�m���7��6�o������y����(��/&+d� z�YI!�/mdηK�x�R�'74S��B�}��������@I����E�}�z����z�ዛ3�Ay4T�Ld�ŝ�N�A�
�D�Z�G�b5dl2i����44�yfᔨVI�˻�{�V"��x��������M��\f�z�wRG������IBXת�`�]Vцeh݄6�p�<�*��ps��	��pg�ێ�^-Z�Y;m=������<<-�{M�y�7Z^�ly7r��G�ǌ���!�;O+z9v�:-��m�x���..�`�t>�m�N�9TƳ��H�$=%�����[��C6f!�!u�2�ʦI�����g9�n�ؽm�x���v]��r�q�����w&3t������bg��I��.���b�o�?@������s��7�U�<��Д��_.�*72$�R��x\���n	w��Q�T�ȍ���"�Bg͖�[֊��K��3-g]q�q.b	2c&m��}����7"jj�3%��yT�:������63��cp��0�j	�����Rr\���Vc -;*T��,�Ӟ�E��д+���s('�4�Yһ�w��Yl�%Mg��j�^$��H�Q7�*'&�E5��<5�G�ǩ=��[�N�b��5S���<�W��w�i�{ʃ��rS�����-W����X&��D�]�Msw�"ano!T-@�oe�4��$ax�y��G!:��AL���'xg�;��� ���Hu�������Di�P�AA��6�J��mHkc��O�cL���s��m0I���E�j��c�>s�&n,�5+�p�\~�['�1u����d��~= �Li��1=S��V�>��ɪm�6x;�~}��eIQ}�>�G����k_�<����3����|,�|��;�a�ڻ��׻A�<��!�J���l��e�p��u�I� �X���g.��)�N��RmX�h�B�ϖ��-��<�xgl,k��|�}E�&��M��Q�إ"�HC��|�� �7��kX�R»�c{�d���[}�oV��	��MmA�];���Zh&�k^�C�b:��!4lN�}	̓YR�6*�����^��r���=��wՈ�{��;��P��3�U��:j%��e��^ϥ �!B�g:y��Ml֯��>hu>T��X�z��P�9'�wH1p؅
��[}���DO\3�u��\J=xn��7�b�H���$�����WT�5�lƋs%�����͇h�]6�<b;�+-�������Y�-���ԧs5	���v�c,`Sa�j`q�+awr�q�wl2�2��㹛�tucwn��I�F!��&L�oO��n��k��9�ګ|��E{�{N!l'9,�贉P�]U�`����K�#U����#�p�)h�xB����{�I6-u!�3�bXΟO�3��9uGW[�d���
�k�/1ܺq�dPp���s��y��(rH�I&3v�
�n�(�7J�[f��F�q���0#1oV��ErH8kr�0$�Z�q�즛�@�5
�E�*S�ל��%�������_��w�T��m�|�p��̴�L��WR�DU�������a�m/vk&�����a�Be�7�@J���0�a8E�����h�qZ�9
-,����}�f�̫� >�Aާɢ�%���@s����w*�I*C½��zq=��(�X�J��eU���m��q^�ը�Y����
,�0Q̫Y�A�Ai&�Y�,rZ��Nr�;��;���-����M��_�Ze*U�r22�%꺴�Mè��y�_D��Y<@��B��r�ɧ�����������O\���31]C��l>��n'�Lv7F*�AĖ��s�T����:� �(�i���8�*�v��ɯYnjBe��)^��[�x�r���u�9/��Z2�����H�ٳܥ�N��ʍ�| je��4|a��Ɔ+���x�b6����-���B`��Y�n^^���o�z��z����9|��y���o������Z�Y�MoC��@ݍ[Q���J�k8���vkw���;Å��2��|���Jϴ�D�%�˳<#V�P�*b!� X0�\�;�y$����.�a-�����!rx�
�t34� �؝�v���bfa�'�8�V�F���e�
	 �]��}�a1ˢ�%�m�,��5#;���7�%�cv	r�Y~���~�{~y��.�����J�y�<�����#�x���:G*|$���kފ�-���_��&PC@�2[mʘ]�/���T9�Bu��8�f�FM�l��#��9&"�R� O`V�ҝ�On�3��TBT�ۃi�q%��	8~m����<�z���5�
㡤j�_ve����2��Z�>���݂���5H�l�ظ��/-�n-�%G [p�-��Ѹ͚��u}��TDR�9�ʚ�L�F$��B���k���p[Y�&ȦG�G��zM�u�b����=d���QA�ܨ�o�ڧ*|��d	����y&6{��x��f�u�W�os<��@�lkɕ�%�g�K�D�0(S�"vfM�
��T(���v�Vn�76�O^lޠ�;8�ާl�,ݡrb[�ڦj����*SӇ�eԻ0k{XZ�:�i�S�L�u o�v׿.˫�[���%�T��
7!�6^�;��c^��y{��\�!���n�$¥ǅ7��<2[5�L�ٺj�2#�(Ԏ�m���rou��\vC��@n�	�tMێÝ^D���O+���w&��QÄ��;Us���e2��q��OB�̝v�׆�6�=<��H��0n�SA�X�D�98�7=3�w:vܛ��Ӳ���ܤq���oI��	�v�G0�8��U���NSPΊ@�[��ڼ��:큻Ƴ�z��0�TǙ)�㳢����)�5�����d9F�5� ����H�j.�ת��y��5�,�s}�vS���N8ǉh������߉j.Л�{}��}�+5�𽏫�_G^�X����J�0R��u.�s��4�}r`�\i�ԷQ�Co'�26"��l����Q7`���It&�c�lUv]du�=q�}���<����\g��� �
�p95F1����J��HE�:x��m�i���lU2�y��&�i��K���#�ۈe� ����ԭ*̲}������F��2���ڑ]�Ub��P�0��<��i��	��4�V��ʣS�����Բd��
þ�PăyM-�3X&{�f�L��x�*�ɹntd�q���L,��L㲹"J�$���W\4�����T�%�r���v밽�:Cr��Ԋ�0\W2�ّy�7eΫ�]��G[�y:n�;���-C�D����}�[F�:�/n��������F]e+R:��ggk�Qz"XI�P�hN�ɀ�$��\
�e^�Q	h�V���
v�^^���}�V\���BQ��c�6����W.�P�T�q�U8�N�Q�����	��;�ڻW�<�}h�F��m'���ǽ��R�\�3ӝ����:��5����#B(8!�JNN34�4�ꜛ��Բ���y���W��e�׎��z��<�w�B��Qטyt�ˋY����g��<�in.��z����ű�ޚ�c�JZ���>��r�����5�#�=��|��N��K��5��S��z��)h��9-�^�la�{;�AZ/lr(���~=�QWd�c8��g>��w9��>�}V�S;�%��_�w�d���l�6�(���]?�.�������W���[��m�.��#��1Q*m����dM��k�V&��L]`ȩ�<��ԡ�,e fk����g��o2�=����+���u,�X��v,����HLI..
~A��"m��t������uq���j=�(��d𹞁�"�,�}���,���F��5�a��'�b7m+<3)����0҂POŤ�ʪ�<���{=��yb�B��K����꯼͢W*uAv��5Caܬ;$�y��q)�2���{�"��E�f.r �z4�U5�b�k�y�3^-�b�r%�α"�#lc��,����z.4�Z��LN�}�@�۽�7Ϻ1���ՙj�Mվ����Âf�<p7Z/�
���n|0<����9�﬩Euhǝ���^�-z��9u��u^XZ�ۮ�t����Ӯ�;7$����C&}��_ni2�y�)󛳉�8�݂mud��9����s�:'ѕx�4k��:���~��xU�F��ܻ�m��7q�x��ct7�Y�Q�v�O+(t�{��b�bn&"`ٜSē6pAn��ը�F��Fm2oU�XwH�(�"xx�X1^bݖ���V�̣�V]���}z�v�meM�R���%�3osT�yN����g�mJ{�V�,���`�]N�`ѻsp�Rӵ�ݱy�u}7k��@�V5��������C�w(�m���р�v��Y�jv�p�,��6fDƓj<�i7��N#���x��)�s^���J�Ό��[d��ɀҹ�NbFƟ�`���%)�F(��i7訔�Ұy*#:��f���3`��b����'8�l���<lމ���Q@e��\�x���l-��+��b�6'�6�"&��56=��-e4V.#m���̄�Y���к�9�U:-�Wk��B�����^�2P|.������o)EYVtG[�^��%�^MkA��1g�j��y�k*���u��t]�����[�g.�M����7��`���'�F.�7PXF;�bF��ܘ&�5o�u�;#6��=-
���ef��N�!ʙ�0@&��������K���j��~�چ�M6�&f�B.�w=�6���Ƕ&�ğV�o�����7�ܛ�.�#׸��b�$��*�����F�,�긴��l�
�''�j�h�[�&��D�I�l}�á^a��df��5���S�4VK>�QIY�3{�:�흦�_x�>�}ڵ��ji3������*9Krgri��|ny糣G���0�#����Y�e6x�f�_l��3n�F�|)b�6��׬Qč��U�"	dbT��s���F���MA�w�nuXu�u��~L}mX�2�-{����+�4�wn�o�v��x�Q�^9�i�����Du9�`���KEcǰ��V�aƗ����O�/M�|بF�6�@A2}	�����s��u�쪡��ޤ&bd��UDB��B<IY�m�534�v���w'�X��0�
W�6�v�ֲ�x�ڏ�)SʌQMx�}��o��͞�㴭��2RC<��,�P2�Īv6��� �Z�����H�X�a�W&]�� ��xg:��f��_^��F�i�Z��\Tg}RC��ӗ���ct�4�f�E�a�Q�8e�	��d��6�b?dg)jq��"��6���K�Ƴ�b�=���b]*�"v��Z>~�83n�뷢ߋ�Q��u�������:;	�dY��Y�ЭsV�u1١s���eD&��~D�k�T=�*�e`aԀ=��@�*!#k<G��8Ϗwl~n�?j�'މ���)�7b8��$�B��ol	Uvu��*�rM�a�7���`�X�±��#�<r͕�J�SS�S��� �wЧ":w����ղ��iw�=&�^�������K؝�/H_Jba��b��y��3�M�%x�E�e����x �M�N��i�r���=Ό�3��vgWs� ��uc/o�ӛ��|O#;jKZz�rS��P��s���	J�� Ci�ɠ)ܾA��M�upi"�ӔIͦ�>��%�;��v��(�qb���]]������EgG9����5
��D"3��������"^e����Fi�����͞�s^ʎ5/�I�w8�xoo��Tӭ>N�[��$�a�P��^<v8r�ȟ^�Q�1�K&���!c�����<.ێ�8T�I� .v��m�/t�[�� m������n���	��ck/e�/[e����i@�P!	��`��%����@`q�;B��5�`���gţX��ƍ1K4qq��鬪��z�78k���p��ѬC��{[�͌��jC,�6�]1�N6�A�g:�89-p�ҫ�N7�/=���p����y��WZd6c]`�8#�4�].����l8H#Y�D4�,���%'����?������DR��K8��S���*՘�{p�Nt=Z,����a{rf�LNlC���{��G��V��8q�����~8�X9ʂ���c�R�d���E;&*{}M
�sX�3�V
���._CF2����&��n!�5�@6��}0r�3���zM�Q�cW�VϏ�Rm��}{x3�׶UX���,��|x���>���i[m����a�m��v�}������'Wq�eEʼ���{kӌ�.����#�ҋ�3��4h�ؑYD�Vz��O~�J؊߀x�=�)�}QZ(�qZM�L(��72;��
�Ad�{n7�j��w�ht�}�KV8����}	w��c��:���B�vޠsZ�y��§�Pl�6�XM4k[r�tk`�W+��`ݬ�qL��6��Q��bd���&uH��:7����V��r�;v�JH�Y)W>gt���;�N�P���]m���׶��)�(�%�v���n��y�=|�C�θ%�3��٫�j1ݒ���B
�u�.�
BD�\��Nd'p	#HCh&bDDo,fZc���8�YN=U�m�Mz���5�f��k�ν�����O�yf��c�!�.��f>�V͟^ܺ�1ȸ��M��@���6��U]N�i�Oa��@�{9���sP��rY믍=�����ﱹ\��[IFk��eJ,�0��8����gb�oN�ˊ�(���2����E��w�}2���t�r��#�9�s۾Ƒ���	f�W)�L)� &"�Lcm���9+<��3wnQ{Q���u�����W��w�'/Z����V�X��Z���n7�LuFE��q�nl[��+{�:o��h��5IH@��ڹ����͍v�EB�K���ü��n����m1�n\$����˸���١B���{U�ręr��s
3�t.��'�e�F]��*�у=g3����II� �n�W���]��2��5��������x�Se/5-傰��V��|�%&|r��^��K��*Oz�������h��H�0ᶳI#����J�ˈ�|�d�::�Ñ]���Z�c����b��:j<,�:�;�O�[H���إ�k���|�U�ɺ]�5���Q��#Ҭ�Iq�4�Ťs�*92�H�3WoA��ܰ�C6��%�Y5=0�Y���"؈3�w����0�a `6�cPz�6����s �ק�2�f��mp�c�*�s,��NY�
u�O����w�VLy.{��on�$�Ch�р�44�bAc%��c�H��妍�BVpۡN&���r�j]�-�.�S����\���*�u��\E��7�
&#����CڊI��FLqF@4�&��qֺ; I3�k��NKg�bD�F��\b�r�������V���T���Q�9Op�j�����|�#��hM�t�;��s7u�b�1�z�w�H����v�+��ܮ{��p�j���sxi���u�
�JM
	A��0���S�s"D�&��TeeR��!ƭ�Ĥ5��u�[�"d\��zy�.�n'�:֚�x��)�K[l�Y��s�$n���÷f��5�7p̍�U��Ϯ�^Vwp�!a`���-�a6��p�lȦ,�\�̦b�nIU[\�2��E��m���h`V�z웆��꯬��hgjGX��7�eE�乊+��.���9[kO=��[��]�c�H~���QT�s4j�q�S��l-��ѻ��£�O �^K��-j�Ÿ&(=d�2�e�~ ��]�M�Co*��o=: �TEE�r�"��j���P�"9w:���@cJ&��渴H�Z=�l"���Գ&�+��"�X�m2����l��:#)l	c����	���$�n;S�"��q�+�uK��j�a��50A:��y���.��e$��i���^}A��^8���m��M1y��5 �="����b�$�Ľ�tOc�<5{�zQ+�o�>
�̬C]s<��Qr{5��f�*���f�Q7�!̯��;>�-x�ݼ�T�D��ֵ`�M�zK�^W��&_��6Xè�P���b,m"VꊛD#�m:��Ht35����I�h�u�?-�]!��x��<T���(YKƲ��7p������c�f���<��K�2�#͋��b�U��A�6�?n�S����/����Y;o��{�+-ep��2(s����t��⺴��w���ov�?������s��;���B�\���)H��ٚ��fpL J���گ7H,hYp!�kb73/`�"�1g&�`�Z,����7��������&A�s�q oҸcv�2�n���J���\x��ê�vF��w^ێǆ�G���h�<�I$�r�]��h�i�ʺ�d��&n�bڝ.����j��9��:��\Y��`�i- iu�5j'$��+�<�j��]eÆ�@A�e��@y.����l�'�om�V���:��e��i;r]��P����8}��9{	��׳kj6;h@9��	n�۶�.d�O95�A��z74��k=Z2Al� 0Xa��N'��2��\���^x��o��պа��pS���VQ�{�q��0%�4d��D���!����>��'4�ه	����H���?�F�n��N����Xw��N����7���N���.�%�{�[Y������.gx�eBi����[k"���l!�imbN ��i��݋k.�!:/!:휂�`�ۛ&�r��n�A]��(9�����M�$"�/����趸4yݫ�|s;s��f�:��<n�eq�U�!Ey���#�1@��oAn	T�4�J�4c����kH�R(0\AI�E������Ò(��r?7Wz�k�I���tR�\u�����Cl��Z��T�>W]�c{�ݒ��S��2���n�.�2`���R�XEm4�[�r��<C���I��Ve%���|���8k��T*�1Y������f��wv�z+�q��=x��Y�_�RO"nW
"}��$��n!6풹_���;����e�d[���ʐ`���͛-�7�`fi��6s5ջ^q�"�%Bt�NG7�P���~�^�4����ն]`��7Zf��?�J��Yq9E�^��XJE��]��Ⱦ��c�pW=J0�ͽ&*�o���ʈ��A&�H��Ť��;��2����r�DvX�Nb'u�e{��a�&zT���i���et)"�5�M�|pA8����3`�ws*X]�w<�(�&[N���TbW
���N�	݌��"��L����+��NT�;W��PFzV�����ᶼN�q����قC���I������rk؄n[>K�冭H{�ӯY��0�o�t0j�&n�Durӆb�4g����j��y�w�ָ�[�"#�n�b�M����Y|��&��ڂB+��1���Pr�,�%�&�8pS�Jm}����3%���v��T���8@�H�I�����⳶z�������75	�X��˒�D���Ģ�1�06�[pGԸ�
'�GN��d��"mGk�dE�lEu�ch��;�q��-�^�ŷr�+A�u*���]3gA� � �S��l�p�:�gz���	��D
�W�puo�xi�J��o��a��j ��	t�˦�g7�}�n�^��~���n�[��u�VK��(����DA�è���*1�T�\�z[A^{��KF+��3}�� l���fn�k�~�6hfh��OSُ��{?�>
h������j����2��⴫'K�=t�mw}���c��sP��/$UC��D&���DA]"؂	�'�:{��n$��(G�#:`�"㖥X��7	�,抎�G��T�r��:�NK}}�tc�Ku���M�\�������6��.y�6�:c;�i{m��$#zc-���tWo#��I�IVө�5��/b�Q�b/:�����W�*K���b�3�W6��J�u;������{h
T����Y��� �8l�5�4Z��{+�9tU�w[��^c�x=�
�ٶZP�`�{Ǯ�Q�C���Ю���F��B�"���j=٣")�	���r)����]<謜{�ܘbH� �D�34��,��ʶ�g����ƀ6���f�*L����BX�E2���A4�FSd4��21mu�3����`��J�fFo����Fߌ^�<�7���mM��}��J���F0_�/��(YF�8�l�}�7m�W,�їƖ�p��Ի7��m��]ڥ̽�}ǚ�ޚKu��|�A�$�q	�EdSJ��4��K��n]W�"�tm��ӇE���z�pNe0���B;<V)UDH���ip�L5�MsbM��fV�[��#�E\.v�-�HeD��Ie���v6mdc���~���9fˮJ�I���3z`9���\���A�qb�3/n����3]WN[h��߃쮤�6�*�S~�Q�O_�Y��}<��4�o��*6�I/r$P�g�Y�\��TȨ�ol�'[�����"6�	���BT6S�!�j�I�V��A*�s��U�3(K/l�n
�Hᔃ�31H,��垽�w��gײWMk�5�Ε�ђP�\Q�dm�Em��ж���=��U�R�7{�7�za2PkjX��']���r�.�s�g��^����A2�X�o&�Gq&#�� ݵ7S������>�ml�����N�=~�U��1�Ӵ�+��:�蘇5-KwX#{��u�>L��(��ߥ�� ���4�\�E+|��/n�ǂ/-fڲt�M�"LN�pd���yux����9<��h�x,hZ�b2�DlΫ�a��J�J�+����5��+�-��̸;����f�a�t�^V;�kW�)5�%�5X�j�U�w*{�����/4<X�
�d�]>�qY{3��a��S[��*�3�U�A�~��J�mRSrN���,�A@�)��{P�Wi�2��oJ����X�H���ht�xe����v�N�B����9�)��2[Ј����e�؝^�ceѣ����1���yZ����H����D�}vg;�G+WS��P�p_`;��"�9����N:=X�么�읠Wnv-�|�M��WV�U�1f��P_05��|ph�Nʻ7�!k6h�C������ؖ�޿���*p�p�$T��mf*P)b0(�^����lS;ث���=�N�1��5+����N_n<yr�-4�,x]��V'=k)u+��(<Ǻ{;TI*t� �����Ly���h%v[��.[5ҢI��H�7V����2��Yv�&�ol��1�5�$o{!U�t�\i��n�v�ކ��W8Lu���O����}Qf�Vop+dS����K�:_n�+���v�}6`�d'�2�̠r3b3n�U�K 7�8�	.��-]]�i�g,��ib�	�iYBS6o|�Y���9Q�6���q����X��Ņ�ܭ7f�*}6�[���3e�c��B��@�b0�7u?k�rʴ�v��n[-`�:�v�V�\Љ�0e�
��S{����s/ńn��-	K�����	m�.ᣗ���ˢ)����M+�:�:`���2���kd��$6����h������r��s���;U�qh�L���ծ�d�K�����D��=���4�<V�ݟ��b������7iZKY��/Fg��uvl,Ɋ�n+ۺl!Ӌ�����N�¶�*�O;�8j�n6E���3���uP^:���ܫ�\gq�M�Lj�PL����]1��[8�w�=s����WG[r��6�kL؞�NM\WK#�75�[�ږŗV,M���	�g��A���ۇ3����t�y��v�ݺT��<w �\�Ҝ	�:�V��[���D��&&�JR�z�5���.T=��ɐ|�v�����v"6f3Eruon�۟���g1�!���9�`м���.����3�;��ǀ�U�=k�!@�z	��z��s�¯3s��I�܋�����Δ����^^#8�ru����N�����s��vܮ��-v�wl\=�|O^z�g�j&��f�pII*��;V\��6ǩX�R�rf+3� ���K�v��d�e@����]�hl41ƛ���+e�j�����x�]�9z��e�pץ�AU�&v��k�fa��\�lvc���YL��w#�t�g���\���v��Շ8�z�l[�}=���0OGvn�p�[��������fqFh��Ɩ0	F�F:Rl�$Ьڻ9ܻ��^	]��1�ƽ�vd̛^yG�[�@W�\jө)��Be��X61Þ%���0R�p�#2u��3��n����lL��C���lB��=�)�n��DsΘ�m�פm�_X�.̄H6l�#���e-�멛^���r�@�tZ�.9�������nrlvn��,���3^n��Z�XAL��b��g.���r8�Ъ��n�i;��y�5�X��>r���v����@�[��csX�F�c[��9��[�N�I���.�=�饮��P���SJ� MD�ͳˡ�m]��e[Oʗ��e4�ivb�v��'X�����g`-g,u"��:�F�V!Q����+0�8F��1����"L�L�J7^"�j��[[�9C��9㍌��⽀�8�F�j;F��\�]�m��nY�oc��`�l0ڻ��&�pe���qf�Ь� j=Is�0�SM�v�2��ҝ����3��7;�y�n9v��G�3�}��v˴t%"7+�v��4�)�kk����Oc;7b.l�9r�0K��r�l�WV�?Y�Tޱ�W$D��o%ɖ6k�6�L�`2a�{:�dv��}F�rNYx:�M��`�.����t����I�B������H����N���[$D7�	�^�i�4l�����:���6���&Z���/���ej��4�4�o��j-���{�<�����>�!/vz���ͶC�I��{^f���+�de:�N�831 ��	ܽc:��ܱ��]�:Ӝ�3�}W��o�к���}ґ���^=�G��{Χ��S}�#�F^��ۃ*=4�?F��4��;�Gp�|�Q�^���J�����!ZO$8C]��^5��!=w�Y<�y��53S�>^M�]�}ba���Y+8_��b�50}�1�޵���������5�Ya�b�����Gm%�j�v�mj+��hJf�W\Ms�Ղ��F�a����k+�b"O�^+�7�ů�YٕYXuȫ�w^�l��Å��P�D/(m�S,�lnю�{:�*�d�
�3���7����Ճ [>뱽rk�t�^���M���;�+0�q*�EEb��ٯ�ި��۔-�����Z��;Ib�i�r��mC���Rl!=����(��N�ԑW[4R�|���l�ec�w&G,��l��M��}���|��P�م��[=�Gk3�ߨ�8��m���ɬ�t!@���]fC�6R���"i0�I��h���5$[{խ���o����y��v^�N�C��&A�Q+��v�(��G�4_Mӎ{�M ��<�}nx�?0��n�,Jl$4�a'�Ev�f��y�ݍ��%�6:I�FpM�u˸�]�ݘ��|��˜�R�
*�Z��`��CK)0ӊ�56��&�tm6�Kr��[�;QX��E*@0���t���\�V�)��?y����:�>諠��)�7���n��Ͻ�����c�ݳ	�*Jv$p0LE��D���\G+nG�E��|����3����N> ��2aT��ν��m����V��.|R�N��^��[���rrQ�]t�U�/2�pReMc�����ٽ���������1�^E(��ᤛ�w���.��۩���2en��X��ow8�����a������C��cx�}{c2� ��-�F�k4$�U�[�O��X��y�]\+s��C�D�[]�H�M����Y
+���k�*wۺ�36,`�	iIÍ\j����#N`q��H�CV��z�ݣ�a��:�nQ��W�o4�$�I0�7��T�8S�J��V����0�|��.W�F���*M�"(�<�[!�絢�
0㳧�}�zy=Oo��c�a	��KQ��a	
ң�ݵm�.2$�cV\T�
l���*G���m��4��B	�9�/��D�8�s}ʩ��^��|&zA��ED#vbbI�ܑ��p�8B�G�oŲ�m��I4E8�����Ln#f�0��0��2�'Α�F�6:dFftL0��=%G���v�0��k���Ĥ�dɶ� �&��xH�����Ų�S�#yY&ͬ}F��Fʸ�7RV�ΘUy�^�S���-P��[EJf�h��aE6�0�	��L��ܙ�9~�K���7�y,C�qf�sT[��Y��ؕ��.�6޸��\oo���V�sh����4aj�A���ᷨ"�pt"�7�͕�m�9c�ec\w�
��,�Y������(`��5�N�ɞ��~�(#�&dL���M�%���I1tW*���#p��9x-+YN�=*�BG���K(
��Rߜ7x�Pd���czz��~ح3޲kNS���smD#�"��J�(!��2�W��g\��v�1�����h�4CF%Zl��+BI���n�@�p����]7���5�;Ҽ���e/M����~��^}y�5�2}z'��G
�
'et2c���W�C)�\�.}<��*.`�|��Cp]Wu�F$6a��-9�/	�w��dܓ�������GR�}b7�yU5"�t�P�������FȖ�R{��+i�β��Z��۴5���[��f�9�[�,:i'��b���p��VpA��C��h��ʻxB��t�TPy6a΄�hV@��ܵQ�Thd �=}\��;V�-%*�]���Z�ٺf��}�t6Eü�B��"�4!�P�D%13A'���F����{�
��4ju��f-��'		�F*;��SC"`�ue_b$�ݷ�{dy=|W+���^�����\�(W��t���Ϟ��Nkf���&5Զ��Z?®��L,��2��c5:��%<[�n�Y��t���<�����CYg��
���'C�-�K7m�c������{��]t�7;�;t���5�ă�������v,�Y�hK`͸���vԱ��M&,\�v+Y����%�[c�y��d���v��;FM�tn�3�b��W=z�E�nv��o�돝O�e2)�����34ҋ���4��,�C��Kh�����z뜣s�Wn�t�v �ƞ��v��JQ�ڋ����ˆW���7/:ܾH��XvP�t����E˺��C1ȶ�"���@�io�?�o[ZԖ;}�Z�ʈ�J����c�PP��� �����9EZ�5��)�	��;p��M�n�a��7�a�m����6Y˄9Y�T��f�2*#4�@-�@1��c��%�3�^P�'9��������e����L�9i�8s�V&kQ�s�{�{y�$���xfb�aH5>�
��F��Y*�
�E�P.:��¹�10��4l`6�S �o�`�bM����da��P���w&�"��,µW"��&����b���3"���ś��������cm�=��M�M{��Ea�Lo/\uTM�o(��=���"sٶ�7��ȁy�s��qI)�SɃe��j��K�_]5������[�`>��X���
�^��+[d�1�u��0Ԗ��\��)��teq�Q�/�x�{�xR�r)��T�(� j�y���'���gy�&]�����`i]O����E�;X�r���߼�4?���2�Q9ܵwPq�p����n/�]yXB���`�z͆b�9؎<彙Z��6��90tD}�t�k�"Y��6Rw�' ҳ�`.�غs9���[k�ٱ����s=Z<#�'�y㻰�:&^����@[�0L���`���u^�k��}6_o�*bհ�L���P�&L�U�N�)]��DA����"iÞ$nv����E���8Ws;��3b-;>��{�<�����g�|u�j��$��������祎�v��+ʵ�i���pb#t�"�$8�.]Th�[�3�Җ^�6��
��Ϭ�Y©��)����M����3��ظ/BU�-	�T-�}Z"�Mp}���v*6�:;� 6��.c�7n���������*�>� [�,3Z�Rh�@�bJ�]Λ�ӻ��.6ݛ�Օ�%�C)��Eo8�J7T�#�]�XQ�#���'�9v����'��s�9�T����H����SY݆"����0Ya��3]���l�Jrz�y_�p���U�^��Du,p�^����
��X�a�H���H΅Q��,Uy�����b �j"
�
��q��H�QώQ�F��������:7�[��B��[��v�>ӑ�;)k��g���[[okr�;2���N��6ܫ�3w��lu���osvt�ŀ�%ϛ`�|;�	ɨ�l��-e����^��9>MV�!q�m,�K�&܀'��cx�y���3w�s0����o/7ci1��*��09�޽���=��犺���?��??�͝ga���ep�7�wk�Q�|䛂X�ʞX}@漰{�Ȏ�Je���lG:%��·Wӂ����,\��6;�kn�����O�ɨ6�ѫYC4Fy��Tuϭ�������T��h>M�k�3�*͍�.e�;P����vn���w����qˇ�goOI�:���UPw��I���b3��*�C�!Z�Y{Bx� ������zi�JL�&ݨ�Q�������3�9�d�T;y����cQ�8ru��&	[��I�Ej��?^�|��j�f�B)&ʆ�L��
�3Y靸ꔾ��g�Ml����A��(}X;��
S/2�ͻw)>�[��z�xOr���o�P���
6��!�ɚ;.:zǞ�Mf�ݱ��Mΰ�����=+`���˺��y�֪r1Q뻣(b�-'{3�;�����Vq�RҾn�ͭ���p��K�cGZ�Y��]�.�l*ZHM��wG6�F�+̼f������up	���R��^$=^S"F�l��JLH�Q&��{���� ���N�����a�\��vfjج̒*�R�N�*�rT*�LY��������e��K1�Q�ݕ Y/a�w&Tx����{B�ۡC�yu��F�Q.�o��4��a
���^4k1e&��s����Ol�d��Z%|;w�l��)K��Oؙ꒨l�6I�	�C�h����橱�Q\=N�s�pvz�̸w[�$Iܝ�x0<�rP���<Œj����� �oM���!w#vg6��
ʰI� ѭ�ubk8��g����e��NU@Qo�W[w�d:z�R�{>]��hn�s�v�c�pq�0Vp�X��mC�ۈL��i�ם̳f���HǸ�"�(����R����AA�F��u�4I-�KΘ1B���Zji�&�n0��a��u,L&S89��FT���3}IH���h8��Xu(�z㆏ ���C5����8.�C�y�v�ߢ��q�֭�Ĳ����˼�3Jwu�-Ȃ��w�R����N���$c������WJ��� 蛜�fT'�}x^�d�آnw^P;��R�m(��٢b��}��v[�,`N��»j�Lۚ�7U6� ��ط�O�v��9"I,�����vu6B9i��f��sn�Fx�o7��8z�c�O���Og�*[6��]�s�xS;%7j��ml�1�ۇx��V��e�r��{g]4��]��TY����t��ۮ��jz��@��қq����v%�&w�d2ɟvݡ�cdxK��d�Uκ��vLi൰�5���j��U�YnR��[��mh��Ů\��k=�rc���0w�����8��n������t�v���n���&��\4=��.?+I��w��bڹ�gϽ������;���9Mv�α�o+��
�з�yJ�H:�A#_\r���$i���Qw�P�w�3`����D��C[(p��p�M��%�D�t�v�'iOT�=\e�61$��1{/�=K�<�����T�o_w���O�z�k~O6G�b����kcK��y�qy�t�s�H�xIR�'3������)�sܓ�j%s%�zd�A�݁Q 4{-�����;��%ۿfdpa��-���J:�Mt"-s
�`�ҭ7/ �h����ypNK�b�uf�)�CT�����fT��W��d?�n�
�j{<���֌4�\�^�e��Wi���J�5�Ys��~z}>�a��gx��X�}�ڹ�Ͳ��Хh�d�3����=�������	��;��0�0�%�M����jJ�Ts�����Oh�]I�,���j���,\�4�N�۽�&��Zx��a�rWe���������Ш$ƀ��|v�c����O^ƜSD�XQ��m��z1�H���c���nF�Ȭ��݁d{s4���PV�,1w�����e��p�ݜ�C}�"��`��B��tj�&��߻��,�{7��M�7�(9��ӫ�jh�>����]R�너�	L$[f-���N�U��\y^�ª�YE\�Yb���!wdMl&"�u�?H��ݵ�yѫ��i���S�I�J��p�9��<2��t�Z�OkZ�{v����d7=/��؄V��*+�[4����*2���Z4�E��������ݒ�M3
��0���2�:���7�+s�Z��B`�@IS��3��V����"߾���||��ڙ�(�0�N1eC|���V����K�̼~���/�_�zb^h�|[6}����M~{֟��؎ڊ{���0�ƯV���{}\���{�#;x��U �A��T$��F>�X���#��f���I���$���&>I��`�P}�G
�+4���;���,��g����1�qtM
�H�8�V�ɶEn5�ϖ�n��|Q��*���v�����`�8N��7/i*���e�y(�/���-=�.��7L��(��LP�uξ�U�������zQ���9�]Ҟ1��R�\����'bn"�p$�«\!�0�����i��ZF�t7�×�
�O]���F^����!ǷN��ArV�vi ev�Q��]J���xՍW���uY-���.��.���-wT�#6�va"��Yd���z��lFoK�f{(�V�*u�N�5tf��V�f��(����W
-^��kr��>�T@��"��sz�k9�@�-�:.���(��ku6Ѵf�D�9��nw�Q��$���#N�Z�����ͷ��1i�%��B��ݮ�qp[��%��$��W;6Ch��hY�S�`��D�g������h�|�a��<���n��Op������E�!R�/N%�%�e��P2_br�����r�)Hȕ�/iK�#.���5dl��y�W2�\�fs���&(�{ˆaY�У���Ѱ;j1�*\,����ðeLh�>+d���Ho������)���{��;�H�ù�Q�]Z9�rp�o_d���hG�ܭV�9r�xݻl���钡���VnWeJ�;/�S!�W�0X��}��t�=��Ui��ڴxL����jcj��]r9�c�I,n��Js��ͻS�5c��/�#��U�S0Q�!n����౭坯)����Ġ��t�-���Lwf�I]�!֨�oWU�u��x��ئ�B�j����t�M<n�y�Ί��7*EOQ& �X&��KG����{a�����s]�e�M'&TNی�{X5�&\.�2���z�:�8�t\�о�R���?O��~L��J�'�߼�\�|�#���<��A�glo%N&�B��v�2T_o`�Sד��{<�UX��V���'��%�{�	����G�-LUȦIjN8۪������@�LR-0̃���6�gf`�*(-��	����X}�Sv����n��_p���┸��f�y���ga�B<�\}emL�OIEV	AÄ�,'	�ۖ���2�'l�c��r��s�OW~�2}�I�?r�H$;"��]lƎ���[�"A�8lJ�t��4��@P��9�&�׸� ��������~�텴v6��8���e�S�%��7���D�&|*b�w��t�����8�ڽI�M3�k�k\��\1p�?}�ų#����
�|(H��(�#~k	"M($����u����R5�q�7��wOf�@�1���٘u?}�QOA��2@���_�$<]���=%��h]4g�5�3)�G_�,H�oh�k������؛y��g--`g9+6�ێ���m�Y)c�B�ٷ�4�1 TTmh9;3F�..]��8VHUn0>\�����1Nk}�S��
~3�8gP�B��[��#�X-H�t��l����(1 Kg�k���à'��f)��u�l៌���т}F�YdP��Oɴ���M�b�F�D��Ǳ&w��~���<�J��9���o��������F�v�+�nޚƽc̀���)D��Y4v�]��4�,cR����Ť��Y�#�}Z��,�����-��t�%LQ
��
}~z�qT��I��G�d"�TY�Բ��/�~ߩ�T�f�G��DP ��9ӮI����y�Tf��UlI���B��2�aT��Y�ظ>5���h@8��>B;뺉�G�3��V�='�F�	��AL��O�0VG�>ߣ	���3鼉� �#���7� �}_l�{�iȓX����`tǄ/}�~���E���R;\���xm��h�d$i3)���~�Ϗ�?r`~6A4|
�/:����wc̊4G1fO�j&�_@#�6�i�ϯ���}�I��3�u���Mf, g�pH����/н������Z�u�en)BI*r��቟�ҥ�ޤ����}�y��u�1�|'��4�#/�^�t��Ix�$�d�r�$}�����Z��F}H!��ك��T~�:@���$�"�����χ�b5	"ȣ�����e���
��ٜ<��T �թ>��Ig�U���:z_��5���>�?,��[��8���@���@��K3�>@ҋ	"�����ϵ����\��5u1v?"G�߸��bkff�#T}�h5��#�Э�4,	+�<Ѫ�u�o��Ca�tm�+e�e�z�-m��V,��N�5�{kd3��� �NVI���%Q�n�2ۋ*L�h�.��D=����oB��Ok�:��6
�Wt"�\�#Y^Bm`DGF��XgV�̇�e�y��ظ�.�Vf5��6Ѳ(g�v��݁�n�,�6-��T�a)3��iJ�(!���36,�R�Q!�Jik��b�[�F9���fv�^�ɹ����Ѹ����/N�e8�U�%����v�M�hde�1֙c����@a�N��8���]��nq�b�a� ڡ�eʸЎ�c��}��4i�Y��H�_U���3ǂ�b�fUg�]��Z]
�5 "O� j�Ϣ���{'UK�| �Ai�|h���8��FpK���*b���W�~��PN+%�[^҇bъ� �;1��?9�*|��Lޒh�oR����=WdH_V�x��ӻ �xI����6.=j� I�D:��T��> ��۬�!�ODZ�,�>�$i���
��΁�/Z�x�n`	��������DMG�c�JDv$�O�D�e�lI$|xYB8"��xY��M�dF�OQ��@�|&n~R4�Ȣ��2�����|8g�`@��I,@ݯ	t@
�C���|��xدs�D�_'���hLG�A|go���"��ax�-W�Q�����'�D��$����ϔ�Gg̀J n:����e@'�﫜�f=��!T2�^ޚ�l?4���"�<�RIA��qRE��>�ԅ	� �?\`ϊ�y�|7`" ڏp�eFۘ�Kkj�O���_A}_?	>���~M�"ae9~�#�*�`�O���,��g]��:}���=�4>�@.<)�g��#�b�K�����̣f��#S-����-N9�f����x��Z^I�y���f�\��<�4	<}����
$�`}��S�dR�¼_���ٛ����`hJ���'�WU�"��u�=��탓u�qB=ĩ��?n���sf���4b�hT��vs��ʛ��\��k6.��m3)�*%K�߻u�-{��|`7>N��^�w6��T�c&�K*��#Tcm�,!EDd�ʺ�;6�����d���=�����D�
1V���v{�G�Ӯ��	{w�`υ#�Gǅ��ߚfĶ���i/��⥪@IE�>�O׷���Wr~+�V�=�b#�}%}n��p��[L$�$�xa �#����Qd��r����#�#�"g~���l�.��>��
5x�&�����O��:D�.)#j�T���N�t��@g�B�����73�P�ۢA�V�
����'d�ܲ2U$���Ή?=H˧�����s�8��C��2>#	!�2."H_unZ؃B��b�9�饳:/L����W|�h���#�ŧ��/�4��ç0ؑ�ȑ�DF`�&ύǲ�>sb8��l Xb0a1aa�)�rl������D��Np��J0}<)�2|ȿ���<��5��>[J@�v> 3[�O��r�F�$�� i��ľm/�t��z魞��b�Z�@g��$�(�uFq\D��X���Y�;!L�۱����nF��[n��Q�[�Y�m��.����`ȿ��8{��@	h�A.�9ɤ����0@��$0'uz;�0N>��2�ĕz]'$���� �U\2�¨���6O��|�Da��h��6ԍ�t�
o��#�Dy
�KZ�����[
�du;lڦtZ����%�6wmxTYAw�i4(:t��ϖ�O��<�����
#v<�v؟|F@���q ���@wѤ\C��S �<l�w�Z�A�ϙ�}9�Ѿ��~q�:}����)>��&���nR)
��|���e1A3+i_7o񥽴�Os6%�}��z`h�3��?M/�{�Q e�խ��?fw��J+���hަhD��S[&����U�B�LE�'FFgu�|m$օ�k�m��b��u��Q{�bH$�R8�a�}!_j�a?D3!��CZx���N-/�y�x˦�͚�������|Wl�X��=��p�gQ*��Mf���?868�#H��S����YG]�$��(��YFYï�����y�B��wo��H��6�,p'���F�,�'�{�����lL�Kυ�u������-�(V
V�S;���7��1X��vA|���/��R��Ѳ��$�1��.@�d�!	�D*bT���������>���^ǣ# ��!��l�����W�韸��^�C�>d��ϱP���1G�D{H����{�|c֨�~��ߒ l��6���(b.s[�b�wR���Yq�i�қF�1��6�bRC��,U<�[�Pؿ>6b���T���57pg®}�2��m}��K����u�G�}d2���Ř!�Ff �ا�n��Q�&_��{�Èʁ�"O���o�K��t�V�hG9-��l�w[������UJ�g3�N	1��&�t�q�i����$iqWc(c�܏��UZ߈��״���#vK}μ6�x3�B�<(�EL=�4}���G�B��3��|����c�{�q��w辯4/�_y���`�**�IY�"���Y��dѪ���xa�wqR���	��L.������4ȓ}�F���7�[�g����w��D�#�>r�'�É!�����]�b4�)b�5��q��B(Ä�I� �p0��	�]bn���6��ÈG�FW�j� YlzO�"ϱ��]�BV~��Vmx3﷐��̇P�eVD���2`]?CKL�]1'y!=�q�B�N���V�����٪�EΎ{����(wU��x�qH�t��O�1j�F�V^�,�>W<�F|��?
�q⟹1S[��s,�"�9Q�k��^AJ�ѣ[>�l|p_��Te��,�"�����,�|Ȼ���K�)�8�Z$�S� ���.�ǰѣs Dw_΀��G�;��>
��r>���3K� h���Bj<:��G�>�͟��f��0jQW&Z���f�u��$�����X{,m�N�s�=(��;�q�)t�]$��ڔ�F��~��e:p�!d�}Q>DM�� '��#�J���|E�i����ςW�@�="l�������#� �C>����>?giءt,�_u�3(�|���w����󕐣r�[)��؎����ƴ�֡������ȶ;�_?��r�e����D�&l�)t��=ɭ��k��(�xF�z���p6$8}!�����$5�g� ;?Q�����q�����	CZ����Օ��ԋ&���Dy�g�L
#���r�5�.�����_�p��f�3 υ��!Nw����k���">�5 }_�6@�&�I�$d�Q�~��uF
1ݴ��3_�b?t���Uu5iKl��^?:��1h�h�rQٵZ�����_���G�G��?CS�<���Ŭ�}j�a��Ui��E����~�K׳�1h��ض�{W�%v+�$j� Q�SZ��HÇ�FWN�8I�$�}��PG�I4���ƒ.��R�)W|�\��LP�Wt���@���:�4�|-@Y5�c�$��'���>��xa�4�}ۭ�7�]�d_}��È��i� ����Ǉ��ό��#݋ Y�FI~p�Ώu���X�_
XUn'
lA�kN���sj�t0�*X�����v,K����b���^dU`�vzŊ�\К�׾v��^��i�v�%h^a�T� �:�q�]��=f�J���c���`TT���CGh�ĥmqW\q��<u�j���#�Yb!	A����B%v�����X���ם]6f���7�������K����-\�h磲{n�.1�f�[�W���+�ۜ{8�#Q���{�{+��kh���Ӂ�q\.��q���f�\4�V]���a�W�#�;5K<���s�����v#��r��ne���.�X�
*]\!hv�b���8�YT�Z���q��A�jFV��Oؾ3M�bb�zzٿ��������>�J}$uʒ)O�܊ �H�0j%@�j	��X�0��~U.{��/ :#�$�U[��D^e����
4��቏g[b��W_$m�M�"���LCk�C�5�[𪾶�O�8D��4S+C��<ς�^�"X��h��*t���^l����_e���|ϵz��E�(����#&=�>*�gB������#�Ǿ"N)�p��kb�	���J6b�&~��_�pτO��� �c��"g(�#�W*|�ۏ< ڀ�U�M/����I�D�m}􀳫��Ǐ� I���3���J�,�g�T����x�#g��y �D��pZ�d���@9�� �|~�*E��yU"��y�2���fGٛ�|8�?} �A]�A���S��μ�#ř&cH
g�ml	S��b�$~��vi�=���C�N���o� �P
fޢb
2�����q����+�7k��2���l��E�0�}D��s�a��t�͑G±���4AV/�����xw��~R�3Ѫ ���okIi7�~C��a�\~*�A!���@`�~ ��"H��,��U����nGbLTZ)R3\����<;.�vYM"���<r���;pku�Z��*��J(��l���~U��N~{z���EH*`�E�,2C��:����H~�<`�ר1Q�"�}tyқ�2�������A*�"Ȓ�du�I�Y�c���9� �ܯ�-�Mh\ �y��U����S%�Jm�L�z"ضt����@&�+�^f��}�� }3�+�խ�e�c ��(4h���F��3��fh�f��!c`F�;P3B�ذ��ij��;PTTtu�\^�8�9�m��=�	t��$�}����Yf�	�uO�Lw���ʾ�^�w\��**�;
� ���w�f�r"��᯳��>���~��{O�O��Y���߭m�(\
իx��<�kH�m*u�щ����(f�~k����^��i�o)����x_G�0t�
{d�.vğ
9���r��z|(�B �#H�����"�F�}H3�$e@�G�*��U*��u����g����x�_�k�޷�ց*K5���N�[4b�����列��d�3F�	��0�& q���X}��{��/*�dY�>�����(��ϫ+hI�,�P���azx����I?Y�P�٬[0�LT_����ž5����]m@�
>�EM��g˃Qj3}�I�q�Eџ�T�A�φr�s\���� 
p$�F��7��#��#��A�M�2�zHG�#�W}/k~+t�0�a�ڃ�0��c�ۻ(���BT�N�cr�sn؀�Jۥen��v��u���,�[�I�D����o�e��Z�ђ�2
��c���4��k�"��Zс�$�57�)�9�����}=Eћ�|t'���4%}��5����ioo��BZ3/~���V�"*��jմ��j�E(��Z�\Z�G�}��n�������&�����9/�w�<��*cc ]'���t�y�C�����8Bz$��
�BO��>��w�=K1�x">(�i�����#k����9-���ч�S�̂+P�}���}u���(x>��DA
�O�=<��>���4Dԝ�^�G�������ǌ;�}Jj�Y���{ؕ15(�&���J�N��n�4t�֊�Ӵ	�Ĵ�!����������O��$��^�L�z���h'��m�/����s�4�3���f{N�1~��r���*��R���]�#>�G�L!����N_T�|}d����u�0)��g�Q��,�$��{���$a�������K��$�h���� =�".��Ǐ���ϱ���O��W���=��Tqg�`�"O������I%���\�kFw�ʄ�QǙ!@�#>�~aؑ��Ev:2�>�*��D�\�>�'��s�1�G��	Θ���S����R��k�6g�D�R��]O����g�WZ���ph+L�)���!z��Um�B&L�%Rݳ��]�]�6Sr��0�\�n1���j�k�Cqdf5���c.v�Ͻ>ޚ���Z�~4�~�?[3��^�f�]�T��}yw�O�X�?<#M�������3�����}��Q~r��>>ӳ����p��E�-��&�M/p���of* $A�T�qO���MB2�[vW�Z�6��"�¶ �����u���������ռC0B#�@ɚ�����s�$��~}s�T�����R}�T����G�}��TY�_N�UIF��h��*c�-.�I}��E�@ �װ8�	>#�U[��$Ν����S���`Q&����׆�EzHG
@L��b~��~��ѝ1S9Û>��S�ߑ�,��=���Y�Z��9�� &n dYu������o-� �m�>;���K=;���3*�,�Ǿ�����Q�����<E)�m��>�&����&�"0o�{����x�̆j��*���T�ؿi��ZT_*��M|zz-#��~g f>��R̡�gN��v㸮�z~;�^�+n��m�;��+i�˾@I&�P���eBڷZ唘u�~D����v7 ���-�I�v���b�"ݘ��iT��촅��%�i��T�= Bzp͇��95���1��K����4N�O7�_9I��
>@��+`���@G¾k������4���F��=8��A�!5�u-)��?��W����m�ƴ��f�ƕm֭�G�:̚3B�7���m\4K���2�ݪ���k��@���v�V��C64�/��i����W�h��y�J.�#���0�\� �$}&O�v> yg��v	 ��*!�}��߲&:,�dQ�� ��vdv�; �q����$	*�����M����>�##��p^1��Ι9�U������5g㭲��8���}s�g�D��"���0/Z�t�"N�>����"E�9�Ӧ�"�|1z�dF�����"*=�D��ܷ��~�/3x�A����� �7+�+�%�A@La5�B"��0,��TG��Ǉw�H�;�L1�|(�����=U�ߌ��E0_�<q�;zD��_p��P>*�&��}��D������B���k 3�w)�� ���å1~�??�r����p	V��|)�{kf-���^v�9֭|�6ϴ���^D�}p̿2 D��kF_�}���+���>�l]3G:DI�%�r�	�$�C6�߰ n��b�b}'I��7�ǘ����>[K�LAU1w����RUYp�2Zo9�u��;�
>| ��r�܁����K��d�i@DN��?�u碦��^�O��$��u�ؓ7��~3�~/�����/
�D���F���4h�
#�=T�$��i��M>F�<��������2Q�"Xp��Tw]���Y�Y�X].Ƕ䗘S9t����¶쪎mK6��'�F\�3V�i�[Ko4�Ρ�ܦ)��;�o�5W˟�)��Ӡ�)�]N���u]��^���dUH�e��,FE�v�]\���ށ�N�M�$�	9�U�(�`�=���󊌜lY{{���\��R���c��nqi
�;7�w0��Pb��L1d�ݣ��ݽi�謉}z�g��`ڋ�ВV��p4�+7q�[%c��l�w6�rM�)��`�Ӆ��i�[��k{�q�B�V��x��X��ݨ��/:
}���#
D�VQ�zi�Z�¦��fX��clpx� �ns��w`f�%.m�T��'�T��b���K�E�­��r�Ej8a������nN���^�W!Yǉ�!��Yt���i�&:_ݷqS�yHkx�Q�BW�㭚P̀<�����#� 
M\����͂h�+J�m$sb��_��jy�I[�zN��Ee�[	a�٘j�����u�Ո���)�l����_D_r�W�\ѻ���S&�x�^�e��EU,�Di[A��a���Fk��w,�Pg�%�̫�Y��h˘��phNw�B��u�����}���o�*ɚ�S����ԭ!-��]��NU�%�=՛��0W;�3:�����N���ׇgV�Y�n�)�8C�b�|x_��1i�!]\O��zf�Cp������Wp>��S2nR[��u�\s1�f�ĳw-<�Zm�X�]گ���u��q�m�4�cۛ7�[h��õ� s��Zz�c*A���qd^�tJ5q�p�'��[,DH1b[��6R�,H�	�0���smX*��)[d��6Eܞ�4#��[����]�룍�����G&훀�1N� u=ih֡ ŧen9n�1"&�|�x;��g�i�ҝq�޶�m���6$b�c���K������_���k�鸽��ls��]*Z��\죨�/�|�ټ�8����cf��X���t�d�l�Z��)rQ��yz'�-��:J��9�v�o6,��˛ǃ���8'Q�s��Wm��m�j�sF�Om>�8W%"K��i�i�����R��N�&��	<������ɢ�E���i�*C"��mPKl$�2a��$F�*m���f�[eX����͡���g�j*EL=Pv{����d���U���i��R�Yr�� UF]�Ќ����0O<�գ�ڂa.9���X{"��.RuO%��-��=���M���+0˩c3civ#��V�F�4P�iEh�]F��Z�[�}�@6������s<.�m�(�v���u��pb��i��t�廜"��ke3�ۈ2�-+f�cHmq4�1�� s���s���4�y�yG���lh��m7%��mh�a&(�m�"뉦l�Mglt�t�q�� �غ� ���,1�qhEe�1A�gqv���Ѻx�5!�ۮ69�v,�#C����UA����Ŭ���p[�l�:`e�3�ȮӋ��u�L����ƪ�^4�d�'k�p�{��7R\���	�,b�7M<���ʮ���l�Y��8Ƭ"�ִe���j��)��:�
XH�:}�㣂��l=�8c-����5Ջ��l�u�#�r��r�K�S���x�u䶕�쇦{\cN�qOl�8���Ůh1��V8C=�j�C��n�,zԺ�b!�"�kY�� �/gq�a횈�����fe��i�sZcw��oh%�Bm2F�K�	)��G���S��y�e���������9G�g@��i�t�}6��zW���! �n�f���b�,�TKc�YV�ݧos\���/��.�+V�GB����Yy�q5�ն�!5z����8������73v�v�m��
N	�urI��{&�����;h�G�nȘX��ϗe�"=��8��qf!J�y�:^�X���.�;�f�w���{-�þK�n�WO�!Oc��Ǉ�0Y�X���{jA;����uw��I9��W��͔��-I؉�� �݄��E.�� ���X���0��q/v�p�`xc�sdv ĕ٢u�yL�)��,����`*pѡh����4�g`C�U���־�o�{BM�1(!�P��}T���,���< �8�n��(��:d�}jsuU�^DhT{�L��Ϸ���/���$r�T�O$��74l18�WM(�����g��O~�>�F��$�A|D�3���2ּ�>�*��D�@���T��^�xQ���0'��Q�3YjApA>j�w�8�^G����@Ͼ�a�M&�ڵ��]H�i>8���G_}�#�lid���ܐ8�f�jdq�H�F�9��\P؝Ϣ7�>����;�.D�����E}�|\důTg��<�����iäI���}���Q�,VYn���O��5*�n:by������R�Ͼ�U��r������#�S�|>��Mĩ�T{܂�>���ILL�i}�����w�OZ:B#vl��2ȳ�<ء��˟�Ip��[���#��'ȍ�FF�SQG�ѻ��6mMs�/��?jf�f���N��k����5�#���}nB|!�G����ix�sO����
V��~��W�8aEYT��|��=��N_+��1s��k-���i��8]�R`��d݋�	wm���fl؄8mt�*�r��|�wC���4}lЕQ��?n�t��؃�S A�)A�o�����|��G��-R�"��\}W�ӑF�"(G}1Tp����$�f	�n�1�u9nB�+��4-�JA ���g�k���FKh���s�QxLzmF�BB���o�|0������Bb�'�\TD��劆\�W�i8t�\�mv��5&{bMVV�^�w1Z S1Xs1rA�F�u��������{�f�:���N:��"ϩ�����gU�}���5'�p5ڤ��/�P�q�!!�H�9ZT���<��~l�i�~�.��{α-�Iִ~��s]Zv��+"��+�D�R��U��Z���9ˮ�����Zۅ �6��߻'ã�~{��7̗�Bݞ���݅g��ŕ5T�������>ˏ
>N�����&��{E1?�tB�d�QYES,Q�w��]O�S6�%��=�|���Q����p�F=�I�D"/��'�j�f�.Lx[��;�Q8"נ�٘dqg����"ϑ��3�nMv��	u��Dlz���E�^}�@�`(M�l{�G\�ZIe�Il��*3G�������O=���-V�~����>Rr�}�o0φQ���3�Y)@�w|�I`"ϑ��8*<l��5�F:^��D���L�B�⨌��=�9}n���(D4�<0�{%72����5�#%����4�rՀT�r��+��EvF~����/��Oo���2�O��r�z�á��р�73��d
��u���\�`�� I�[�*\ $��@��O���t�����@Y��
7P�z�D }9��H��#����3��ؙ�ퟪ���u��&6t-rP�8%6��a�Dq�Q���(�n
���8A"ȍyk��w�M|����`�	:�x�������>�KgLa�D�d�&��b��d}%��q��L� A3S�1�`8i@���8OL2'��f�z~�n�X;�����L�=�/��4(B�|�ЗN~���mx�!]z�ً�x����������m04g?|!��؍���k�����;�ώH��.dw���U+���Fvn񇁦Ժ��{'5ŗ#4��B�����#�W���߂z Y=ت��C:x�4��τ�bc�9�kgL���y3�lT��A�J����>�W2E*%nYĸwĉ| �P(�ۗH�N�'"�����xB�]�4cf�P�����pgflT�N�饯���&���W�L"���/�ch4������x�lJ���D��#���j��@<ɂ�DL���UZ��<uţ�-��Q-�Y�*�� |ccI ��H���D!$�4�G_�3�@qހ4>�	8F(�rg<�����T逡���넭�Ow�D�#L!�Z� #��lQ��U��֋�}�������\hUG�j�/;HN �`�9^Ӥ�fnءjbk�z��V(J�j�gR��Q@4�KU��#���>t�|�vB� �������4��.��f��4m���9��A�7��/��pG����DQ���E�N|M�S�3K���P#yͥ�'���1�l��%��pR�S1� UDE�o�>�>G}�$*�cv�����������/���C�36=?۱)�����D��*$O�Q�{_~��om3�Lj��}��r������׌Qu@��C�>��A2�Yl�.�B��&eC�C!�6o����In>��E��L�m�ec����x�׊��}?g=��B�~�h����5���k�hfA&%V�?#_����o�ΐ��ţ?
hЧ�?�p��r;��V�lM_��*O��ס�8�D.7w�^�0�D?l� Q����T�$���
>�ٹ�@���\����YΈd�P�6�;�#��a�B���/G<;�̕��l�l�DTyJ�|�ޥZ
�\\�B2+ї76V�1_e;c�lې�S���ƫ�wS��t�(r��{� a�ז;�}�9ɛ�Cx��N�LSA�US�Q�g�yq�i|l�{�OBfW��R,��&�3��{�@&�Ww]��$a�P_OEqA�}%��!6�*.����]��R���Ǌ�U5#��/Ȓ���Tث�QP�r����[��߲��N�����nq�Ic���Z2cpv(ޓj�&Z�����qe�RIg��u�dL�����'빵AE,��,A��*c�z��+�FG�(�B>��(�Uwʀ�؟�\V�qK|��$�~4C�Ge)�{�g�<��n�f&bګ�зi�T�jK�K�y~kFhF�娠�-
��ߋ�s���S���g" ��K�QC]�<���K������fY5V�	Qn��_w�t�:c����f �Da󞯜�>�@�J�)g"�4��>Ȁȓ$����
��ik>O/�>Y��>D�zIS�)� 7����'�ٞ��χ}�q�T">��H�N;4:�
?&�"��8|>q���A�K�>�~�2���"�}��E��YG�����u;Qcn�����F&f��l��I��}��޹��y}F�2����E����M�n-d�G�߫�{Y��Ȣ���NA~ n?����zG[� 3$
��uݑg�T��b�+Z����о2��ݥ�0V��x�&bg�|-i�o�>ϔ�H7�J>�|������7�����k��͋�1Bᕴ�M
��ߦ�w���F��c��5^+}���Ƣ=g�p���Ǚ	Ğ>h�������Lg�UKP3�����[���tmm��I� R�㵏������Y�vb�ҬݫY��m�E������]��絭5�UZ^�L��\V8���ko]<�p\��y�s��[lG��M\3����dl����nu:ݍ>�/Rgb��UѰ\m��,���������Uۂ�J]��1{,̃WMF�m`]�M�`�fvF�X+qͤ@�Xla���Kr�[�(��b%�5���_����-v�.u�sv�l�^М� ��n��24n��%]�Xe�.�]�և�.=�B�|��6Y�m-˞P� ����I�z��#;�ǭ��������r�����*%��y�hK�����k(�p�št϶�f�L��_�jE"��HdDǾ!���dwB�\��Y��؛���D�|�"N��������#�>2|��f��H��g-�u�:�D����x�6I�O���bH� ���>�� N�##�E�r>��G��G�gϷ�����?}7���<���r,��j7^xfS\Ԣ���ޚ��R�<@���?w�coTu�|A)���1l��L;5ܪؚ��wL��J.y��
���υ��dg�t�����r(�V�DADI�G�'~����w���g�����}�u�ȉ;���l&����{Ƴ�x�^(S��Z1k�����}�[X�,���g.�M����80��L���6=���9������m�@)P�W���Κ\3����f�.i�ʄ1���]3��x�o�A�A�&>n/���D���φ ,�D�&Hߠ)�
�b��"Y k���n�p�����iC��z{>&�O݂���]�>"����}0.~����2piu�N|Ǭ�D�=1DJ�Q���.o��?^`w�u�b��ܰ��81k_���4m�?m�j>�.ڛ�(�#�.̪����A����]e�-��@�#��Ԛ���f��	���C��k#4Wf�R�`��O�~�_�{�TE�B���YF@�Hn �|>����}��K�`�c3ʵ,���q�s�Ҫ� ٘�4���mG� _�뽶/�O����8��<&c��5L�y�'������|T�q��d2�B���
#O����L$��g˥���A�L3*�#c�`މ��N.)C���<;�jk��v��PTТz��˺���tÇ%��!�����AU�����EӶ�!?4|�y�m�.��*��RfƄ
w���hB����n4W���@�k���bm�^0(�wR����l���$
�j'u˃ef�~�?3�h��������#�[%v�t��&�AZbm���$�$�a���B��dYzO�hѻ!p8�>k����q��67���-���?| ������&�'!�Dݬ��Q��h鲜6g�N���[ �s�{D�P� >�t� ��H�M�أ �����]r�
:T�Im'�6:b�����F�}��v���[��S4�	#'�Ż~�5��ـG�*P"�}eA����{3�P��t �p!d����g��\U��'��%�H�#�f����p؍���o�2+J㵎B�q�h:ض-	B��`���_�yw�6/�^i�l[-�w\0�7��{;�g���R}6��qD"A-�1ߏ��蘃�{mPA���f�m��n1���t�i��܋F����y��#L@F�rX�b?w����ڻ���n)5tD ;%�Tɺ�v-����N��<�7+�9V{9ڳ�H/U�I-��о0���b��x��̚���Y�o�B�`&ءD�;r�W�齈`�  ����"�� ���q�[�{�/Y�v�-u��&�m-s{�5��8 u��0�}�hϧњ9 9��������:���%�����0L@-6! F�;膾� Q����|���FWX��& �/�l(�c�9�{��~�L�?6�0m�O7y�|���X4c��4��2!����s�����|���d�z��篼~��|�ƄG�\_o�� d�+��r�lu��`�  ���F������is���Ʀ�!t�o"7n�n`�o}�ق>�I@0d���@ȇ�BgJ��ﭙB���2�����F�n�l��07h��3�0-��3+�#�i�u�N�W����%A�;	����;��!���>葰�	�U�I���FN�Z�ofL���Z�GJ`s�zi�ֿ_��5��n8��;"�O�������.��)Wqkmu��z�]I������Y ��yM�z��)���r�������ˬ؟$Т2PM�φ�����+[�������Dr�B�������}�� �vqik��Bo ����~V���㲻f�o�zc¶#�Z;Ɨ�kG	�_�r������G��*HE>�Z랆Ï��|G�{�_�_44�z!�Z3G6����<��.�|c�k���05�#ٱS�����2y�����A���O�������s�ri~�&� ���b��k�wE�#�^�^ ��*X鹠h+%䴬�]-�#U�QIe�#�A��4aX4d �O������s�Q�i ���� � ۻ��������p�� �@�H�H?;ߕz�'��^N�a�˷�����P�&��C�~�����E�� �`z��]mM�����#�2J�ێ�-�L��y���D� +����e�x>�TA�A�f��?��|G�m3e�DT�b�E�
�	��6����ML���n~�ޞ3�fQ����W��A����|�' Y���U��沲HD%@# �Ui~��U�F�*����|aѡz����lcBй���{��s}�<h_�'*�f�������s�
vK��&��.z���(�S�Q�賥.�ϻ�9��ؘ��!�:a����Ϻob$T��D��� ��tZ���ة��l�}w��H;r�[j��r�����:%���_��:u-�$Vv���9�$�BZ���x)�1��W���� _޴�=6.�B���T_Oԍ�}g�D(�2͔t�j��>���F�=(����#b�0�X��3�l�Ff��ƅ�m��ջ:o2@:p���^m�2�T�ۉ��r;큅@ޯ޻͠803��ZM	�M�b}���?�V��H��|���6%�g�i]{�Q�;�M��Z�VĊ�GK+>�U�B�ߎ��ڙ
 �$�\��}D*�r�ӯ�����,��>kF��)�Q�k���t�����(�h�p�Z�Ǝ���������/��#=z�������OYU}�<�s@����oWF��i�h���fI܆Ú�@�8����Lzp������&�G��0�B�7� �s��[0\(1!G���j|-���n��{r�D���Ͱ3�b$�F�=�~�U�(�Fdd�00��4\������mz��J�M�]-\:0/�B��A�����Kb��h�֏�b���^o�5*�K� ��
�q�EǊ��1oMlLi�_��qpm���]���J���ъN~�qok���x[;����9�$p?D�$�l�d�R�duYm��8a��EE��T|f=����}N@�v�h��Mw��A&�O��Q7t��d���1�H=���@���!U���>��(���	�i}��-��(�np�h����ݕ7�Os�۰���`��6�2I2~�Dd�bA��6�띊�q�G$���遟?~����+�1� �(���Ǚ�Z�ܪ� ��}s
�@Gvq����~�w�Q�Ǜ]u�|L5��El [wՙ�@�F�D�!x~K�c:O'螼u	�y�s�;�LT����k�x���gZ��u��	Il��#��P�a妖���kF���&j��SHI�h�����������T�w�d�$A��D�0(�Tm��w���ܞF���b�P������vkgL}`����-�)�� z7�}=��ؚD���r&�Td�R�6��{�N`���.��6��X�N{�L�ۇ\��$;��"���V�K�1�b�h���80�=u�)g��N޵،ˉl�)a�F�:m�#�m����,��e�]n�؀��u,��Ha6��Ǝ��������Mak�iSlsm*IHA�s���uss�k,9s�F�[::��َ q�\��R�䶩X��ҭ�����db�7A�lu�C�ׇa^ `C�c��v6n|��xL�:����赌΄�c�*����=�C�}w[j��^�.7a{����ţ[@ܩ��g��R&�\�"������[�QC2�	���ǿ�6mm �0���v�$s�J��s��9�]��}x��a�0I�T��"� ���\�`[:�N4���šo�ߍ-/�æ4)\�sM{l3a�߷��T�F�a-����W蘵�����`�~}|�}f���p�\�a�O�_��q���.~���Z�����6�8ؐ�I�G�?r�qi(p�-!֘y�\���n��4$Y�؀bV�I#�67ύ5ד�Z2�5��&�{U�V�$-��#���t`�S�߉���|�i��QġHK�N+B�j�=ߔὋ�����s������y��?_s���AwNޛ�gFC�8�	0����ͮ .��!�j�0�ЁR�Q4�K��~u��:�����8���nE�6hGo���z�i[�x`�����Ъ a�E�}k�)�[F��ܛŸ���!m�$��`hZ>�-�߻�����V��x��?����nZ2���9���R,��`6��D�k[�f��j��.~V�����7hobG�qEL�g~�;���"�:7?D��AZW��A�E�!$GX�7��0̪�G�Љ��"cZ3�DJ�59����@��"�S�pbbиU[?~�]����A s���[��q�c1���k�}?~o5���v��Gm�����lQ�M�#y,��ޥ^]nh92	�m�#֖62h�V7[���/�4H��0M@�g��k�-��� |o���� I��rA��a$vV1 �ICi2$��]�2	�\pe���w��}j.��D� �ɡhB.�s�P͜��rA"��$��~���!&X-]�6�����}��{K�`� (�$��:�P>y��8�|�韸���!׋�AŖ'�%�օpla*[�˲�[�W𐗷sunZ��s��h�Oc	�`cا.'9���#� �������/߾�� m���
��5~�٬�0(I�A(�"K$���9�O��X�;)}J�}�
��@A
���� �P�[5� ���ڀm� ��PE7�~C���D�ҕ�\�O�����M�w��:�7��M���<&�0��ޘk�O��}����苴+f��>��#9������3CU���޽l5dL٨� (�k�چ�������k��U�ϟ,����X}�"�;�`����h�
��z*���ـF�cm1 ������[1�U�G>�Й��FL�_~{���ء[T�4�D�_���O������_w�Z[��֙�kQ� ��3
4 m�F��?V��8���x]����0�O�0��b��O�~����<L9�%3c��(�a���|x�4i��-��b�#~۪U�$�����������>���mmo���hB �$��Z 8ٟ�I�(}���k��E/<c�!�Є�I�F��w_Q�����h�{F' �+S��n�1 �ŝ^x�\��WgOB��β`g�`��t�-؎i���� ��W��P'�>�e��?F>�צ����CM�~����孜o	�{ZBm����k{kXxg��#b?~�?=�����ѽ�Ϛb�	D�`0���7�ƙ�?�@b�ٓ�tzl�9�=��B���jvYf�g�"���6�� }��<�$�_F}�}��"�ML}���I=�6� #���ב_�3߽�����{�ߍ �f����=��_ܚ�u�����m���֚u�؄��T�~��vi-�р!s\{�?��v�#�ϐ��`���~�^��V�[k�v��#<>lMi�@�dl@�##C��߿M��ip'�<`}p�$�#�>�eeo�;-o�p����.o�|9�^�:���eL�7"##�i�ŗ�^
�ū�����P��2ֽwR���V�X�I,��y��柕n�X$����c�0�Ϗ�܈��ʭЌ����m�F00�`��s0H�N˜���n'�I��&f�j(w��J��8B��7�B��̼�b��	ٸ�����gģɁ��ۺ6u��ݛ9����-���2��������	u|�'M�ne����ճL�s�	J^��$a��"a8�;�$��/��}�Fw�"#iu���,(�v���f����V1j�;����,e,�1��1Q���i�o���ң������_A�*s�F7uz�K��I3ŦR��aٺ�X�t�u��9\�:c��x�ၳ�e�`]0�,����Y��MԠ��&�",���	��N�|j�l:�C����89nj�on!�qqiZ���ҫ�S|hV�h޻�q%$ �dei�����U�0�O5�[��op�*(V��ued��n��ଽ����7���nX=�����x�(�[9m��Lm���j�e�4�J�gj�:�Ӣi��nf�$\�fn��]z�Q��5t���Ln���|��a��·9��U��gs��#��8$��Y.v��v�c[h���&��PR��i�a]�ws�V&Lv��
=��o��"��(��o��w$ �P�[��&\�Oo���J*�����
W9c�L��̼��[��"��1d���0�����o�d=���X`�Nd=۔WJN���ͭ���^J#�Y+qK���;s��M�x�A@b_�rkh����a����3�n&
6�o���ќ���7��O8	j��6�Z���L0�rϾ��j�-갮YհB�š���5����9�kZ-� m�[���� l���"=F����-�`-6�N~�.�� �u�� �@�8�@�-4���-óSO�� @��/�����X�y&Jm�y0#ĂI���TM��P�4^0M�����ƀ#�{l�
�$�[#c��h q�	����ڊ�_o�뭨�u�m��Ǹ�q�4`
�IϿ$�t��~ﻄ�Ȃ~��ڈx��B�4|!�4��v #���[@|?7�� 6�l@i�#�kM�b������G֕>���`y�F�c Z���ߵ�ێm���No'm������w�9x![5����h�U����H6�n
UYU��F3�$�
�F��m�`!
�����t/���[� /6�� x�_�5S�����4�aZg������i�nD�M�����A/ߵ����׸�޿�����5��k��`*�sk֋��B���[&��q� m�5(ŭH� F����5`XVR2KV�� ��` ���nE��6�cޮ����`�������\B�i�P$�H1����m���T>�����̀1���A A�l ��:�j���n�j7����oI� �y7�p6�&� `a�n0g����kx ta�I7�������V�v��$�>I��ā Лh4�a�w�J����2堬�վ `$��A�� Zi�B4� A����k��[@��dQ�e� A����H>��ۚ[@���0��`~�����˜�N�~!F� `b8:3����{f]�z0�3M�ЀQ��+��LADϿs�[��!������ 
�B����]_���n5�bxӒ��C��ؕ3(�����]�_b� �>����  ax@�b[���׋KB�uȳ���TY.�������Dw@��YtUq'����W{v�!CW�9������ޖ^Z*��θ�9Oz�����⯱�3F���OA֖c=�v�юx
>+schg��@��}��b�I��I�,6Sj������e�|i*,|y���%��2	F�dGLb�m��������T����ʉx�k5��[3�t��q8`p�b�K���f�����Kȃ3�y��E�_ur�?j}~�R����n$R60�W;��qj�P�l���G��kư���[��yp����eE�TYW���h�g�J���U_>��-��k-iI� ���|������(bФx�!��/O>�"�ȩ�Ӱ�m��n��,��
ÍC3}��Z[�L�b�bLKb~�[-�<<��``,��3����5�Q�F� �$�>��) Q��YU� 2@����Mgk� ]��}d2,��7ﶵ�G�1$�♔�e��b����.��3�zg���F$�L�ϓ��l���X�f��&(fd/��i%�s�ƅ�#b���$�[�>��)G�j'�E��8�98"�v���W�� �ad�fsv���u��V��͜<x�u��,��8��lmȪ���-Dr�Q�Έ 2<K<!WS��o&%��� z�D�� Q}d n��<޶<�'�z�o|���x��4Ĵ��г5.�$i����:|>kv�'dVw�\BJ[��l��y�|,�fw�ۛ�������if�阠�E$����_qk1q30��M�=�������z��ZY���,����h؁(.j�{�f-�u����j�ģk01/�ޟ���
��.q���f];!N맳���h��6�vL���.��r�Ŋ�;���&!�Ԏcv����Cy6J��v�~WӦ�馆����@�B�V�$�H��EF�2f6lX^8&�h=��1��F�/D��c���8�hh`P*��,��q
E��ٍ��c"�6�����#`]H-gG2��1gX:^�;���ls�����1;A�[\�#(k���[�"�Wu46%iH-B�jg�K�DƮĮ�-�Y�Þݗ[7�j:D.�u�O#�7 l�F���>it�-�n��۱�!m�
�J��5n��<d�n:���a�g�����~����;td���Q�n�+������Y�H134&,����љ����{�\���hK��y�����}4�f&b����b�� ��޳Ykg�eT�7I�S'<$��}"�{̒��l�@���#�}�D��ϲ25�	?|&�GX8B�נX�f.�0<����Z�G0�!�������,�pTI_w�ZX�8d�@�q5 �B�D����k���ȕt �<�qvo�H�,�&��jʻ�bZ1A�1'��Qq 합H�-��.F�&b�4�i-k_ik3b,#���� ϱ���C÷f�����9�?t\9��b]��2��ib�y�X��_m�+����w�gL]1k���^M#d��?{��H��gdd�(�!ȥ����q�kko��˧�'�@�$I��>��>�U}3X��%�(����">��Z����Ŕ���C��xX*lo@y�&H�&,شfQ%�m?,VF��2[^�-��j�S{栩��x9�r=D2<�z0ĒG�Aˮ��{t�[�kqH�>�"(���� �쵬[��<^3�\O��&-f������{�i��b{i��$����PK>��f���7F_*��'r|r*62Ja��^`�V�fyQ�wn9��t�(&n�L��f�:9��V�b�iUI>Y7����$�Ώ�s�Ж��kU��K`-���%�>��Lf\x��c35wn}﹥#ҕΘ��2/`.�!G��r�Vl�W\*g�����6���:i%��鋽N�bZ�h���#ďY6�l��s�2e]l��*�v�1���Mܙ�
�uN�e��\����co^��I�q�#U�c�n��Y��Z3����w�Z��1M�p3D1.��}5��]35����ǲ,�@Gg{T�$��ކ�����Ntĩ�TĽ�u=෈�;ۗ$
 \R������'�@�K��ϡ8�����}Ɠ�� ���&���t`*/T���S�%�ncjW�O� A������oP���H}R�l���Ȉ���Q����_I0�:MWxH�,�޵>�4|d�-��B/<�__��pCy��L�i/��>�gȉz��(���F��nuǠ�Ku|$>@T�D2�Ñ���'�0j"��٬ٛ4e1w]QQd����͊�EMj��pX������a���z=�xO��1�y�*�XF�w�ǳ�tNiY>& ��5�7�f/D҈O�ŝjp�y�����kYe�Yj�Q�\F-M�\�H�m�Y[�����R]ם�.M�9ܛ���o8��Ix���,�;�${C̍��g�I�>�r�2�G���!�����'73sF8껭QE)^��&Nf��kIl��U������^/~7��hř���������y�%�5=Dx�����x��� ���f���j|2��$�>g�"A��H�=gȂo`y�g�r�w�$ ׋>�n��{�\3�����ί�Z�8��8Kk�D�b�ct�,
(C l�R�}��s1�" �B�����U:i���F�u�Fue����<���ԅ���t��:��2tYh�+Zt�[�V�׺���V���:E��Ɋ�Sk<ϸ��r�t��c�С�QC3]�Il��'�M6�?v߰|ASpZ\)稀�Dx��M���ڙ����Y�b�8�dI� ;���
1��D����emS(�b��[5������$����r��#4� tvڪ��|	����/��m�;���*�۬��%�2�o�/����T���h�D��d���Xi�B��u�`��o�`A���S�q/oZ�i#|Xu��*[z��uۑ��� �>D�� @G�N�� ���͢K?K��\�D�Ge�0M)�C��e-�7<�[�<�����̌�^�ٵ7j����M<ؖ��}�w���,��0O����M���d	Q���=����*1�x�|��ч��&f�Y��s5��p�Ό�+����>�ߤ�NɃ��`�4�3��ط�`ɢ �|4�SJ@�7�Tg2��;��dD�� Fφl��=�$	>'ڠ��Q9�J}���y:�L�[��U���3K!Z�U���< ��YF��{O�dN�+^7Gl�鋦�ۯ@� 2-�ڑo-�>Ch!�1"���5���� A=�M[�[3�-s��ҍ���!��t�I��{��,��9��n�Y@ځ�b�u�>��	+���r�t��3*�|���!���h���,	�1�@
� �fs�#Ơz[�GN�\���G����'6ɓt��F�Șw���ن����.�+��vD!�۹�ݹH��K���詶Pw��c�{v����`��S#w*��x�Zf��s*7v����8l�����@��;_��%��4��X�X+<�z�-�T�\��w祛=[�[��ڠٗ��e���Y��f=� ��sR}�<
"��BJ�G�c6k����H��ޚ�w�!����n���q�^܃��mϫ	`gl��A�鶱���slͭ�h9��.�'�'����#��L�Ʒ�[�>ɪbH�lE�Pv#˦k�{.DE�"�pHEl{s����ɉ�����\x"4Dl�]bƛ=SC�T�$�d	���)2ȣ)$�[2u����h�lI�^�S^35�X���mc��*4yD8�g�B=}2$�ee�&�>��zb�>�XE�/)h"L�R@z�"})�YA��0v��vđݨ��|	�>�ݍ�P�T(��Ϟr�}�R*�. �>�" �t��w��7�+f<ݲO�y�U"�@>$�ѝ���}]�����K�[�C>]d,U`�n^Ta���َ�����a�n�lH����1�0ppܙ���BH�G�Ő�� :�;Y
�1�
&"�{-�ۣnˈ���ZH��Ċ�C1F��UBт'�r|�maejF9^�l�}�V����֖����Ϟ��Q��3�'���{0(�D�۟�M��̽����	C�B��!�w�I����C�G�Q����{%�ud+EW
�1�F��^rKr�靍)�g&d��FoV����3u�m��oƝL�	��'SF����+�����Str[�3[�>l$�p"���*ں����F���8�u�L]�Ƀם��eҊ9댙�[N��a�;Cjlq��g�ɓ��;N�.9�	^�Q�W7�!#]	B������;�#j�+hl��
lr�seѦ�u�V���|����(6���12Dm�lu� ��r��3��p�s��n1c�o�Zݑ\�y�uas��S�Aڛ�n�-ۛz���PM���[��,֞y�!t�l��ô���h6�Q��I���틡	���]>��zM|� E<߾t,X��1Ǹn=$�!{����M� K�ŨO���A�XF�R3g=�����_���6.D��%�xEX�52��H�ۡB��
5���[��$ѢDWV+U�50fh� -�!}U��9i��B��]Б�z�E�,	�g̊�
}����A;[���wf3أ��7"2�}���v
X&�Nڶ����H {`F�ɚ ���8�L�}gH��B$FZD�1x�j��j�f�o�"	��>��a�d�#g����Dz�g��h��x����$C��վ	1,��G�W�����G�DT�B�eb�km]w�].{�2��( &ƙ=��'rd2p�>ۜ�P��2�ٸ�����R�3�/�Oz]8D�»Y���j�*<O����ԋ3X���ϕ���[��5�y�����Q�xϡ�� D����L���q�6R L�P>������6||L�q6�v��U|��r[ne���t�ݸe���F�6$��ЗMhˌKXa?I���#?�'yg���v��m�2���h��������#m���L��,�kz�lwO����(eP�� �;(29��2r�M�,��q�t�G^t >��(�KUy$��;b��A�&���o��u)�L@p�pqkkҵ>'�;+��K�(��.Py���3���������ⲎP�I*���r�;ncD�ʍ8�I����i�%2=}�il�ݔ輯��S[�������>��b6�8ܔg���4�L�3{����	j��٢�NE�}�[D�ښ"�A��uBu&`�#Q�/��䊢 ��P������B$�KH�^��>��ᱪ����F|�7�Pl��t�B�5o�X$�ѝ,�	:E]�	 V)�$�A�O�̳���$�;��	-}37�yt�1s^�=PQ_|��٨TV����Y�ػ�s>���<�X�9N!�,3wۚ�.'�t:��^��l�e�Tف]r*�E鉰���`�HG�T��*ɰ��HI��\�;� k�F�l����V9�Z@���l#
��9Y���vvm��&���E��(k��b���k�~����A���މl��|m�	'z��𲈬3�Q�,�L�s�$F�Ï��G�e/h���:�X���� �}�}��UʥCN�9M�Aw�F���;\ējzkk�z��'����uկEz���I�@���n�������39���V��*�����ٝ{^b�GEJ�[��sS��@�ڍ�V}��!L$��]�"r��`�bݭ
I�:N1њ��or��J�c�@i��)\�eK�X�H��۔�nv�͖��#��Ǝ� ��TRD�(��5��soH��	�68����	��V��[,��pbK�T���P���LNDålY�A��U�LT���<�l}����&�rWkFӋ.{ �N��oV��̜Lp-'�6Jl$�a�UGF-�jYr�A��)�X���l��]{�J.vd��:d� A݄Y20�U��X����X�z��Bp2�M�w���{�N����u�P+ʝwWy4Ib�Ά��0��rX��Z�9kZ��sz�b�!��-]5���Y�?�<~�<�`����՘����%O���_��U=b��M�[pYm$s)�~��ד�e������2Hm��e�����m܈"��d�[��������^��v��x%�W_=�3�۵2(�ҽ7;��EҘ�Ȃ+�ЈlD0�p�p�mU},u%:�&���P	�|��A��GE�NJ�N���k�I�Lp��D��!N��c��)���c���|R�l�A�ݵo`�|��C���<�N�3��`�<�%K?��U֥u}ir�r���
3VE�6n��C�\�C�%n��M[�b�ed-�!oc}���U�{/��i��-�E"KFm;�C�:��a��e:]Z%g��[��KQߪk��Q�˅���hQ�k
���&jx�.��
�f��N�EW-��5���
�%g���T-�**<�0$�o�1aA^w9�۔6��-u��\�=\<c\`Ǹ��nی8�D)#��X�X�d]��l��:��֓��8s�_���N
���˓���]�5[�����m���Ր{]棗ٽ3�1H��i��-&�Tb�/�WnġUn�. �o�R�GHA,���䲠l�) S�&z�YA��v���l�"h��	1#���L�ཱུLD=���B=�'�wu� �Wݾס����t/.]�j��;���dQ?*�,e��KMU�<��]`�.+�|�&Q�]�$^�4��6�˲��G�`�F*���ƣ[��f�G=Ee��(�枨����`j�R����[LI'�ȃuozޅ�&M8��ӻ�`�_�3�ř�환�f,���,�K3f�fbY��1�f%��3?�fbY��3���K3f�fbY��3�ff%��3?��1,�Y��9��fb�����K3f|�ĳ1fgٙ�fb�Ǚ��f,��,�K3f�fbY��3�ff%��3?�fbY��3�f%��3?�fbY��3��3�ř���K3f��d�Mf�n����f�A@��̟\��o��C� � m� @�PQB�J �h�@
   kBJP UP(�� �H  �B��_                        �@           h       M�˘V��/;�z �F�'��z7��נ����Z�o ���)C�`�z��Ex�S�37�[�70�=`��:SCR	� �QT{ezx�.1�r*��΀x���
P��    �       �{����J8 �P����q�RN6��s�N*��PF i*�cdT��� .v₤�⦱HP�΀     � P�ԧ���������1R����(�X��Jn p����D� �� 4]����fm��� ��
Y��m�v�P
* ���� iN����=(��< :護��<@ b�B��)��(D�hPX `�Z���:kE��y�^s��iLCW0 �����E+�         s�
K�ͺ$���HJ��,��0�厀Mb8 (���nnt�$��	ِ94� �b;�=k����E@	 
@\Z�P�]�t�
� Ϋ(��n�R��͝�EG\�kB�M2�p 8ӵ�K�H*��*��**s�ld�h�(
 �� z      u"���E#�\���s�����.ڊ�� ؐ�Y۔��^���';�R�#��J�� �A)��"�Ö�@T�@�]�h�)M�u)�d� �	�I틌5�q�PE���(� ��;�;iE�2B(�`�D*��QU�hT�U
R�         �J]�%J�`둲��""ź4��� �(�1���\�$�3vR[��*�� ���L�9��ۍ�T���.�V�4z<�'y��i�M� �� ��JKs�^j�))r5��N��Sy��Qx���ru�ڥB�X� ��$�ͮ͌�%D��RW,�	�s�I^L��a�EJ� �?L�R� ��d�R��@1��&� '��J�z�	���5O�$
�M��d` I�@��5)l#36.�0�ى"�����<� jBHtx�9�W]�n�c��@ �$�
� !	%��BC� I?� ����!$d �HHO����W���+@�֌�~���;��@�ᛘL-�[����̽�2��Pe���𥚮��-���`���W��b��y��`{35��?�L:���q�h�gll�e�ү#w�3�B.��_]�e�2i�J�W��v��[t���a��ք���-�e@�ۭr!�we�eCw$��!!m༞�;�G<#FM���ccJ�Ƕ���)�z�"�P9��"+c�e��a�VQ}�u^
N`ݦҙuY:�j�'���1)bA�6�!+��⸭/C��T��;�1S8�Z;6dt�-1 ���J����S�������;�va��ͼb��ڼ�c9cS��f��	w[4�bڠ&#{����c�e `�q�E^Sѷqk�^K��,Q:��e����\
=���3{��j�-�Քԭ�.��ۋP��MLϥeÁ� ���va6�͒�FQ!В\�f|��3p��"�WMC�r����'������+f��ָ���]�IrP��a90[V��X�^��)Ⴏ�dP܂ͤ�Q5t-�p�����ܢ䒎`T�rK�ۏZpP��Z��'zYx��Vi�V�S�r��A��B1�͊m�}y��d�R�a�&�F��vq�V��0� �m�F����o�R��᫸l��Cr���J�X۹4��@a�(d����$��.��y5��2˹&��1�jcN]И�ICaZ��id���j��N擔nՊ��͟>mV�B�mR
f�uz�lj���P#�m���dF%�5L�37�u��/���j�a��)���xj�E����ʛ;�*Z��wn o�&��\�y��׺�a}s+�3h�{߼�d������M�O��~�,lQ�����yl+܃��Ʉ�_���� i~i`��)���Ws%`�@�WL�Y%i8Q���XTi���[?9TF�0I��6#m��M�*�Θ7e��G/��T��}&V*���^5��+3&V=�38wCm!.��"�t1VB���%�3*B��<Sׅ[qe^:H�˕�	y�6ڹ�wJ�\��K�R�ͺ8�n�ɐ}.c:*觡�hO��
h�ٙd�D`�q�����
��A�
M������޳k7
���*�e�Y��b'nV�pE��-c3��Sw�h��^��b�%��a�f���V�mDSf�kʛBj�������cQ�i϶��ɐ�ӻ� 6���un�Q�R�h��8��6��"���A�>n�yW��R�ך֗@f]�bٵI���f�榠�5{��2��ۣ�/sPr�b	t��#0��`e�m0�P�c*��v��4��o�']�x��;�2�;M���$�b�9�WC-�wOL%��+j@m�R�+!5b����؍"��7B'[E�5�Q��y�'���T�0�6��x�^�	�f��c����Z
b6vfU�e�F�CJ�L�JZ�����^��V��"�J�ʙ��l�����F�j���n��ml�Q� ַ��pGP#�6��\���C�R��r	pGv�b2)���R�����wF��1�g%�pX]�j%�`ݘ'�F,��h��z�2����
W�	��c\1�z���(*�"��h�~�]���X�w D�W�l �7��Y��sk�����f����3h<7,�je\/�6������	a\�oj�n� Ʃ=��B��VN�&��9���S�$Y�P�
hQ8h�b�7-mk��|� =�G��嶎% 7B���8Ә ���H���c�P�DQ&�ci|[L���i^��#(�{���X���O)(MGi"�:�0�V�pl����e�,�x~��O8���Sw>��r�Ц�z�KX�8e��MC
f�]�1���Z�b�mV��ݼ!^��.<��sYRZ�k6�*�N��#�cy�5R�V��47��N��C��C�6\���Y^Zf�����y8زU�%��ūfC,`�3NҵP��Ҙ�c4��$�gP��zn�+��F�L�n��<^�t�x�\pE ò�fc���.�7YC2ޫ`J���r�ѽ3cܖ��[��&�.f�j�R�:�!��^����ߪ�{��G�!Fn�Q[$'%�Z�_tp��(S�/O���T'�ѷ�N|��p�[̃nd��
���@f�=f�X��c�{ .͋U&!� �Lܰ�BHlLr��+^6��&̉�Gr�]�պ�*�sV�wj��<O_T{}��廔����#B��ӫtVd�ᇬ��ݛo�ob�sVQ �b�$��0MqK���{�#Ѭ�^%�]�+�kVkWZ1��3F���E�\LoPVp�[��(K�%r�.;CLf��)�S�Y�h���Rk��:%���a!�wUAX����윺XeȫI�kU��� [�)ehb�rPQ�*��ʔf�m�f�j�n���m9�j�.� �,��MU*�PVƯt�]$э(]�����y[{Q�>T���.�R;�i����i�y�aQxJ��L�����6.�<������f`˸�W��d�t�R6+tI`�k5H囲�j6�;5>
�2�!e-�r�6Y
x�	�Z%�v��7�R��46X�b�M��CHE����S�i�����0/���a�x�pO��o-���n��]]i���Ԡs�a�z��%��B��Tt��JV�s6Y�i���h���̅Zy ���fp��n�%WDX�ykhL�e歭8޼!���/-�ǻ�ڦ�P����{s�㨮S:p3{S(��(�:�4�-�si�6�F���w�z�X+0���c��-���"�R�^�PZ�(a��Z���RUv��	�a����O!���W��;XZ��
i�X3Z�.%WL.���X
�J"-�� �ۡKl��Yt�5��j���i����mּ�wu���1��Y���OR��,�xT@��d,��HA�.�l�U����ֹX���Ptt,$5���h�LzJW{i�@�3/	X����v�Iu��D�Lڷ����Ŷ�b��%b����ԥ�ea�������Z�R{]c1�v/�i�������fL�ll�ci|^$rEq]¯%�Z�b.���v��KFӒ��/�B�k�H��Ǆ���]�(QW,C��e2��Xm��m�������2�͂V��x�͑^Vn���Z` :Ea��W#��7N��e�������7s.*܊�KyQ��55�B��n4�d5p�4U��d�h��:��1H��6��������͓sUY8�5��nk��f��%hk1g�ܘv�X�<p�f�n�;�m'J���5�k��[5�َ�_��ǗYFA��n��AwQ�Cjm�*�Ui���Xʹ�!I;�u$��	2���Ō7u�
WyN��d9u7< �P<(�7�ܬ��V����B���ref D���j8�����om@�l�髴�)���
��Q��)Y�VܽSM�n[-�q|�e][yv�3M��t�e�{�iԱ+ĩ[m�w"_Gmdͼ���6�!��%�oo��̷�{i|����,���{�qSj�F����ˬ/�?^��ѷf��pF�f-�V�j�H]ʽl{��J�4}���+z��d���ں.��D�*�f5t%f�¬���uQ�����O����1� ��F^�a�30P�!Uu��)���h<{+-(�Xq���2�k~0�����os)�:읣i]R;��ܳ��W4*�¤۸̒=��Ƶ�'G.�fPRX+�
zj��,���I)HJ��"YY�$���/Pї<�v��M�����p�H�y/.�5�Y�f�1��Nꕊ6%�����ej��ǚ�2�@.V�߶��35Km+ɹ���h�ڳ��ZWX��$fJY�Ц��1��eF�E�ۢg/�Oi�L�܄�^�;V�*�Yw�R�5�XK9�
�x��~�׉�ia;t�];��	㫗t�ذad�DA����{ש�U�B�A�w�����eM�X2�T��MGk���l�����ҋ���i�+�4���>�A��
ۂ]�;��t�1������h��ˬ�1Kd�Ur,��8�,^��Y�Ŵ/r��gv�7.Z��ʎ��S/v)��V7�5��Y4p1��j�]��9*�Y�/(8$;(%oF �c˽W���d�`s1�[�$)����u��˼NI�V��Xj�߲fdn���H-`���@�mej�*aF�`Z�f�KU2Gw��(�N���)$Vdܧu���=Sr�V1��wv��:�+��s5��L�At#4l�n�Hd1��2�ܑ0�i�ZB%	SeP!�o#��k߲H
d����ʽS@U4M�l��c�Up�Z(]�Eމ��X��(!���unKt�����l�&���S�6X�>��j=W��tD8ʨA2����5�┕�o��L�����N�M�w���D�Bl�ɗ���2�� �:le`��AmfN��nU�ۅ�>6��
�4�)|�j��&@�<�!Xs-�z��T�s1��� �`�:��P��@&�ufX[͕�2����,���S+�*�����m'+a��`�T��O��Ʌ�4o��r�
'^/ٌ�62�Uxf0V�N%
�t3\ܡf�y��
sksE�w	ۚ�e�ہ]c�u��4��m��#RʘԒm��n�b>xk,55�[v��yu0@mYjl��S#m�6Ռo������R�7n��k�z�jM){����;W�t4m��&T��������n���RTrF���ޚn��n���ز^�sDg~/*+DE<�k%]�[��ʡ�N,P}j�m̔���X(M�T��Yvhfl��Tl�,ޚe�CD�E޽����aO��nS ��e۠E�����ٮ^ވL)�n��&M�;{G�͹Vrn�o�
�W��P��CE<M���J�-���-���ֳ��Q�e+��m�w���Kλ��y�Ȝ-J�k7hZ�cs.�/&���f q�qz����RCq<�+!�Ћ`]K���r�c\L�6f��EM9��"���fKi�4d�i*cE��YG*C�N��Ja�=u�`v
O�b�U�oֲ�~�oMf�̠$�@�I�Y���-۩�V��z��x��3���K���6��CHf!�.X,�!K4˔�aL�j�%��:�B�T�;Q��ˁR0���ӕ�%6�ؐ�&ݲof�Q��7-�����*���ke���ݧSmb��Z�u�Un�J��x�6d����̬��Z�`6r�ڸkFi;�[�h`o��4
�i��k:y�\���ܧ�����.�K&�ђ\ٻJ��6�Y�rn��4`�b�ۣe#j)��d&6J��6� l���t�+5���V�4�x���� =ەw&
�,�sj�E���-�EZ�u�ۗl0�}�f�[3(�Q�@�9%-�M�>uHX�l
LšDP�v�j����ʳ5&D(8n؍V�qդj�J�B���o�lg���ٖ+/6�]�!P@��Ԍ:��Y�kB�vD��dqDT��襁�-�Q�fcݗe[fʻ�V�:4�p��2�ͳ�I���xI�&Vu��ֵ#� ;`�:��^Fv�ћɛ�W�.h�����F�NlF�7*	���̸w*&I�7	4�˦�;d�eJ��*���Z�8��ʗ��˺�����'��x/Y�6����X>�K�l�C3�3P�oB]�mm�W٭K�q��`���*]˛M�7N�@�u��fM�C�f�K���Eɛ�;Y2��v�Y�QD�� �WnB]MP���y��ٱS�Z��wf�IZoA���o~�1��O.�`g5��U,ѯV	p,T�n�Ѻf�[���
O�.;݊�p醳T[1���ՙ��A�;��O3���?!#�J����9t�1委j�Q8m�zkP�u�K7��e�q1����@skrG�Id��:74�lu3*j�wp��:Kv��!j`����]ڸcB��	9�uz��	��n]��ǵ��FY{j��b�};����c+�V.��s2@�h���Nݘw-���RM�P)$hJ��<ܠ��^S��(K�,ٮ�ײ�VS&ӸB',�C�lr��h;�3m�eV��z�^1��w1�
 �B�zY2�n��L
�sZA"��D�j],�.��gY��wv5,IH�m�2Z���� �J�iZ�SH�We�Tu��2�GH;��e��f� %94=v�g�
�U.����X�Y��*h(�iZw�Y9���	�ȼU���i �ʩGCBbWWxdج�k`9N[&���0;/ ��/4Q�p�����R���P�\vsf�Y,�B��L ��*�_ 8���):���#��T���f\ȼM��Y�*[��u<�0FT?���ϪX�&�t���F�+#��GM��|�j�yRz1�ܴ[�+1�� �D�{P)�{f�kV/�Pآ��O(,4�ɕ�n�̹ۢ�-Yܽ"B[pE�7���B�&ŀ�نb�5�[�;cPc�b��ˣ�l,�&i/b[���$�R�ˠ\9g^��zP�9�B(�RC�j���zI���XȦ��v�*B�
hٮ;�ʈ��V�urD�{B�XN�p�T�<��:���W�is�175���E��ɒ��F�a¦(�U5KYxZȬ��f,��2̻����z��&��͂G�f���c�=g���} ����n,eLl]����,pn?��3%���퐝k�B�������zmCB�ɣq0�-�Y���|�R~�lxa?F/к�XZeec�M��܀�ͅڭ����(,�Ƕ�i@\�-CO�)�m��c�0�)�,t��_��?�bH"�~�F�FF��ڮ�m����e˧��˹�t��=K�佷o3�n�c޻m�-�lZty۪v�xzq���S�&3�۝��v�&�r��f�A�m�sgq�`N�8�3��u���V����_Y�c����8ޙ�|���z�Z�R��.��A�^1nv���7q��g���]^�n,����ֶ�q��k�����jl�㶲��4K��m�Ș�u���I|�����f��9n|t��Ze�� �Pu���{\�v�=����ncv���V�tt�1
^���W���n��]��;n{��^��Fzy�vm�K�ؽ�^d�ٞ� �6�i.�c�u��8�.�m��"�k.x�tv���D=p�&���+ZV�����^@ѝ�<]l�f���o���N6m�۱��l�[4�=��;=a�;���H��-t[<0�c	��q�Ps$�O�Mţr�S6O��W�g-��S�#��q�����m��w��u�وw��|�۱��-n7[wGvXm�Ν�]K{���7]mɣϑ�;���U�ݺ]]f��i�#;�sے��m����f6P�YC��1ǒJ�g ���	�C������.�t�v��Z�]r�\ݺuŻ7=�Mǒ���/l��L�e׋�"�еq��4v�8K�糮w��/N��;��v���rs��Uŷ�0��v��v����
F{[$��]�S���rm*�Z{rt�(;O)m�wh9�L�v�C�y{];��\�Ǖ؏1Cn��Wm�E9e��ӶkP�C�cˍ�u���ݛM=���ٗ�n^�s��,b�vQ�G'eܞ�l���E�=�=�^9S:�现v�U��$s�F�;�X ���pfT0�hw4�<��g]Y�;km���6���K';9��U��Tm��j��4�6�p�õcO��셻lv{pX��ܒ�#H��9Zm;W�������n͵Y���\ysH�N�L6�.M���	&�����1��g��k��R��x�m��^���v|��ѣ�`�<�a�n{��g����W�������ch�<�=)�D[k�����-�2v�.۞׭Þ�ͪx�]c��	��v�w��0��c�pU��v;;h�u���l�N��ϋqho|���z��Z�n8�7gtB���p��x3���ψ7<֣s��Lu��r��{uی��S�:�n��{t���ـ�D�8��װP�nО����h��^�����s��#��>�O'*�Ӷ�Ϯ���:e�Cɱr�:G���x!���.@�G!"\�(�3��#/G�۲+Ӡ��x�OX\c0�k���T�H�۴vKZ������a�/77:N�8�����j�ƗK�sgN�n�mue�j:�ո���ε���x���C�mj�N;[Z�Tp6��W���!r��m�۰8Ź��cmv��N��ck��)ǴO7�>���/b�<��N���`���@]�0h��� ^_F%�7/�C�1��8�������pm�����c�����S,$��Y8�	p�7nt���vݷ��^�ݱ��Usn���[�<�>��\��Q�c�v�SЫ����ٍTv��<�t��Q\=��8MT����;kF���r�aJ��9|��앍��Z��r�m]��O���Ջ���㧥���*װ�\%E�۲G9��o[[2����ݪ���x뱊��e��<�{\��s{tGE��%qo�u1v��k��Qڷ��'f:�N����ñv�P��)#���]r�v�N�ۃ6�T]<������>۱���ݗm�nyC�lst�*��UOb�iȝۮ۷��]d�D�D'�re�NX빧di�Փ���ʝ��d������ɵ�ny\�kqn7��yV3��7[�rtB:�s��l�mV�f:w g�P`�\g$p���ؘnܽ�Mn�nڣg���[��g�T���:ˁg�[[hvη<���m.�P��VVM��Ş�S���W<L��`�z�&������>�۸�\����iݶ�;���;}��׷��/����z���랖�1��;o�x�9��f�)�p]u�KV<�б�ysǍ+�^ͳ���F��K^�tc�[�w7�n�{vzܔ��X�hd����fy�y3= ���7j�]J���׶1�4C=�i��+���u�qOX�xьn\�c�r���@�c�8���\��pK����B�'�S�`����=G[Z��k2s���ú/1	����g�';m9b��.ֹ}띜�CcU�K��㰎��d������즸�4/n�Xݞ{v�j.�5�M=��
S��3�Q�����w8����t�y8�;��ly���r�1�b��v.��m;n�q;�9��nv�;qƒT��p�� ;ڶy�g�Cm�P���dwO[�-�&u�-���NQ{�5#���ql�n��H{� z7�M�x��1�)�p���}i0��j�.FӷS��	�O8��|����ol�m���)M���cM����ڰ�d�������{���1m�Mn�m���9�s�"��s�]X���di.I\k��<����n�=cg��T���h��D1o7�������'F��NLV�fŭ]��ۗn^��ڸ���������u�ر�������\��;�[����sq����4�*��Wk7:<��؈��}e��ƹ����ֱ��Ͳ�/����(dރv�򞣛���ݽc�����v]��on�v�����>�^�dT�e��#�[�&���7�;����{[�֌����5���˴j���-כ���{74�������������8칛�u[ڋ��N&��c��N�V�������t<���%��3:�S�q�Z'Ec=k��u{\x�y^�a�p�tJi�;uŅnU3\���Q5<�a�a��B=	�!�ړK%�ֹ� g��9���n4/���6���m�!nM=W�mn�us��N�z��nC��cWj���b*;x��-ݭ��z��ZIۇp�*dj�;�vq6ǫ�n��ݤ����Vqټ�^pv���S��h۱�,�g���qv��EÛ����������`��F��oE2���n7Gc���Lˌq�#f�m��9ݳmy
���>{uK�H{F�sї��N�u�G=������)�n�3���o}�����ex�.ۉ;^�ٝ����k�=�U������� ��v���Mч�u��WQ�g�B˱>�y�KV7�t��S3�WA�|�[�u��&]hW�w��o%�� X�^�r<�y�G#�!��)w;��L�e)W2��E����������7!����˺�d���H#���]�0���Dɯ2��ۥ����N�:�Zw$&�Xm�e+է��<n}s��ͼ��z��2�������q�_6�q�Qخl=D}}����Bn
� �	��3$mF��+\1���xŰ�g�b�#�mG]���v��o<u�fzt�;s>g�E �9���޳�wF틯L];���J�ɞ-oOa���]�ښO9���Qށ/��r]���5k���n�[�Ͱ�z��iJX�}l�Gn����pg���s"e��zp�k�mz���x���l�85t')^nt�<'Z�<e�Cv�=g�����a.�zL�=�TK,�l�v�NЏ�X��-��AڻD�\�`�W�t�
��u`�Mɗg���gc�{��G�׻.�v��\�tK�q�1�j���� �vݹ���v���g�B\닗���:�[Qg�9xu��͙��:��ն{\�����K<B�-��@�댏f�����;�8�m���H^:�=�����z�Ev�y��/������*��sk�s��=����(=���<X�װ೰sE��7��v�#g�u�j�mMnݪyO��⃎�vѣn�<��P�"�#�<`k��ax��8��+��n�9�J�O<n���a��DoOg��v:PN�ї���Cw9�vw!��Q��sW^{����gcz�;B��n7Rd=g.ٺ�2����t��71�s�'/I��	�>���<�n[c]\[�n�]�U����3�[=v��Nx�]۴��f79�p��j��M�ֈ�)���m�+puÈ�]�Y6���wE\n֞�n.C���ю����6:���X��m����A��n)��'v��l��{�[nc�9�v��\�;#�8-��mk�� v[��պ�OZ:MۮBlm�����y��.�nثqå��[��71����(�Jvzzp�`|h(���!��:��b-/ǳ�s�b ��dG�]����,�6����+��%8��Ogpgms��v��ٓ��{;���v:�m�kh�so\�nޱ��Et��}�����ư먢ތm���ņ��i������Ԃm���;;�l�3�=C���-F���2�^w�^��#E"^z�έ�q#��I���u��sz9��Mێ{um۸�=�A�ƃ��vn�GnL��\p]�<C[�:z�TJ�''�]V<Y���8@y���/�����&:\�x5Ų���s�mv�x���9E���=�<gE]���t�|�ixL[�� �<��v���p{k�E��.��ە,y�s:�m��-�G���8�ۢ�ڷTN�]�L�y�
�̺xuk`\m�N1�g�i:����÷֗���َC�m� �u� �=j6S;q�h;c��q��v����_P8p2�0'�4bx��'0���
nu�lc�	n���6+��psr�eGm�h����;v."n��vq���~o�Պ��z�����g����an1���nl�ڲؖۜs�F� ��߂=����i`H�wW<=�Ж�W[���n�nv�y����y[d�Inw&�v�����p���^�6x��l�޽n�-ɥӎ��wj�	�,;��k�<gptG)�MW�r�S�`�ݖ����D6��i�Sp+�W��;u�Z����v�bwr����,!vu���z����?��w�BC����@�2S��z�~�rqld.f�E��s�#FvN���v'���=��7bճu�&�;Y�т�g'c\r�ll���;-l&���W��۶�Z%�
tWo<[�4����Ә6ܽ�8���lLd�qC��9�޴�ή9 ��p�E(\n'I�x�# �{�+��T�����U�iֻQ��l���X�jܷ\W
o^��=lA�kd�G\�8�y/ pK���CeS;�ф#{=]=�֛'|E�WEۇ�㔬�`�z�Ղ���]xn2q���s8y�� ���xq�y�m�'c@瑳>�4 r�ض���Ęz��n|��;='b�=o\m���ś0�9f6�ܩq����˞��i�e�ŝ{{r�"V=�h��#��x�Y��=s�-ٓ�{��ݖ��q/1j���1t�������tzL����:��]s�(x೭�ǧ�v�m��u���f�n����=Oa��.wB��Z^���:��:�BA�g���w1ڻ;D�������mn�2��g8{
^q�91�vz�=������y]�V���s��1�ہ� ��m�����{]û%�i7o���mhϣ�'Y陜m�I�O�8��z���8���ֶU��SZx��.�%<\C����F�Ocp:8DF���3�ظ��dUm���M�`L�����ۛ����#��v�!ft�lmkO.�s�wW]�ގ6�v��m�;��b�m�r���&/i�nOi9����'�ѡ��v�gt+�c��J2`g�����s҇煝�ť.K�jb{ey�Ϸ�D�:OO��3�{<q��Xb�v6g�3Ⱥ�N�=lݹ7�S����<�kn�KxI�������Ͷ��ͫp$uĜ��ڀY�o5c:��S>ڎ��7"���<��\Ǯ@���tmCgR�{[�ܭ̷'Ѧ�{�*Aطg��pμr�*GqE�g;�ڝ��f��m�>v[cO�f�Zv���NR����s:�����;�땔�VXњ �@!HB�@�,��)$	n@ZzǢ�'%cr߁4�H*ʈk���e�e�n�j;;8�N�䓌)vN6��f���a7=�r��or�0=�쾰�;Fv6ɸp��x�p��Mn3�㑵���@1��E�ۋ:{q���F#�Y]���n�y���k��iϞvϫ��X��Έj:����v�L���y^�f;]��{t'C�Û�Q�]����N
t�-ڬ�V4�{��z��p`�'�g�)�)��g`�plv{n��nw��0���$�\V�/�5�����?\�%u���i�ʞayS��a&�y���dkz{U\����']�Ii[�oT��hq��Zg�j�U�4���v�*T���R�����ag���5�Y�* 2���cU��q}&��hq�F������>8�m�����ߴ<Il��i��
r���z�x��;����];YV�@�g���cY�nSf4�e^�f����O!hi[��W*������z��?���*����Ep��s2f����7�a4�-+���d���f�e5�7'ʵ��]�ɬ}���m�m�_+��T��n=�浓�R��V{�@PϮ�β[MUN����\�m�e}�m�?g{3��G��m-?�[������x�y�}�d��C�����#������J�Xb]�hĖ����8���z̆8�Цi���O{���{�9��M�TLN�m/*���o�l��/yd=�ֵ״T�����g�(���,�hQ�yeT�"�;R?�rO�{p=7��OIZv�3���s3�P<V���>���^������]`�׃��w��z�@�~�q���;��V�sty�i*���׽|z�j�!��n�����u���G7�3u����@�:a�g��f����d�;�{�U�㒲�p���8�L��Ah[����S7\�Wv��5QhU���]ȃ���+
��#x���ў�)ء��^|;{LJn;[�҂�(�Ш���uޣcn�����{�oϚ��W3�F�u
9R�o�5|��D�b0罼&�K�M�l�oj��SI�{��nc�-���ۧ}�[�ScKkJ}��ȝV� ��'n���h����b��s~�6���]�Z.����[��̿j��ߝn����'��O!Ɠ�$<�k/�5U2��/ޢc;�\<3���N]am�V-c��nuۈ:ַ�ٲ�#]{C�3k�(qHiԛ�>F���n�؀M�:�X�G�L`XŶ�d^ �����u�R��w�=StWv+]ޝ@��_h�Öi�s��TJ�TV^7��y<��U3�c5��*ku���Z��d�=d��r�3��
����q����Z`|̭}z4m>C�M�����/}��.��ܨl��WO��{�멌����e�F�����
���x\�Q�Tѷ�˺۩�[����㵹�˶��k.��|z���ҸWhy���P�S�6�m|��1��8k��u�Ħb|�32��A���q��)Ѽ,��^ (�"��bC;�u��T�M��%2s����U���UVy��i�%���v��Vc��ϝSt�ܶ��6h�;�}gM��i�{����Q�q�ғL�}{ӠY��E��Q3����x�4~`׶���0WڇՈ#�19�����،-�#��sl>~Ld�7gɧ�[6����f��i�T���>un�l��Y�v^��{��ڔU�{�+�_Z�����V�����dc�8��Yy�H�/xF�m�EN.��KӮ�y<��b�k&�k�<�ΜIԶr������I�4{�8�R{����3�]��>d���q�e��6�L0�'��t`Z0B���� �>�[�6ÒO���%$�{Y8��l�S+�������$�����BļX{(VZ���������2��i/u
q-��Ag{��!Pۊ�[MՈ},��������{��&ҙ>v�P�eǧoR��q��c�����`c�/|��m��9�Φ�f�P�\�1�q�NP�!���AmfK{(e�0�"eD�e�!�ŝ�>�Ӹ���%�4v�u�9՞��@kMϞ=h��^��I:���=���?�Q�ԇ{�tѴ��Lf&��E6�h���18��aڢ��_�Z�r���ұ^���$@�_Qy&G�[qxo_^]ߙ)8��H�G)ޞ5|��yYwy����u�q���{���S|�_mH�S:���������^=8��l��x�*c�P����e�����]�)�*��w)��a��?��F,�5��w�W&�e3����Ʋf#��uxï�y�|ɷ�(��w7����Sˠ�&��R�U��u��@�kg>;ݜ:�B�A�;��N2[|�2u�;��s�`�j���CL�8:�7�X�e9c��a��5V_��6�y��=��O+�=M������Rh���}��7D�}tE-=�y�^_gk�ЁDG#�x������R:Uz]��K�S����۹*£Zւ�.���<�۬���J��y��2��d=K�y�R���&V|� �N���z���U���i�}Si1�=׽�R����e�C|��g;�Vt�=��^$w�ө�Q�Mn�;�����ܔ�<�}��,��c��s��K��<��lۮ啪#��>ox�	ݍ4� �r���+�5R�^6ַ3q�1��WXv��p����0�����7YD�n'�A�/.�t����N���l�_f �=�^��w��dR�q<�}za��=O}{�w���l�B�C�6��5�@�x��r��;[/�Sx`��r��8��8�\���4��sY��~U��ԕV�skHz�����!�o;�&�S�|������l�_*�=�'�C?Z�V~o:���G�yރ�1}���X%�ƞ�T21�ps2���F��N$ˠS��7�̆���D�&+ew��]ϓ�Dǉ��o;>���I=��aI �\�ɺ��)15���-���z�*_������U��֍�[U�Wlt���<z������Z8C�}z�>B��^�f3�n���u�_���F���-��`����s]��%��j�U
/}�;�sT�톮��e�x��_T:���޻�!��·�7���-�����2[Oj�1u�j��C�ʠ9j����iZA���{:��f7�����buЬ��-sמ�y8�@�;�:���l��2bb6�P�Zh�I�*�$|S�.W%���
2���r��l���^��m��{O,*>`n�1r:�ϭ�Z8Y��䡑���u��3�FW-G �+�BZf����eD�[���0�������ɻ�5�uS��:{pqky���T�^��NSmM=AZ�v�z-jj�Ig����#�g��,<������5l�q��3{����'�^3���BX�x=j�rBu�Jp��v�P��l�s��q��}��~~5�wn�|H�x�UI�r�0�s�kl�7O�^��l[�7Y��]�N7��l�Qky��9�Ɨ��=�QC܉8�;j��s��ǩ:�h�e���m���8ߨhN's�<��w_;�i�Ǟ�=K��������}���WT�2�gw�6ji����������~C��O�[C������¹���O���o#�A���x�aI��'R��̋<���dg�U��l��������P��h|����u~O*q[C����>�s�}�	Jssӓ�Y{|���Tc��`�З0��I�_��Cl�w�\�t�x�û�ZK֯�/������E���0Y���d��[Y}�'H��V���ʛN:��P��w;`d�*�����58�Ԙ�E����$9��6F�/��G�}dC��*�_wZM��;��|u!�n�>d��_&��}�B��Z�J�Yo9�+�����:]�m+B�g�1���xя���qs����i�4��ɏɧ�-���9��e0�%'�߷Y�׷{t�s[����X�-�`>��jʇ����l�[�_�c�q7���m���f��
u"��Ơɣ��1u/��(6ێt<����u6�و{V�ܞ��]�c�����x�J=�m��%��~{��gD��c4��s$� �Y�}�5�PL|���^�n����GY�e�F����s]��z�Cw5a�s\��I�h�-֨��z޷i�.�\�+/	����R|�����fs�5)���j�f�[B����̘����vh�p^��؊Z��eF^�q�:X� �ŦB��q�c����d�q���
�u�w���f�%��f�w��@�)6�E�g}��N�o�m�M8�<�xM�g��5��/6ޞ&&34��!���U�t����ziu���Z�o�н��x�i�;D�q�W��`�0� B!��v�u��J5'�YTi���F���w]M=C�bbm��M���Ѭ�i�0���yZg^�X�߁)�Anq��x��2/]n�[���|G�#��
�H���	LY��Pwϰ��@�R�eΦ��uB����2�X,eh7�=�����Jg^0�(��5���I���Nぴ��6�r+ a%�~�0�|�k���v/����;�[)[�yG�&&��?W�|4��di 3&f�z��U�K�:e{��w���pۤ���x���(�~b�5��e��T�V,������WF��M���*�w�/dDnv�ueyNOh�s/����J�׽�߰��]=��N;���D1��c�9F�w5ܿ�l�B����w���A�l�>����8��y�~^�P�a�?hKcT�d���?uuKX[Y��q(�!x�������Ⱥ�s}~�9�(��1��y�n��5A��<�Ӵ�N��d4#���m��6��u��Mn���/�l�B7|L�m���P飄a�z�8$�6ahO���Ci��4���y �{��ۭv�f���Y1�&������g7͝�m�����|��{��Է�K�L��̀[�n�/&J�u������̪���E��L�ɰ�J���5��f\�4"y�>�g���?��U'Z��"��(���5KHo�^��ѽ֍θ�����}�8w7pj9D(���Da��?}1R�Z�t��N�U5Z�&�uG��A�n�d�k7�A�R[>@��^ϓ�m���v�#���wgk��י�tX�D3��4��Ԃ�{:�6�b
�ke̸m�)�e@�ֽ�R�8����z�kz�Mոf�g�Ϫ��40]:q����8��&+������;r�vi�(>@�ɫݚLf��[o��=_�kՃl��	Z�3�VG��;2�����b���F^���=��+��>�<�dӳ�,��8���8�qү�r|�v��o�}�[f�a�O��2�C_V�8�oz�g-��f��¶�%��O2����W�4_�&����Ni�t�4�R�uE%j���u�����$.[�@���g�'�<~Gȍ��>T�/��g�-�~������)�Ҫ&<vΰ�V�0�s�.�6Õ[ކ��׻�����6��s�=na�2U�6�^V��))�&وv��Y�&j�4�g�feN!mv��~����]΋�;M+���7�⚾�����"=J4��{ׂ�F��t��/J>��s.��j�4�nټ�u���׽cT�wrc<���M0�-�;[ֵ����O;�ˁ�љW�ǉĪ�DS��0�/�C�|�ٓ3
�~�/LZCʔ�S�Z׳��h��0컟K5Vln���O�#�������������o2+�y�P�i樁۸w6�����t�t(;7꣗E��Ek*�����i�*[ItPR}���H��>`k�X��yc���������u����n��+��ZN3��y�L������G���h��<�ua�;�.0H��RW�{/F^x���� &-[p{nm��;Fx%���gn�;�����I��'�-tB��X�S�Z/��͉6�ϵV2bu���5'��'�0�JN�����L��iY&�G�r��q%U��ѩ�}���u|(�ff:#�?Y��m���+��"����*��ms3-j�/.��en��M�G�i����&����Ρf�7M
#�	s�Y���ףP���S+5e�-ƞ%%wW���:�v�n�H��7�R�d���g��V�\$?����MH�%8�V[g�x�;�%��L5��f��L�[I
a����f�A�A���S��Y}�Vl�!�߽�������Ͱ��z��q��7�ɚ��lN{vM2�[�.�f67�XT)�_}dS���M^bv6M���_��D�l�m�+��~����T=�1&�����i#�?B>Ƚ�>��ϩ����򘾅��p���N͏v�%����hov�=ˁ��f!��^�̯Te^�fVfb
m�Pi}U>a�R?[�����O<���N0�X���˷��e�W�ܚ�o�)}�1ǉ��=����w�ij�ڒ�ZT4�5{e���������(�~&]��^C�M�p�:%��e�ñLǛ>�1�����L�D��r�����s��s���Ђ��xV����H:'�jt����ߺ����9��a�hE���;^v�ۣ���w/=�����vxx�nh��<{k�<q��Qv�3s�t�S���h�vkh�����ܰz�e+��8�q�l�G4��4�G��3n�9����+q#>����c�Gc����ם�湓��z��xW�s�f��u�"�!&�r&@F�[t,Oj�9�*���mX�]b�kf<s����sۆE�Z�s�"�1�Y�I��4�b����^s���ms��1���>�>,�D~k����� �a�_}�����
�,��l�q�x�U�J߷��{�7�j�畚a�-�U�&ҹ��ѵa�>�8����T8j�2�n�A��9���dx�.+�@���l�1�[�Mp�k��߷|Ka��O�h��j��'l�O%]x÷ZN{�Ӡ���S-3�}\a�v��G{Q���<=��S�e����>�����h�-(��Hz��i��;V��n��yW>g�"��\@?k��CZ��}�4���W9{ؕ�)�6��S�z�*r�zʛx���-�����h�1�2���C��ٶ�"�}���u���Ae��m%�8���W:R�u��~Wt(������|H�:�^��<�Il�;��
L��p��f8��RMo���^���r�{z�$�[a�9�����x�t�g�I�����V��t���՞��m4�������@�E��䔪��+뿾�Jgk/�6v�������8��7�Ѧ��L�R���w�9�rV�6e&�z#�`�{n��e2�R��f��l6ӻu�
u;��g��]�[V�~��������,8�ƽ�j�����q�l-%�ɞ��My�b���1�1�L�k���N����}w�}Q2$��Z��u���m8�:b��Yhm�}MaU�����Ưm��KC���R�#��[/Ӌ?8��gg�����w�[zb��%^ܴ�9�a�,�W}�xi'NWg)>hǣ6�)}�,�)
de��o�~�����u��~�u�p�{\�0۵kw5��~�΢��[>Kq�:C�����{����O��eT(q��AAm�;y���_/uz���p�8˥�Gae��X��ˎKf���R�N��y�m8�f�P�Zq�{���Ւ��t����y|��e�󧞠�o��!��+*�[f�����Ę�S5��Jam����Q�|�n8���	 �C�}DCG�=�C�wu��i�q��� Dh"ȇُR���{S�o�5r��[��1��1�f��8��|�ʦ}z�Oȣ���4��{�h�a껇wX�1�96�0���FHg�?a���R��OkٳA�CəP��|y���#/��q#Q��tV��Da���󻣿T��5�{�ͅz����VJA��?{��"��`���,�G�T�s���.���׮[�D��i�H!�D���u�������"�=m��`��S���l�V���t��߭��}ָ���*��*�4�u�ֵw>N&�\M�B�T)6���z�k~K����9�6�>fj��aҫ*UK�G�+�F�S}d��{�4&����ڬx�g��a�d�n]V�]��e��y����^�<���V��׽�}^=���l�i�k��8��CL��>iި>�}�A�aO׫
a�:�۫��hm�s^��^���l�iķ�ٞ��-o#w��m�c�m�a��ZRU��ﹽ,��a��;q4���3{�6q4�(1���=�!��v�ilW�WG+���L#lM��9p�H��:ɚ^���+�j����X��;�0b=A^W&�ʶ6�Yۃ*2�'����,�p{`vf}��H�;�Q�=Y���p{���VI�[z�	�����_m�|�ao	�����w�x�����n8�X33�:�*��%s=�x��%*�X4o�7nt��Nd�4�n*��z��U�1�tZ峂 b�gk���,��u����a�(<
;J�K{�M�:�t����1�<C�����,\�=�:���{^PKS�F��'�*9�U�!�րt��	M�ۄ�ԭs��w�{G�	-�oK�{�6f݅�m�2��.dB�W�R�.�o��ݐMĠ�ܝ��v�wOi�x��m���.�q�md��T�����4s��H���+�'wE���o'nX��#��w�>Z�H(�L�(����3���N6�1J=�V�c��P��b�`��uR�m7N�a��{su�X-/8�`�-�o/Q�1eq}4xx���\���7����7�;Y6U�5�!\��/pa��m�z�=s��a��x҄na�v�⽾,m��A���_ֹ���_I��:h3W�e�8�usu!��<m��vu����֮�.'�bt�_@�a�FNkn<��[9�J:���Yk�������`�v�^`�W4��i/�%�ӸǊ���q]"��/"����\�T++U�l�S����LJ��c6��,�����X�.��pC2�Y]x^V����7�U�����Go��G�#᪢
AH)'�2���I�0�����f�)
II�����RAH)0B�TC�PJH)!��0����}E$2��S�H)!�;�{ ���R� ���P��QUR6�IUR
b$���� ����4V}?c��xe����.�)II!ʨq�$V��
B��]Q ��UH�k���qܤ����
C�D����-��ˆ3;[����
AH)�B�S4�I �5Ty�
AH-n�7D���I!�D4�Xc
H;�}Y�
ACL��H}��=�=� ��
H)UR�) �5TAH) �2�7tKH) �/5�׽�R
AK�,HUQ ������Q
��) �2���R
��_U����eW�U[`S&�I!���Rq
H)!ʢ
AH)�D�Q ����Q�0���
CUAI) ����}gj�^]R�ce��y��wE�>�Y1 �*���Xj�
C�DJa��RU"� ��RAHePm%$��wP�S#[��z �:��
C�D��R
C*�) ��Jx����D��Rq]Xo����w�sl�e$�y�齁�) ����Q ���ʢ�IL?0���wD��P-)&!���Q- ����7�.�) ����j�) ��U�9�,��R
CuDʅ�%$;T��
AH)�_~���$8��h���;u%���$�� ���RTAal)9��
CuA���ƒ
Ae�e_����u�����,�+�K!5;nz�GV�-dZ���'�a� 8��������YlŻ�*�2�� ����TAH,i �2���R
AHeT����SH�RTAH)��)!�}���AH) �q�� �̔�R
CUD��Rl� ���R
C*�,V]$?����k�
AB�RC*��[s�P�
H,4�R� �bS�P����Q ��$*�;�%�?4�R
C��x��) ���}y{Hj���R
O!Hy'��)��RAHUQ �׻�Hr���R
AH9�}Y�))%!I1�1�� �l
H)�@���R
CUD����i!�����Y)��R��W�e�ta��c�R
AH)�R�H)� ���RU&�R�
v�@�����[M$���肒����R� ���{��o���-��p1 �*���R
At}P;�AH) �5TA`<�d�RAHw|�M삐P�JJ@�K�N�R
AH(~����� ����
C�R|�a��R
N!ˠ���4�R
A߻��D��Sw@ZC�D���
C*�@�e�R
Aq��Rk�- �;˲
CUD*�) �=���{ �<��
C�D��R
Z�s�5� ���R� ���RTII ���_V�+�5yeZՕy��
AH)�
d�r肐Xui!uD��R
BꤶRAH)!���) ������w�Ri
H)!ڢ?2RAH)UR
Af2S�귀g+��aI��� �/3����R^���R
AH,�cTAH) �.���Xg��u���n��U�|�R� ���Rq�}D���AH)�{�{ ����IUR
A0���QW� ����ۢ
AHr�
��bC�D�$�����;�RN���
AH]Q�d���P�F���X~a����)4�I!UD��R:ɜ�X�����ʼr��Z�{�
AH)���Q �+�ZAHj���1) ���I�}����߳5��U��0���RTA|�����P��k��+@ZRAH)!ʢ4�I �5TAH,:с���RAH)��RAH)!�����AH(q%$�j�) ����Q�c)!�КO�āHI��ޚ��Y����P��7��%��M�i a������f��o�3u�2_J�$����pbv^]��M��R'25�fROk��J罣�u*����o(wf<��}Z/��_|^wٟ� ,�_u���U�@)��Q4�@�I��Ē�6�V^P�Y�f^f���a�	���H@d�jI�$RC�	�T�u����u�K`C��a;���>���Y�?�L���)r�@4D09���2-�k|4��6�y��;4�Sگ!y�W�����e�=$m�h��n;k��$	F�[Qi%[�}ո��.i͗��[�9���:�CU�(���9X�ԙ�+�j/��go QmR�8$*�{�@�qFҒCW�mK��O4�csy�����
��)Kr�7r�HV�(����ʥq�R�;��3:Y��_z�����R�FFD��j7U�Y1*yŃ�]�1��K��Pv��5ю�i�&;ڱ��"B�0g[����y=�&��hYk,R��M��a4�[#�� eE�[�'�
6�zGY�`7��E��M�Y5>�\D8𣫳�x>3�'U��P��nI��ç�yy�u���=x���㋬h,Սm���$q��_����8�����m:�'�{MP�nB�P����1O�B�Y�X�
�A0s8F��b�Ws�)�7��������s2�n�\���	�^�9��CF�n���x> ^V��i�v��o�N�u%�V��\7\�\t�ۈ9�n��ܚ�1<��/m�;^��dW�l���.�����>w=Eա�T�t4����۞��ˌ)��j{'�ɼ�W;�;`��#�u�۝ƌk�ڸ����1vt2�tx��6��x�;;��d=pS�.��l�&dJ7 �v�f���Wf���[���h�$u�t��ڻGX0� 	��z��ZmH�Q�kqj�bU��u���V+*�Ie��Z��=C���wf�*/S*g�}���C}$��%׮�s��u��
��Q��]����+�X�$RpK����&/�KZ�㣠z�C ��玱@u�vIm,F���^OQ<�T�gz�^8p��2(��{.2=R��X#$��0Ғ&q;��C�o���	��t��S�i黮�>�я(�Z��nm��3fEJ6Q���(���Kl��$e�'&BK�w�<lֱ��m�'�ݝ�Y��lb��^E~�W�#����#�4���Z&���ǂJ!��ܱ�7.�-�+WȚl%E�	es^�$Μ'OT���W��sY�����楶�px��Ö�V��~�Q�k	�(*��EvV��>��6dnH�s�(WJWTMC��l�۵��p:ֈ���9I����/~n�_n���2�n'27ch���]�rG���[��̑�m�tK�OyOn���)-����9��f��O��N`���;,�{��L�6]�fֱ�;lL��p�sv�쾹iF��ӵ���_P�Ń�٬	�F)b+�0�aN��U�*�X�7EN -��#Gun�Z�r�ߵ��ˎ���Pg��Em�鄭b*��!�x<�h$�9Y4�׷&[����f��'�������mu�o��u+�UK���Y�.���������M�nv��>������s8�A��1IF&�:����!g%����pE[S=�S�������������<v~�Vi�ǻ=��@�[jL��_g�r���
%��yab��d�L�<��)��kS�۵V��L��іED-.��$�^�}�n�f,�.}����ɡS����'n��ѹ{k7�]� J��4�:2]\#�������n���zk�����L�y�4I�+ϻ>vWS�V{{p�o�iݒ�q�v�鏹�dk!e�vzfK��q؊�����)���E����p�-��z��&g�t����r����Ou�6�1���k��۝r���)MnS��PD��)�a�,FDEnЖ���t�R'�rMk�[���Qwg�`\s&bW����쮹�����̻�	Gt�Е�)E�X��dM{}��6�])>u����ku���V+펆��e ���i��}���K����Q��ݥ�q��a/���n�.��&J�/	�##��"�j���֐���9僽m��^�p����{h�{ݞ�պ�Nei�:�߳d��zz|�Ь�d�`i��(�zuQ5�$;7����^P�<�.ϡB��:2;��Aq۰p]p�ul��y;�����������w��
�b܀�~7�[�������q������v8٢y�6e����vl��lV�"��*�Ո"�7��=���5��f�׍;!����{=y����l���]�6������ߕqOR�2x�U_��`J�x��E�d ��R�g��y��A��֣��-��7wh��zY�k+(OyRW�}I��+d���v�*����(�����<&��Ѿɣ39����꫻9�����7��,�u��=&��un��5�n�*[b��1V	5r�I%ħ*O��8�j�)^��z�x���J���el6��]&�V��h}�A�}~^��bo�M4�;e7�l�Gq��uv�Vd��^G<Ĩ	�X]\3�KÜ0�"�hq�<ʚlS����ޛ��t8T\�r�cECӢ��c��e�#n����E`jV���q#�_Wu���2��6�Y��Y��I:��5A��α�>�&Ҽ�ʇY^Qj�Tq���I�����U���n���R��q��-�l��c��OtݚK�v.DT��Y�T׾3+�T��&�zx֟8�O�����W��Ղ���'y��B�K1T�}2dV�&LM3��[&J[u�ߑ�r���46t�½C*M;9�����^އ���{[�(�ߴ������FrZbC�DLq�-���b��^�o��z,9[}u���Q�ZŞ8�t�k��N���j{���x���� I@��"/�I�n�����p��=�%n�Б^m7N׽�L�v�89�[�����L�{du�P���J's�u��q4Bd���f$^U۹�3E1j��<pN��%1^�8X�]n�ż�S�:�(Z6p<[{���a)�9��%��J�f�+"9�Jl:���_}�rd61Y�unԎ�TJK��4R+x� �W,��UçX�&I�s��[�a�.�\���ܾ�ĸg;��ߥw:w:��1��3�l=�:�^j��q!<�f�ͽ�ݦ=e�^���L���q�ӱ������z�����p�m�N��iN�`�zc8�����\vV�s�����B�[�[k��ݔ�b�ƃ��9y�@�ɶp�]~��m򕞒��k[��-S�맞Үv���஺5Fցi^Kk����Eᶍ�ln6������wn5gy��-��b�"s^xa瓝�
k��%�Ev�Ϲ&n�z�Ę!E8x�������]/{��^��K�4!fY����t������כ/\)�[oQ>���@P�B*Hk�0ɉ�u�[�h���#ٖ�@��[w�zu�����#����[�콣x������3�@����fyQ�!�&�p�N~�B��죝����;��
�=+&��rZ�w=��݁ձHݷ:�˰m�-ֵUY���A�k(��xr�~��^QBj�rLN���ݶ�TS�}Y�ƻ)�2�3�^r�պ�FP�|���3��`��O��g�󜱋0vKIE6�A0˒��!����/��.�#�a�m��9��MMɖ�B�����i�q�{��B�/[bد}/�3[�n!2�'��r��۫���fg{>Ʒ& �g��ϱv�1;`s��z�Ս����M��_���;��
}����y�ݬz��9�=�3O�.��8-K� ����ņ�R�֊O�d��!�Lq�t�\��<�������Q��UJ"��r�цT	�E�r��.gf�`IG{���R�"��[�殬щ�]�9���f�2/.I����>�E��g����?��.�.���Ie+\��ȼw�pS�I�/os3zS�X'���ZA��i�$μ2ĥD����[�<^;}��{��h�{����¤��ǗG��gF*���`�;w3僔����P�T�(�z��M�wo��n���v߼�MEP��$ʲ��-;�0�)�יQ�#�}J����f�u�n�JP)����H���b�_U_���3�T�{.Kα�`�2ZRh�d���;Bǟ��[�%g�c�]/<6:�L�re	��b�
Ik��<�m�b�h�@y����������h�Yv!0Z�Qc�*;J�9����g����ҋ�^0�C�d%{ن�/P��d>�&��=�P�u�W]�8�LX�A.3p�p�0��%��[ΰE5;t�Z���W�Oy�jk{�A��p����c����[F:���pgkY?F�1��R,�U�����}�1��W����j�.�ѓ��n1� @�6��	�?1?� z4{E9�A�ct�4M�>��M
��[���*9����ɓ0o�I�=:�����ߏL$�{EQ�vF�Q��q3x1|Kn��ZⓉK����.߃O��Ǳ~�����x�|ۇ~�O]�{��T���VxS	�b���1��q)f(xT�`�V�3��yy�v����0r5QT�'�ټꁬ�o�MV���:����ZܻYfR���-߶��C����}b��g�k�guԹz�d8ݱn�z�wM��dcrF��F��Q%{�ǭ�ܖr��ŏw���W��U��!K�\s�s�dh��g�}�]�m�s��Ԫ��\p���>)Hd�~r�M��A�ʍ��zǠw������!�Ԫ�x_	2m��f��؞s��ԿeP��J�kd8� No��Y-��-RK� ʭ��3�¯}u���Ȼ�_"���k�ں����|�Ł��^Uۊw��nm�R�k��dޒ��P��L�\!��O�.��n�2�^Z�S��[������5�z7�>�I읪V/8&�I^��s�P������-x*�u�L;�[��X;O*��t��*�kWR����%j�DNYֲ�uN%�1fL�Ӱn�C>7oVl��=�����^=|A��<$)a��둾���>=w�uX�gJ�%�H�����I�[�S��2��
��-�®���c��X�=�頫�6
�v�P�Ќ(R�����Ts�W��خ�Fe�Υ��������t�,�uAR�QE	-4��'۝�������Z;�[ݽ�^��3|5C�CG� �+VG�Rh���b�&C�A(c	��Ez⃫E�{���.�)�>�}��\���H�n���`'�x%W~�m��G<ω��RM5+��}}[�)B~�5�W۪~0�'���+ol�&J�{��{���=�0:{�J9��m��c�<�Har9���I��|��h$�U�Cw�K��"]�k7���D�����ix�t�YG�����y����T˷Gi<�y�z�TۻQ���n ������PS-��N��E���eA���Bm���'�,O�\֟&���Qmm*Ͼq��z#X�)���W���n]T��Wkl�h��2�i�-��F��u�����`���e=��)�w&]_E6,uZ��g<m޲�n��qp�$�U�ı�J6�C��>��[]'L�pH�����o��9:���Z.+v���c{E��!&�GS��9�
��;�Szyh�Ѻr��R<o,Ʌ�n.�,Vk���t�Y�C�9�_�ppA�/2��k���r�Ѹ�]c�wuV�.�E�<|fy�ɬ&57���>u@��64i��z��� ]Po�]z����Ŋí�{Y�{��bh*��jb�M�jӣ�r�ݵ����]_��(��33-�B�&ҵOg���}G�rxn��Ep�xt�x�&A��p���_ ��+�Զ�♰�j�;x�t�gL�;�{�_T[�˭��Z��a�x�.��>l�Q�y����ECM���Mv�:���Wg}1�ޫ�
|-u3���Y��qD=�4�:�험�/�2��Ah�}q�U�l���7%��C�\vMb�OK�W�j���X�TŜ���rޭϰeuN�PtF�6�B���PЕ�M�o*p:��%T�+t��P法�VԦo�'�v��K�8 +�+N=�Kub��S���K)!uǮ�Qj��H�ꏘf��Oq?w0#J�jFf�	�YGh�R۳�8�=��c�r�5�����)
e��O{}p��ɖ��>��+�<�(�8�'v�ᾴpu�9���p�ї��� ٮ�;����{���\��0�+�l�5�t�͵}1����aud��p���x( l��X��ojS�9��ڽ�6�\��ף���̗#�i+R�������K#����tq�c'Gsu�n�a۴�C��>{l��V�u�El��=Q'��@�6���C�1QH}���g�y�Sێ�l)Ů��]��<��ӻF�	�$X
ۋ��d3�ǫ��,�]ԏf�;<�\�/GC�q�]g�Nݗ�z����v�erѶ��qf�c��ݭ��{$�y6�׃���)om۫�&���2s�!�nzLݦ��ܼN�S���]�=v��9�v�;r�k�������9�c�y��x�m��ຏC���-éW��v.:/1���y���O3�ۖW�d�W�x:�^z�Ǎ�zC���V���V8�W�s'0N�;�Pv�Y��s"����h$��]���q��O���K�:�g��5xl�ZE�7kUփ��S��vw��n�mv�v�պ.�n]'<�WX�mv0�Wj^+q�ou�,�1�����͞��Ǡ�tQN����/��f�c��䗃ta\ ��ֵhB����u�s(oms���s����g�q���Ⱳ�����a�f3F^k��@R3�ؗة�eqq�;� �mpeϷj��Qŭ�4��gv�>Ru�����B��%=���2�UNV��R&,ۈ��X�ۘ��7U;����Oj;E�C8�]��uΎձ;zt�8�e��q��$:ln��{l�JƬ�b�����1�I{sw*�k�� �y��-�.����cAh���pqhݹ���&��t����n�r�@��6�n���������.������/=�rf��9؉��.�u�7�	!0�t���tf#��������7"��G]�n�;#� �ӑ}<��7`�u3�t�
֎0�{n�A��k	�^|��{ ��w6��cG=N+�Yڽ�a�ѳ���ݖǄ���- cE{h��ú��}�Z�[UK2�l�.��h(��������B����q#Om9�� �:����Y��<`�\�j�1l�O6lK������g��+�x1�fź�������;�6��>�vۭÃ�����ô��ӥu���kn�M���FB�2�X��#;�v�˺8w]�7�T�c�G<��m�\�z�1����n"��׻X�l{n�h끍�r�v�J�1km��j�Mh�`�eݥ��p޷n�Ã��*�㵎�����X��z�Rq�'��9�;޹�oZ�ge�ͤ��6�V��,�Ks`I�S���#)	�~�xR����,Q5�u���fk�η��{�ދ=Lu����X���*.P�)��kk/��f��H#�H��W=wx����73{�'����g'�:�l�+/׍�5�93����ݣӪ�¶��|E�ے��t#msqO�܃|����㴽�C�|諻�]�GY�;�(f]_��x�}2⭜�TDŇ}0�N�z��ԯ˕�~�֥�+c-6^}�Gw�;������Yw��a�y�,�^m��G=�p�ĥ�z*��kڵ�@�Z�w��YTĝ�-1(��aBd��p��̪�쵹��^��d9�X.����"���ML��|��d&W���z�;�6��W��D�c�<���֮ ���\������lϠ\l���e�Q�� x��\�㮝�]YtC�ܺ��&��X"�U]et���z�����{�l^4슩��{�`Y3���*�d�=.�5w�����P=4�.�6���@޷�Bl�(@A@�ۂ�_ޕ�[�����|�;��0����^d�乵j])�K���#�Jz����4����թ�okb������t�yz���IrZ_�,��G-��_N�_�[��K��M�F�)B՗4��5<�Rr!-|��ʮ5�B��k�ߍA��?ͨ|~[ rXv/�����43�F	8v�ْ]��n�7�:\��uޘ�F|�B��������gxJ�7ܵ�4c�5�W8����T7k=�#��ׂ�>dz�<0c�3�����oC�n��n��Т�*�����w�tV-�x�3�u�u���x,V}��`�~��ӧ��N�J�o��<�O/�t��R]t�bC6��ӵ仾�J�9��б���FA���[A��>8�[E�nn!����X�`�D>y�bÞ,��n&S�fOUU!��W��,3��kX���=Ԟ.�=�6���b���ӝ�뱅wەu���Ɇ|�ʜ���W���r2�9ŖPw���.�x7<'�����:��T4�G�Dsh���9��&6�[���߷��mH��=�s�k��X ��BE"�n��-��?_8Vc�;�0ػ]�{J�ݙ��*�n9Мy�R��Y���:ٳ��R�;��M�`Z4�)����\�\:tJ�����c��s|��e�­Hk��ڜ��G���޹�\v�A��I�d5-���%a2I5�Ϩ[檰U�X4+̛�iW�����[B7^Jx�0k(e�}���k�*r��7b�U�I��L���$aJ4�p�Xo�_��@��xL��HJ��F�7�znv]/7��Z����*:��e�#�v �!E�i����[�.�~�l%"WіHp�A��]S
�/h���TT�p�����9�@;�]�\Z�������n�\�%��^uA��]�ȱ��<�ua����	�!�LΌ�J�����Wgja
��i7|ҭ/�ډ�ap)�S�	r-�b�*K��s��.��&��e*�#�9�q�t�逯�{5��uzD�����4YXm�\0v�E�~7"kM_Y>: h��Q��(��q;���[�+���#�q�~�O�ն����ɗ�����9}!"������֫�z�5wtw���oAJ&�Q�^���&ܞL���}�*g�a�g9�dN�g�sF=�B�)X/9�Z3�變��yjoN��E�.L�[=Z:,&���t8:�6l��sv�E��Q��[��a��p)'��D�D���n$m��畽���4����h��ěd@Í8��x#�7s�٣B�<�
��G�|�g��r��F���Ttmg+�~�ѝOƍ�U��K.�.w�3m�N_.V#n�5CZ!�Bp����{1շ�/nq���0/��H��W�O�~�O��?&��ߩI-�'�;�y�<���t��7�͒d��oz��
�ƽ���]v�O#���{�Q/A��*E"~A�T#��������sd��ey#DB�.�C�?41��k�M�H�V��s����>B��YI}�}<�����i����19���S�i�>x0�="K���fU�{�W�=zu>��l#�*	��GZ�sA���r�I��p�`O^yʇ��:)$����s�������/s����9ý�R;5���ɺ>e6&�n��^���,K2�]��y�~��;$�=gl*@��N廰��_�V3�
灿�i������R�mw�l�ײ{9P���3�o#����V�^Y�V?Kp�&�,�=��XLwa�!u��i������HMA�2�V�-���=���`��
M:��3S
1��N&iԟp�	�����ѱz���J��'6p��GI,���h�y�r�7T�I�en.ɣ�Б�{q�-���j�v�[�v�41Ѹ�M�*�<G;�Ջw�0[�bH{�9����	�w+�b9�탒7[[�S��EZ;����m�[5�_D�s!/=x��
��Ͳ�H[�S���?/��O��ͨ��ɬn®wFp=8J�F۝.͒.7c�3�*!+�N�mFHJq�vq��snuw7lIm�����4Kۇ�4�aI�B�>�!̜�W�gj���!�Z�����}�7~?~���C��,*�ݓX���MWIΒ�'�&��5��j�CiY��������皫�Z$���@�!2H.�f�����^WS�=��+s{4^/+�G<���1�g�^v\�G!YS�Ӿ�����O3�s��pR��5���z/A��ap���MD�)��^�1�4�®�s��6�
瞵QC�[[<�ޥ��2��r�w�' 1Eq�V��)>�9�hg�C���D�e�`�e�^����V+F��~a�� 3>�~��>xu�ɕ��㋬�a9�ڍk7;�y���\��a´��ͮp߾6IJB�*v�i�w}�����/*�5�$q�bӚ�����D��;˃�.l"O�g*�S7�PlD��oU�WV�#w}1mVP�૆��=N�6gyZ�ژ	�I��2��v^my$l���쪧-���f�+��u�8�B� ���~�6��j�m�M{�����}��"�8��&�3�CD���O ����=�Ӹ�ȵ쏳>K�Z�I ��U��7H�+�M��fɠT�]��7��r�wZ���
^����A[[3ڃ�=�6�=�1ug`�A�H���lu>'�v�F��깐RF�w~w�ڶnȇ��	���dQ��}���,����\��=�:�'1���{^����Q�"�&�-��kֺ>�"Jf��9��t/٘�3�����h��-��oV{��<�������nL�@y�Q׋��ک��}���j��T1[�:n�q,�����A0!�]�K��8H7^W��a�n�P�-��R�cM�[���;w���\v�3������w��m_>�+�'�����(2&ɐ�ؐ�$��ɹ�h9��d�YĆ��՚;�z�{(>�rL��Z�k��+�Q~�ūMd�i�ݧ=�[R��Y76�E����a�*V�?z���:�����b��n�:ݹ�������amǷ G�۵��hG~}���|�kHU���tyC$u�Ҩ���Qč95J��9w��%�J�>�:�*sPxug�E��Gֺf��m���p�᪋���z%8	&8c
I<p��i�F����a9�>x�k%x�zc��5�قͯ�A��0�V3�!2�0xȡ
�<�op��v肜�S�D�j"!�ڍH�fk�=zj���׹p�gy�P%���n�;�c�Z-��s��ٕ�'��MwF�Ty�RY2��<{M�tF����Y�C}��^n�t�b�v�f�.���X�s7[�
Aۗ}JL"�p��64��uӼ��ob�ļN�/=|Xܵ��b��^=����Ïq-�Nl�"z�������8��V@DU�ӹ,��Ѷ~���xVP�-˺�o���FTfI1M;�� ?&ZF8��
vU�_n�E��]�V���(�RwU�n���F��ѢC!��<;=
?>츖a&�nQ�(Ug��n��u�F���E�
Q����[��j{aV��8��E�󋂃��nl�x�&��B��4K�'��m�@Is�ۮ�2Y1��n�[��'�z꥟e�t'{�1aʬ�Fa�?\��ۗ�8�f3���]VsX$�,�E9&ל���aq�S��(b�ܛ��{�;��~�/�,b8����zp��z�;�����Ǧ�!C�Eu�z/v�!FV�{�[�ţTZ��8�*��(TF�����e*R�y2����-��t�HS��I~���|��%�3M�+	P����gw�*ʼ.R���������
�SJ'ƭ������ReЇ�ʹ,�x�w�zl��n��H�M�5�_:��3�z��HաFZ������8���{C2Z�[�����tl.�	��WFwQ�/q����mH�*I"���w�E�l��̡2�Ӊ�cV��Vc��{+��r�O����N�[���On��;�w�t?Q�m��(Eg���'�ݜ�yTDH�v���.�&~��{]���ae���&�C"��yf�s�<��wj+���w1s��M�f��\��Aj9�eux�=4�����30[�p�G��Chj���7h��'t�������iU�LhZ�.������rq�^˶e��K´e.h���%s�	�u�5��m�����%5�k�����oۥ�X�-����J>����I���{�痈B �ߞ��q튢;�awy����_h}��y_�Dy&@��?-��S�� ��C������=�[���[Ú'�����3����aoT�,v��+��ȗ��T��u���}�����	�]}<XE(JgƎ]l����j���|l�<�Ø!�Aj1z��W��	�7�}z�����]~�>�K@:��� �mw^�/�/hd��ڨ��e0�L8�$�cIǘHZR��/���f���c�Y�BN��X��u�Z�5�U�}*]*k�ʠlC~��"�u��(�qut�ڣ���gн�[��O�����:��3�k�ɛ�F�C�u�X;�}3���3Un\�V�;ǥ>��K�6�o+*��g�h�f��ۧ9d��M�|���^�G ��N��n�n�I<M��u��y��n�#�}�h�λ���b�;e����<�Ѥ���4�g�uc�f�s���۷���<[��nB�n���g}�]K�ۜ�3�rS��+�ٵmۮ��qt�����ǻ�(Y����/j��z�Hu�m��u��N��f㖀����e�;u���y�*գm�;�8uö9릔�:�q���t�A���n[�i;j+p�m�e_Y;9�齫�S`��T�<{���=�pH�N9���\A�]���n�!���3D�u������6D�7/l�|50��;�V�bT�o��^�"�2S}|��.���K����2�ҍ$L�\�4,����1_|������[лU���,ؗ�������g��N�٘3�̛�g���g[��e����3EWBF}>-�	R+�FO1F����`=טh]�Q�E�6s��M�yE�@ �lKޮW]u�{���'���>
{҃_1>�wR�t��,�F�`�j���e�R���3V�C�ҕ�o&��eE�����CȚ!���m�x���D���B]	�L�g��׸��VC A�D�Q��(x�j�q0�E�la�^��z�q?��[�I���X���6��������{��҆�Ԡ}c�]|sŌe��#O�!�W�d������Һ�9��]��D5�!�A��tɼ��:k��������+&4gۍ���t'�mkP����-��w�F����?{3���N!��0�g�0�T-N���q�l4���v�>V��p�Xd�0m�O0+/��-��v��q��w��~�-,V"�~�SKm�?�܂�����|k�,S<�ە��NO㰎���`�C�p�ý��Y�c����f�\:�^I't���)VMZ
�o���o\��Nz���o��}>�uwRʹ�U�5�����
7�9F����͌�mg��y�s��u]I��yr1��R�8��((Fj�V�0�W�ra����4���Ʃ�ۻ�{��}��i�V�lT�J�-ο���ꭼG��ҁ� ��d��E���D^���Σ�ɽ�B{γ��-5���W�7�9Hn�Y��D:%�=]~5����p��j�E�Ǉf������߳�q>�&��������Jl.�V�=��ץ�>����.��Y
�ry�Y�������^(�|<�՜}hD4����1�`��(�k֪��LJ�w-?���х�- =g��j�����6���<*���3���셽�@�iҪ(K)~e(�-���q��2S��^���*F�drȡN�4iZ��G��=o�ҳ�gYɑ[�NEN3ie�ٲ��S���V%'�Ui��D�F�Hr��l�a������X2�/:����j��r#��~��S�=���_f�י�'$���0�-�"��X���v=�4�(��_�t�N���'K1i�x������.L��y:2�1o�	�Þ���+��C�e粷�_�yr:�7���6;lݮє���vn�/jX2��}���0�+[ʰ���`M_��w�o1�vxe��a�X�'Gρ��p37V���`����7�亲��T]
�b�9}Y����ӝ���]�/��Ь����v�&�x9�6���.�>�G�K0W<[r_[}m͌V����͌��z�H�ţF�v���|czu�9;�p�Vwo �ϻ��1�s;9G��=L���^t�t��׽�t^Ih���b�uܯ2Jӻ��f�\�i8����t�I�����cpₜ��o��vk��u���:b�ɃE�V�1}@i�(����/���
��t�F��4�P�}�q;[F�s5�я7}�.ΛSї�y�u�&����L�J�'����h�cwle�Vis$��*&"�ڒ��g�mTє�v����࡫� ����O���L&�{Օ4�f�)�ge̙���lH8�kg�S�5	%5d,���D�.�Ǩk�-���E�����J�N)7�`g��n�SG:�y.[꼐ts~]�v}h��mE:��^7�	���&G���r�ND�j�?m���ݩ��W���������R�^�]nڹ9�pi}�"Ҟ����n�^e�m�bL�$X�LE��ӪW(��]XF㾋qo�z	�����v�Ku�͝s�+e	�u#��v!��
��( ��u�8��r�fԽa&w�����P�H>�y%F�.��/���0�R�v��yC��������K/�"�	]����(�d@�2H�,���*�e�Ȟ̞�6��bl]�S��%�w�¨�$�oדv�0�>�o?XV��p���dy�0��l,��E�>���㇈��V�c��N���9��U7e|K�6 H�� 2(�va�$�A�a����s��fx��b���\��7�i���(�9S�:��l9�n Y�|���p�n��w�p8�xPb/�i�$3v�^m��s⇧�a7��v�]��{GDb��pnR��)�.A���ԟ�䫾��7=������B�أ1g�Wܱ�݌Q4h�U�J�î�l��1�d���y�#}���"E�0�<�<8�i�bd�㯍��2�$Q�}���ia���)�6\!;�b>�iڥ��oz�� xVß�sw
p�`nd���1\�JUm���>����4�����D8I�$�C;�����@���_�����p���s�R�Yk�߽�K�8x�=X􃹼�vl���C���|H
�<�Y��w�7�nm�ϼ��
��һcAhwWg�'�a�K���5�ִx���n��s�ة`mŒλ����Q�.��n�f�����i��4�5�Ń^7�����q��D�<�e���;�0TIv!.���.���W�'\��\jY곣+�rv%Y˺ۿ"I5��u0m�1Q#�g�����t�-���L�v0�b<̯�ϖ�A�����Xha������{;�g���j���_ci���:�)Aj��ʉڮ4�b\E�ͥ��{��&y�x��F+>teNG~��_Wo�������j��ج=lh�+r�7>����d��R'ܽ ��a���_i�/u1��"v�'/x�
W��h.p�%27�<HcE,bT�X&�HV���W��;/�)����-*�Y�i�" ��q�B��C���
\�)xٞ���p{�����x�P���^5�#_Y��'�#ko(Y��AD$(�e��u�t�R�dZQ�h��[0���of�{iC�Yk�w�j�x�q��}Y��x�t�q���q�g���r]{��X�\X~6�s|�Y)Y��R>��N��{U��,��Nӥ�F��Q�N)4��yLD9!��g��G���"��ٞV1sG��vC�>�ǐx��1���~@���s�X��ەi��Ҩ��{xk�>�Hiv+w�lM�!�;aX)�0^��?S�2���6dw�?"+�~��{�(J�W��쯳���]��	>����Z+��yS�[Y�Bu�#��Vy�J�V��4�2�W3��F�/ūZ����ڼaC�$r����{�[�N���L�'
b�~z��R����仺��*͑���m�cs�v�f��+�oT�^�!`�"��˫��,f����k�ڟk���#�Wt����k;6q.M��͠{q�����"�7.��bpa�Єg���cV��t��3�
禇*kk���,�bLU��;q���Wu6����`��v㫋���	����u�ۣm������˘E,�l� z�vq��8�v##�-��o�m����&��:��<ō�lYy���`'XkZ��.���x�~|��?�����N��}�k��`Y�Vc��o��cj���e"A~�o×���Yk��9�f35֌Xg��B��M&?
mE[+��o��?�Dwy^o5WZ1� *uU�k!�+՚#WRu.��F�*�����WF�QAT��L����}�u{G��B�4'��Q�k
G`a [H�����o�"�����_a_��_`��~�g�>{��u��^�^���TϠؙ�~&^g�����O{��[d8s��ڶ�଄%y��ʻj��L����x���x�����ۍe�+O^�o�u��]w�����՜~e�SL�xv�5���\��wݮ���x��DJ?�����پ�[~b���~��>4~}�	�R����=(��YT트;x�����'+|ha��#����U[�i���a�!��f�A��h)a��s^��\�O�c �X��`A6т�[�qn��v]��
�0�n�uX3d��O�"R�����\ �u[ʆh�{K־-n� ���#YZr/����4t�~�� lN����GR4B�W�[I��?�D&äs%��!HL���_>֡��r�u�*�"�z̀�p��QV��uM\w�
+�າ���}��S�r)k$����d��E;����Y3@��WQ�L/*c��<+�x8��n����qX��<@�ڄ"W,�)��j?T��2so���p��}ccAFdp�R:$dL��}q2�wwx{��dL4�lf��w�>��^$��8��M�a�Hs��g�vA0Jb�U~�;2�&ol�8�C;���!i#2�N+\��n{���4���5��O����WwU�j^��a�)�,��h�KcPn��R�H����U���:Ƕ�{�437w������}R��.���00Y,ȋ`���!��#
�?r��r��\����=9f�ͱ��h�ac�	�	O~9���*�ґ�a��Q�T5����"*�ӕ]W[|S���w�axʻ �]��4�B6�\�W��h���5�����`5�V��5�~�� <�Pay}�]�ki0�Ez������ϟ���Z(����\+�}
��������=7�Ť�G� �.��Y�yQ_��>���G�8��k�h7~`)jH�YFw��Q�DN̬�����¦W9w�#�p�6~g�{���a���-����"����?���,���|k����+�s-X;�c i�"3��X�nYFQ�8K^-�@�m�[�3^[��!�E��M"=b?)����F�]Q"�&���ًYh��P�p��.U�B��.-*=��L�DØ�z��v6���x,�'���#��-������m��<����WW{V+�_=��E�<���*�j��+�7�k_��u�X��S���v,���5�gЊڡd�(������o�UT�U��g9-zʩ�!�V�zW�6�� �o`��a�v_��t�=�W�~��P����\q�i8ˉ��X6������N47� ���6����.C;s�?�������^�^{:#����<,� �T~���>�0�(@��dvj'��'�=��f�q������sm����e���f�����f�Upa����^6f���n-]��z������/�6x�G��ʅb�֨�Z1��;΃��KO���Ѡ��v��8��#E�!�K�wA�m\���y����T}MH��y�"��ٟ ���y~����7X�,C1�s��j��	���!�px���P[i1A.Yxz�ȢH3���A�U��+:Vԓ���m�%��5UW<�
��TjK�{aF�`M�|n쌤+��;�ɟ�pQ�q���)�S�R�;ƹ{��CW�a��	����`9��$�n>��:KPD�5�"�n"�e��{��_S�X�q_C�K��A})ݎޓ��ⴧ/��C�e+8M�5��V�s�Ӓ�t(�}F��t(����Pq{@�2�.�3ZD<z�b����A˻�{�e*:��~^ٕ�RJ�EUm�'���C��5d`D ۣ��({Mp>lF	r7 j4�r��v˘��o�亞١d��,���R��;��2v�;�4\����m;B�T�4e�����4��E�hY�}h�_�Գu�����Y�B����(�£n7e�t�\�w���+�!շ�s�\�yS�f�b�t �'��و�*D#J6�F��_	�i�)VKk+;(��Ȣ�YB��
�}�ޣJ/��W!ԥ��a�0�wf5g}��n������a ��EҠD#���!@�d�TJCY�!���ן�u�]ܙ�����u/�:���u���;kMh,Xa�N��yc�Y`2	���o}�����0i������{�M�P�Rq(���V#��b�YW2�W�x� =N��i�b����Z�gz7�>�a��ޅk&�x�z� �l��ݐ��{3�p�'m�DP7����uz�	�
2Tp��
�L,T.z�,i�"� qU��XB4d�>y�;vn�,��eΫ5�@u����/Pu��@a����D?1㣆
m��P�S���"�P�V�FE����ŘQ*fm��%���>�4�,���� ���+�j������Ğ�@��$�(� 򔄭��c�݋��iY$��Q��9;wKi�W�����'0�e��s��^�o/�E�Y9ZkQ���p׻�KJ���7[[	���H���Ji�痝��}�9���qN/+.��9܊��O uҚԫr�d}�q������'>���QR�d�ˌO6՞Q�n��ſ|��#�.G��,�q�5�p͕zźm8�u�x1�QQǎ�ۮu�]�c�wr�wj�M�g�4�x�a�z�����̦ 3�,��=Cu�3�ǍnW/]�4v�͞Cv/mE�͍a�&�)��ayn6�s��Ncv����O+0ѡ��g��v��WU�U2���*�y��O����;��M��e��R���ﳆ�C9�J����V�B6F~cP�y�v.؝�;j�!�ylv]yWZ�P��e� ~>PyUǜ���-���E!��O�~���n]&г��}�b�[����FD�2E4<��D�K?q�o.�G�q���yWTa�ﳟ�=d����������O@h���j޲MF����J��%t��p�*vY�{��:�FD"�w��U+;g�p�]�t�;�;/�7U�L'�ڗT-�/�@�:�IW�k�?�F|,�6E��m��`M�H��k@���W�C��s� �3�p�?a\���RD��U�׭WCIB-�,Vx|�?�����A��V� �;��B�6?-A,?yyl$uGP���;�Ɨ.@B�]N���H)מ��9�x���O�տg�Ӈ�W}��֎I+�r�ԽSᮻU>(�_h�Ό鄪�&N�@Y��]}�����.�C�&C��q���r�pѻ����8�����cs�+N}�I��D��Q3/G�k)a�������_:���>������*��p@@����tbw�њ�"Y���
w"%��]U~;��Z�8�M�E�J"˟4)�V�.���;"�����X�%�f]��΢K��
O���j�({j��֒�Ñ�v������g��C�6�goe�ۗZ����^�v����q^fO'�@�soֆ�4D?.��@�<5Z2�}Za�Fu��f1-2	���i۾�c���&�R��:V谈�^��������I��������b�"�x�ew��/��'�Y�l#ݾ�@Y��bь�aOw��F��t/P�Uc�����4Ir����x��#�e�ZiGN<��҃��+��7��c�1v1&5z_��U�v�M������\_���+Im·����h�;I+-��v�᫒�����:!���=z<8���ik�ĺ�B�X�Ce��]��;*�l�Z��蹌����r����?~�}p
4�3\�����}K��S�#v�hH�yY��o{t���P�������4�r�E�F����}�w/�b����TT�Q5K���op����n#�ɯG���K���{��a�X}T��Em~��dS���x�󿲐��6h�4�=7r���G�i�Pb���o�S�Bn��(ܦ}ض��fn�j�����w�� y�'�~�P�ĠI�X����GB#���  6��%|,��g��V��V������r��*V�C�V�Æxi��V��>�J�wh�5X�4�X�	�ZX��/����]<��n�^fl�ѐ�B*}DT]w�+��G�=�ƾ��Wy�2����Ř^�F�E�[E��Ь��䐻}׭��w���߃ͅ�\�4�#puH���XU� kva��-��ɴ��~D�c7��_iJ��̢~�dY~!�d�4}.ՑR�:���E��ʨ��x0Ȭ� 6G�36�4��z^����BK�e|a�A&�s��`C<�t�ϟ- z�e޹��-�L.��¹o<�We//7kۆ���hwSX�������xՖ����R���L�Ԅ�L�o������*/��`Z�:]�(n�)W�(�4E�5��Ѓ��� �|bp��sw�3���Õ��ek�Z;\��=��T�i��-Cd)Z�KX�qC�x���'�(��O��k�l.�ٻ]�h ˵~K��^���n�g?[�� Q΍;�-3�9zS���Z��y*z+4�]�2�����{HO6E]��l���|s�i���*�9��yO�c��qO=B��b�L��^��ү'&��y����V�;�4��nFլ�MX #Cʍ����zX�W�R��R�a-���`{�0b(gN��
�5\p��e2P*(�r��6��mB.������	Ph5rg����}q)�}YF����~Ӈ�>���J����_2�?|����s�� wU\����D[%���[i�{\�-�wd��&�eٲ��������<����޹^ <H�4vS��e�7�X�^�:���o��ʽ$����� .�7|���&��wD�quM�Q\:;f�Y�D��ݩ
�v5������o��N���ǡ�I�B�X�O����}7������Oa�?oc�*ȘDL��31zA�B���䐮*T��jT��]l����Gy}�f I�kާ�2�=Ucx�hc�Aٍ{����s&h�p�n98o�
��y���dd	���;��jk��v���l�tAϣM�R�b�o*u/Z�1k��4%8��9m�p����:��ba�E�o/�A7J�mNIg��w�y���@�1���V��<��;�:{�3'n���|P��շ0��}J��ht�!ʂ�8/�D|JQ�a���A�z�����(�n�ӵ���Y��|�C�&��+p�����v�B+��FRF�d�|�t�5x��d^���?���5xP��pٖ�1�5H~��[#�2�p�d\Wk�wTZ����:oܤ�-�ծDm��m顦ߩ@ug\�9J<���"�Hg�u��9�i��_�}�L~�d"<��|I���8텵�lRH׾W�iD+��ѓ[�Ԩ�Њ#ڲok���?Y�(�.�v^���7�kOU��նx��J]�o�-ڜ�%�gm�V�͚0�����[n�p"��dM�A��-�Lf?oW��>u:�n��1��{m�ţ܎ٮ}�g�b�~K�<����0���C!3׎��CH4��o,�x�},m9��K�H��b_]׻�m��es8Q3.������YD����+�R�	���A�d�z��8i��7�:3f]�1�������"�!2g�Wm�t�έ�K���!��4r�d�՗�0��Mـc�+6�)��\"� �(G���uʑ�ݚS�\-��r�,U�H,$�c|��T�t���sMiM��a��U�D��5���.�˶&�5�Z{73�M�&���Q�˚]�?(��;�4�	ٛVG�X�W/P.�i��i���j�Q}�\���O2��W�Ӹ��-�sw;
ՎS2W T�=�N��qd���g]�}w��/��-�����O��%	�u�����/h��Ŷ��C��;��-M��GY\lܜ�K%���lD�����4<�焹��W6RN���Ԗ�f��s�9�Ko`W�sՙk8�7�ض֗'f֩G|��V��̦��Oe`����'�^�v��������.TS+c�u7�վق��5�($ad����������iҭ1,�HcYD_ܤ�pu��3a�Ɍ=�ݝ|�,��p��,�o�{��UOx�QqD�&�����j��ћ�k�v�D�;�������
ˇo8s�m��F�Wx��{�vv�թ��ކ�� :ʔގ�T}��^f���	���Hss}���MT"�=%fev�]Yy��ޛjK�~�ifd�ϓN�`|+�e�nAc=,���j�u�]{�/\�gN��1���f���,xykt�U����oh(�8W����嵨 ��૭���E<�ϭ��=��=�������n0/�ywj#�3˽u�E��$���;��-��l����뇺���^��`��9�Wk*`܈.�y�3����μ���;C��c����ە��Z���ܘ8��q��mvǖNvsR�,mm86w;bi��ۅo\;Ԯa�W.i�X�\�σό`��7lX���8Sm��p�.cȳ�ힻv�牞k;�n5��=��=�pO\q��^`��$=�ͻv�nI6�3��n���y$�Fnk���C�v�c:�uù}��;۷��,3�rs��ĝ�=k��%u��I��	�{q����rg;�*�p�׻q�67,�v{+�sڈ�E�kEvP�]�=e|v�q��ljѰOb�l͎�o�&�v�L��Щ�&cx:7/�N�^�Ō��OX�6�x�c�5��l�mmٰ��ܹ�V�b@�Qۇi,��썣n�s��]X��g����Mp�4�&;n�m�n,�T�&8��4nޕ�S׆89Ӱ��k-�
�n8�s��[=qk��9g GC�����r>x�I�6îln�%��\�OM��D�v:�6⣪N�B��ۗ��D����֛x7\o+�t/���NE��v���v�\s��g��Av�-�j�q��}ul��^ ��súu����O	vʙ��y��9n�"�g�낽t�cGk��ns�<Lqu����4�񫰎��$7�ꛚ�&���k���3�.6�kO����vK�8Ÿ=z�e��8 �Wg��nΚ�<1�6��W�G�$�x�0�����šv}A۫^l����(��s wK[8��m�����[#���^}E�u⭰s����ڜ��<p�bz�9�p�"��fݍ�nA�X�u��_7YL���m�p�]pu��lw��b�ض�'�t&�[ѱ�d��+�hn���WV�;%ҩ\�������pNY����Gggkzͺ�5=<�u�/�sf��wi9��]ln�q��cErv|7nzv�i��G��Sȵ��0n9 ]�C+h���mўwl��p`ۜ*���2]m�
N4[��t��m��ۯV3�������Ѷ}���^Su��
�-�Y�i�.�X�:��=������9��mO�l�ƺ�6@�5&�̩l�'/�۵��&��@��g\q��a����O�p<�*+Pn��-
��y�9�޳`xl[��+��E�	���um�L]��3��8�ۧ-�VmG���b������DY�	��EP������aH��҇�C����@�g�{�[|����X����ˡ�m*ƾ��֬�[��?n�oɃ!$�e�$�z�*�pGw!]ޘ�;K�$+��	�]п]:7u;d	�eI�7뭅���DT���"�UT�#�ȨQ��=�W\��x|Ɋ#��7����-9��=fHŪ��@��_^ta���_QC��5�.?/��I�{ A���u��ʳ�����K7���S;*X��}��M�o�|�d������<tȬ�A���b沛ħ�u�
�}K|>C�U�Z��x�ޔ�Uм���,n�����6A�Pگh��PM�N��r��C��ʫO��SyWT�ո4����ݨg�v����=�x�9���`n�AK��p�s�^Ώ�C�}�o���3Á�y�,�7�ж�d���:��u�>�9w�+��%��+��[�
�B$RT��tǃxSۉ%7h <��s��NM{6|�Ϊ�%��H�ݶ�޽�4(�@RBb}=ʳV�ix�e{��v$ܨ�$n���6&_���p�^He�x"��������@�#�䰺�ȓ)�AE��e8pv,��0�`�Ŏ��4,˓��ݵ\ǡ�>72�3����lB⺼��C�zC��4�/�.��;C��a����A]ڍ�t��P�ʻ�Rˏ��ey)�U9�<h�����g��Di��v��}B���?c�����H��e߸?��{��w�}��y�*�4Jk2|�2�������
6�A˚���-|�n�	}��o�7�!N��=�/����dQ{��pU�s`N�BH�u���z�?C�2K���8XNE��6߮|�\{k����u�n��B`]Կ��!��댿d5gZ;jr��^4h�D}����!b��ˋY�k�TZ>�Q��!�e��2c0�cm�__���H�T���r�>1 %�KuF`�����ݎ�UC�H�'S�7�|���M�ڴݑ��n?����Gk��n�'4�ͪ�QE"$��ʶᵚ�u�:uج��s���I{%�%�c���5�+�!&}#R=�N��.T4	^�5��XUuh|�n��䆕����_9�����.WC{�v���(��^���_�~����:G���)�AFI���;��dcc�?]잒�mmy	�Y�6�Wy�)o���+�š|>����� "�Q$
=AB�We7t~�'���v����i�b��$��f�P��"��'���>-��� �p��y\�of�+�Fn����v5��£۾ٵ1fs]�x���Ƨ&��٨�&>SbA�U���3�K[�;N< �*�"̵���ԋ���ǌM�+8x��/绲�p�e*�����"�9��~������H�cd�Xl�^x^��F1}3~w�ܞŷ���_��~���-�&���:;������w2|�!�����\��+�.�5��zV���I�Hc��v!�i�(�}m�}k�b����}w^j�^���寂�3�ޒ���k�@r5J
`W�p*�(�"b�?�ut�@�=N��D=�>�&����y���Z����9 Ara˛�ޣa�;5�/c���;�M"�C�Q�n&�zqDڒNQ�J0�l�*����� "n_��r�&eк�|݀�|W܊3�~Y��px���~ྐW�m�j�I[�Ě08�Q�(�b�"������o*�a���^f�{|{�W��\��Рs%৙�B���/�񮴧/^����͊������.������qAq��8��ךk�zW�����'L��E�R�`��S�Ko;��vΙ�:�h_K<��oH�^��w��P|j="��쬣�xh��0��ء�F��0\.#d1$����nu��,{=ދ���͜*��)PCԢ��Ѓ}}���A�S]�̮�5�Q�`��6n�	��V����bu�߸�μ�6w܌G�����B��}[�1}�M�s�1�N��fΈt�	�۴v�[2-����b�C��u.�����1�"�Nw�hƌ�D.H��E*�@DWZ����j�o|�����5%�s���8򵧈���E�4D��U�e0�?2,�]��j�����ε1��g�
�S(6��!���mu�;6��&=s��S�3[���ǐ"v�"(Q�ݲ��7�gQ�"�=5�S0�hC��}lQ�	��q�I�~�[ֈhҝ�����7��de�3�ġd�>��qW���,�́?�lH� ;����������UOEC���B�rX�2)}���\~�ѯ�������	�[��g��v
���*�+'����w����6��JF"��^��F��-P�f�u+��
�C"{}���ƵY��^����Ƿ��?u�g���Dq��	�p]W�|@�žT}T����A#(�p��4N��'���0ǭ�H��qu����DZB��nҭ�@��SESH���تœkmWC��%V��෇��9u��#��P�Ik,vV��z>���/�wnr�J��u*�1g`؄{As~�;o����LT+�!��� ���>��L�B���쇝�L8a�6�R���i�D��|������g$=�J��[�ܸ�<�[�Wf��5�m^I�p0
��`oa"n(/�dgt�g;PC�;@v��jV�ѫ��'���[v��S�>r����k������j�\uJ���u�{�g�y�t �Ѱsi��jn��R;��l�ok�v��=�\q�]�s��sqr�:�rm�<��c�=��:ɵ�9͸�I'����X�T�r��u	�����r+��t��G��4ł��P��iR��Zw;ך�\p67n�D_[׻mȾt��9-��p&�7s� �UnR���ޥ�۞ͤ��Xٹ�s�/v���G�ɑ��I!`�#!Gp�^�_W�8H*%���+�Ɵ��}T+M^�?^gzV�da�t�]Vb���-]qݍ�VN1Ӻ��{�ا����a�6o/:�G�@�A���U��&�Oe"������^Ր������P�����R�x�R �L�[�կL�[�t��8��}[�����N�G�K�}𲕵g�`� n�P��K�8�@�ER�;���/�^�]��=������|��w��g?\��2 8+.��6١����t�-��a�S$����kT�+�t��''nj�0��yu������$��<�v+��hpH�h�aMWC,�2��}u���E�X����_YvM'B�. �'"���,�����O^�ܾ�� -�4�aCl'���h_V�9u.��}T��/���/M�;�=u��T'�ME}A����\��ܠ�Lp��(�`����;wn�nۖ��b�7n-)�xz���ۀ��-�������oG�u�������(T�CE��[�k��!O'JW��ＹV&�3��I���~m�y��DBK0��zrM\,B"uRSJ�5Ǐ�f�f�zk\�����;���,�L9�-�}��h����PXv��C�=�wM >֩�jn��>|����Ὤ�[�힭���I��{2Lӑ�e�	�!�����u�7r�h��@�D,޹>����V]=[����GW�>���G�l�q���u,6A��W۝}�x�tTNn��W�0��~>��6���[��k�q��2�����F�\�&�oMF�"B�mH/c1<o)F�����n�)S���a�٦��gt������Z�������A�'��]י�̨�.�v��]U�0$;oA$x�'Ѣ#2EC1��$Ut���Õ�!��;�&b����K�Ɇ�B���\��L�� k�b���t���hTuc�u��=�Oa��ԁ?��:�U;S�ێ.�v��s��<�6&�۱�xW�
K@��9��>'
�_e�0{Ϙ�z}���1�P���t������ "�u��3|��I��Zp�r���&��2�tb1��~F!Ŵ�d�
;+��Q��'�J!:������WZ�V���"�Vg�X�C$ʌ�_WV��̅wUZ�Җ�/�+��y%�6K�^�v����
�Q�d��ڂ�����M����cY�WVj�xVy�&����{f���CM;v%X9��m_�d{+A�(_�x�$\'�s}�����/xjs��?8�^{�c���<�Gzk��P�;%Fȗ]tK��}��;}�Z9li�&ȃ,O�m�ܗ]�i��E�u��{�^�����اsB�\�v��y厝+�D4m����~�B��4]4E�s�]\���U�YD�
�܆7�P��bS:�q������`�fF:c��K�zxit�m��n�W�?{n�k�T��*�s�/DOPb���WVC^8B9Ys�5�~w]g�ٙZ4y(���eRV��5D,���n�[ۮ5Vzѩ�;tln�5�k��;�/k��d���d�l�b�m��˜�Cv��kS��)��C�Y@߽7{���̝��𡱽m��XB�Z����u�<����m��x���	 G��Fe/A8o���u�׵u�Moj��m�� F�p-s�X��8®oR§:�mm�3E�U����gw�-�=r�P_<!(Y1$���2c4��1��]}�t��l��`��<�Ӷ��6ދ3�mze{��?t4[5������;�_�Rr,9+�*�n߮��I��b�٦>��c�r�X���W�=Tw���� ]�m�>�����Y�Ӳ}U}s/|� �|�ånB�;�8Hr�m^������k�i�R�v��g9�j����5�w^lY��/�ex1�6[��v��h�k`�]�b�k���}d{��.q�E��P��e�࿬��z���{s8�ي�U!���ٸkI���ɫPُ5}t�˺����\�YEG�w;��� �s���^=8��7fz�����R6PøS۝>$#]��v&�tsc��ä�RM��7nn�D�PF"b Dۇ�ʦ4~w��Y%�ty12�"q��{z�/X�rE|{N���[�ʱ��h���P������:�p��VbD4���d���6�rvdڥ+�n����1��5>]�h����@9~�����ER����P�lҠ���k��9��N#t�vBOK�U��w-�	�u��Z"A��!"73�#�u���)�{�����3�/�bu��=O�'��D��,zwu8%���;'>�p��yg�	V=���`�L$�q������w�}�iQ�y�gd��1�$,���ͥu��e�o�UX�3�|�#� �9��{���?ye�zKypx�j���o���H�$�G�p�-;zu3��?��Ofeߦ�L;���i]_&ݕ�Z���{�N�T*�������Y_vv`���",?R�>>�o=���{���[�Է�t}���r��5�8�1�z�SA�H�'3tkX�q�ޭ�w,Q�nҝx\U�G^��}����q�Gr᩷2\�֙Tq���2з|d��b�t2yGcn^�ޓwRv�z��n+c(���w���
��W<a��.�vG�zzw���]d��b�g���d�q���W�yL��	�^N㎰{\v����ur��m�<�m��\�U#�K��HV�m�8���FY�ɬ�N�5���耺�;s�xxҽ�8�ۍ�uϦǣ��;X��7Z��d.�=q���m� �c���.�m��e�-F�p4wHgΞ|YuSv�Fܸ8���a�v���˂��8�Rw�~ο�����^�դYD.=�ٙ[��Ye��.�`�rs������9]ݲE�_��o+��{$&�^ʓ�[eQ!�!�$d)��(���E}{��:ڱ�~���
�HK��j�aR�<��D��Ef�Vm}���+����i��+1_+�����y�nO��79���be�
��ే��;s]��C~#Z���ng�7�w���b���.�Y�������p�~�Qb��G
5�A˩^��\�
`���Y�Ädr�X7�Tc|l�s����l��^W+�暯�!i���
C��#c�PH�_�u�UB�%� /��#Ϲꑗ!0ai��x4�Qxʻ�!5��:���q�(E���=������_o��~B�O�=c��΁�ύ�Em2F����Szh��.T�e�q���L��hlT���:5��rF7��D��/K��+��۴i�d�p�����}˻\���Ƭw�����ꆳ}������[8��C��1D�K��!��%\�<�^]�u߫�����#N�X켦��d"�l'�a�	���Kfsh��	K�0��<Y�-��=����]��5f���t��*B�x*;�v�I�M�Cά��1`��"
�w:�`���6)���=�Y@Nʶ�����;a;�]gOʐr15�Jq+P���p�wl��U*&�����> ��Ν��^�R�*�&���t��dk0KP�jH�Y�EY.���={ҳ�����$����~G����Y�^XJ�L�����Ӄ3�A�k�u�mO�J�1����P'	*�N:Kn���_��ȶe�zh�w���a�dA,�Sޕ���R��P{�-Ww_٣0�.��~�n�ۓ�n�&���'��:Gr��Q��31�{�<���=�(����h��z�"?IXȔ͎>�`�W,��R@�G�J�����5z���ocϻr��*�2��P�{�Аme	D7�4uv�W�״��F�T���ۮ��q�:^���QJ�U��5K����/G��{�4���#^��GՑ����}�(תx]�N�ޝ^]��,��f�$�f;�X��t�!��Co�`��i�n�����8~���s�������&L������E��V��S�l����u���>�T�3��f���p]s����XV��(Ў/�h$S��^ �nw:ux���@��D����Rx(����wEg���ֹ|riK{!�'X�OK��|w
�^:�^D�������$��B�:7^�h�9Å���{Vp��Һ�`܅ۀp�M�@��մx��Nj7y�.gc�O^�/�`e���t�o����g#}��ւ�B���{�Avm�dM�+V�$J�t#7u��i�	n�V���U�����ӟ&�n��'-�D���W����f�̳m��-m=5��J��I�Hs@�<�51���ϠV2�[�I5ٺ�4r�
4o��ܸD��/�:rAV���ħ�9C��7;G\�����5�]����ߎ^���3���#"㡜���ff����B��Q;XQ�}MV5��+�`a��U�=X"�<���[Ę����giZb�ɓ���&�������j]����zb�z��	6;{iQ��m�FpY5�wA�/1b0Ee�`��Tbb�^:}r���],oh���)�lh3�<0�Y�7̔��+�������y��Qs*����ѐU�oNF�5&�N�h��HC�%��M��r��\�/9��E��i�zz����d#G4�������z�k�+�
�@ڜZ�ER:6���j8,��;1ϯݛ\�ܙ�'9��&輮��3q��㝵ʶ�X�N�t�L�"!�a��jm��]v��ꙻ�FřY�;���fN}�v��L{�l�'��f�B�.��eJ8�!�nn���0m�F0h�CA�u឴�#ȭ�����=�X�eVݡ�r*�
Շz�ۙE��T�lS��kƅw]���Y5��*&�q���w^b��g�m�Uݕ�Au��a�@c"8LI�uu�o��}�sE[L�Jy�u���f�@����wƻ`{JZ�P\��[����Y��h40n����~�u��"�� �)$�I��!0Ce�u׼����>�̍d��ȫ��6�$���Of�OWیƬ׋�v���b4�zLԪEm��3�qgۺ�H����=�㊜���u�mV��]�Ǚ�ӷwN�M��ų�Go��+��@�o��N���<<����l�,І��}�/kZz/T}�L~�k��
C�gPYF�S��ׯA��	����#V�,׵r�6�U_� �l��o�ǴG-z���[�U�Nʏ��Ŏ��t*���B��T�N�(����蟙~�3~9�Օ�S�FjB�"�:Gc���ժ�`�P��v�^��/6w\~�|�R/��z��Vx�J���x�c�Z�C�WR�=�B(���+	��]��W�u���q4r?���{�Bq4|/a޹�8��ױV�b��>�W���m죦Ǖ���̹�(�MK7S��T��5p�۴*��1k�2��r�f6̲h*�\�㻗��6����m\�J�Ys%��,g���nL>ժ�Μ�"���"���n>۪f�F�)��2�r$�p��ú��+�?<�s���!�Q��5��F����_o�C�|�x�ol�c`}X~��O �����ېN_2�22�7[x^|�Y�	���Y\����-�����<㐷�֍��*vͻ��=�x�q�a�li�v����~E��,��_����#u��=�t�"�w���XBa����fu����]=�(�CK�+I+%p�3J�<�D�����%#_4`���Ow�M�o5RY�����Cp�_yu���9��P�n�."�+1�Y���NזIA�vk�g=ݜh����ZW	�]�VQi<��|qQ�T�)(� Y�-���\��>�[���Y�V�&���->�Q��u�^�&�܆�kDyq�-`���-z���������4n�q$�A��qOYcٟY#'��E��u��h`�5���r�P�a�m������Pd]��VM:�+�h~E|;�����M�!jHj˼u\zM�'-�k
CQ6�W'G�%+�e�P�aV�ǁ""�����C]���!�h�V1`�wwOF�̌�,���$�=�+E<5췆�'�/&��y=8m�e��@��,4E��0�3�*U¨J{�o�Y���=�*�zC�.�Qɧ��V��Kn1���,M<@h�P�������tK9����Se��ۋ5��Ƃ��{YPS��Q�מ3�l�V��v�������zN{w��y׮�#A�b�`��k��X�qms�����M�6wan�ݶ5�:�<��{qtr&�n������k�9ȉ��텝%��mv�i�7a���3=�3�����hݬ��@r�C�Vb��m��e�/ɢ뭋�1���7k8xn{#�=E�;,=�<p�t!mr�iz5�da��w�LM\�����0���� ���I���k�=3e{�)Y�wK �U���ډ��ݶ���w
�/e�y����O���kdc�Y�m<�I�d���^�ܸ<>��L�tt;���7�!�U�5}�m,���!�-�C"�[[Wu���2_��5f*����S	눙l��rK�;#�u��	�mԵ�Q��2������T2���/zq.lX7�Y�tf=���Dd~J���gtg}����ek;�B���D�n<��p�l��Wc-����N�V,����R)�׳_�ǥ���>Ǟ-xeH}�9�}�����Ω�;ۦj�5�b�kل<LI�GFG��g<�]�	��o���s���G��K0zS������{�]��x\��:���.޼71OT�t�W/f�q:�:�1�RQ��sn��OmpY�S��p�n�:h; ;��㊲Z�>�����V��[���G�?]TƲ�S�ǧbn�5ʳqo�b�{��}TV��-�G)\*�n�</27u����r�:�5��M�����ѹBf�(�V۩�830G�{�/���<ƎD��;Q�R�Cb��7,]u��0nM[:�
�}B�r�xȶX�c/xl��l�۹�r����}�-.�=�iR���ݬ)a��MPs{���v�AQ���+��?G�i��bo�ߵ��d�J~!NI�)�����9A��v�쮥K|�*�1V{F͘J�v�Mj^�>�u�(|�-v�ٻK�7Y|,ތ0�E�щI���.�=��Z�)�zQ�9�+!V�f]t�lPۚ�J���s���e������F�hu?%֫wؽ}�Bn�Нg4���Z�n��Mt[��Z��sY�-��J
7��=�����V�{*�2���=~��ㆃї�.\�z����3v��/E�k�I*���5=���I���z7���X���܃�3��\[F"IH��ISv�}�74������{�UG�����2��q�J�5��B�k�_@�ϹOo���g�A�u��\v�]����,�a��"F�k��*%-nV�-�7��+��gV����}��ޭڕٴ��P��m�un����ૼ��;�� �yN�HG���7u������=M2�K��P)9f�~^�yhN����Ϛ�][yj�
��& �Ѽܽ��y�9e���O��FOl�%�᤺���`M<x�I��Y��,o��n)o]_��]����b�k��F_�Yr�KT��%|�z�}�F�xR�}:�4&ZV�M5�#N<ϱ����3�ק�;�jU�B4��vt��d뺨�w;�+nb�|�H��ezvXxrZ;���(Y������8��.�]�R��x���Q���۰臨AF�>�7�B�zѐmU��c̬9��L��uQ���~��d���&q��eG�	��cos�t��:
�Ik���t�/KX�`��q�"(BB%���������;s��z��6
�n&�v��X(���yW����]SC��h��nzUe��*����{(5;
�
|P��s���s�R�����칃�y㜺�A�!����4�f��y~��"q/{p�
�����oR����<jx>G�Y��;�]�c�ܢ�"��xon�;�{��⼌C�Jf&D�{��[۫��'�c�,��cU'�2�]3Yz���v��3_3���G���r�Y,��?�@]���Au�)b�Wy��֜�{�P��yLC%�Y�]·�<����7�lP^�j�3X�.�,n��U�t2����\�fE��&�u����8(��囻�AV���,�w�>����ֽ�x�ڙM���V"�x����KC��g}�(P"L��qk'ݒ���t4s�ծ����e��`�e�}�?S���5���58�����܋�������&E�h-"��"a?�E�9u�O]�v��u�����w:.�����<�q�v���9S���������o��y;�sgM�^�^([sʩN��6"͝
�x����W*^���[���BHw�U�&8���!�+�XEQ���i2��۹3ּA�k�t��,�c�~���C<����Zr@��vC�@������Tl������  M� |S8�B�E�v�ڳ5��wp�Do����=u����l�5r���GlW�}���\�6�^go�6���. |������ݭ�������G�����{���.'G�G|�Қ����뮋��h�x��Z���3����o�7��	%�˹��>4à�h����UK�뻞^\˵@QAe�~ʎ���O�<��/Ξ���Zx����ï�Co���#�n*"�7�q=�����P�=B�d�`�J���ݗd�s���3��r�����EvA�ҳ��r��fY�t�	�n]�������5�H�΁����B�[Ci����w�kN9����8'&�U�ݹB��9ۑۻmصkQ����!vv3���ו����nMF�\��u��h`��!�gũݹ�)v퍸���[����#�(fB;N��X�6�o68[���5�4�@��N�X^�;'T>m��֗��:@�7"�����8��8̝�lm�m]m��29�nny�P�����c^5��r�Q���=^�=������m����ocn����s=���L�b$r9;�˺�yu�҇�;���$��ѫ�<�T㨧�]�5JW=��ho3�I��k�zw���A^���� >}�	l[.�L���#nk]�vf�8������GHu��7<O��2�Y�继_��5���ה�8J���&�j���T�i��#ӽ�oJ��A�**e�7��{�H����w����<�أ��}��֪���`�.�۽�=a��S��<�]��f?x�*���y𱍷����57|�w��=�}������:�vs�y�vA��e����i?b��Y��=W{IYHcq��zW���4T�[��$@W�e�Ow�
��UB�Y����@��b-��?c���Q*VpU��^)%?kx������5a	w[Y��9v���=B�NBb`�I����+���Is{b8�s����(
�f7n%�&��|CaZNEsiQV�r����5���ə�{%�z�[�^T7�k�L��}��ϧ|(���\7ӏR��*��B���Wř"�g����g�4��WBoVm�heD��.���k�>'w�\�O�׬k�u� gr�-�+�X�b�:w6:�r�滕����q�Nok6_oSi�A;ˆ�7J�[�;�W�̫�z���ו7gh�
��=A�9=�m���oWb�y�X���'������J��wOQ�F�`�(�(�x细�#:y~w� e�eS�c&�6�\ʼ��T򪩍�0��b�0�*8�����A�'�w^Op��j��w�G�9�_:��p�Q.��8��OY'*q�V�ۮӲ�β�]pdP!�u� m�AFZ.Ay�doIy���*�A���Y~���7U$���Q���8P��wKw|�=R��ÙY�)!�z�I�����T�К3������<y8��\nH��9�׌ �Ν���ݲq���Mn��S�:�����,�ޱ�+�d�lWmd���CJ�Ƅ��o�/�mz��)<��*��mǲ���wAE��T�����ɡ�H��(�i��'���H��n�~Ę8��ů��z�O�%���s'����T�mp�q3�50���B�A�Z2&�l���ʡ�w�(4��M����m�|y=�צ!��f���"�j���Z��2����V�XՕ���H����P�ulm
�T�[9���i3[�7��M��Vùy�#���˸��ΞζE�$0P�	����UP�n�ԑ��D��w�܆u�ܡ�����'|�f#�Z}�#V,��F\�M����xl��__��;�%d����Y!����v����~�0�.9��f�c��j9�6xk��ٜD��U$�����������e8d����+�}���nvػ���]�{`�����K�8�x�+��=�������T�'T��Z$��ߕ1I^wۣ|2���s4v���9;$&緝,:�{�L�òo�Qg{�Z�Ժ{��h�35ղЪ֏�!NRQ��M��9M���<�J�V�W6��K;b[����	{m����\�/<WYi�/�����s���Gw����ڇE��?0��"VH���M7 ��i�F_o����v%糽��m��{���g�bt����62��^�5d���L͔,>��"6��'v1'4���sj����]��Z8�z�e��F7z�gU�O{Sʷ���P�^we)�����Ӄ��tqD)����O>gUMN���j�T�2�Sj���_>���$�D�
Ü��,d7΅�tЎg�vn�ܤ�X���;�d?@�9�G ϱ��S��|���)��t�֑�-̓�3(�=v�ޝ~��n�p��#�=�������xm�sʹ:S3F�ΡF�����	'�uv��+l�x-�����wС{F�h���]F����`�𥅴�������.��=�r�۹�J!�C��~.��d6�0xo42���n���hiڠ�<���thy�zE�E�k���9�r��G^K_K��~����ѽ[(׳f���cڤ�Sk�L���S7�����#��-f���ۦP�x��^��� &8�%iә��j���������8�v�t�8^�|�����Cb�X9�1y�|#�Hh�V��q��
}�1��Y�A����L͋���׼��Y��>ֻTP�>�6�}K9���¤ن�����N��׽3���<�sZ����@pu�H�]��fƞ^�����4��]��#v6+���>����̞)͎Vڣ���=4sVr��9\��s�pӚ߹Kcޮ�� �ɖ�<�[boTH�%��V8]��a.Y�7�d��W��M_�s�=���w����\���]� Ϡ���x*��s3��>�t�ݕ�i�Y-W��1�.!92�H֌���gnS�S�� U�Θ�=v��R�N��u!ʇ^\��..�ui�;��۸�$��ӻ}OP�/��q�Ge��Yݩ�ףh4\)^QOOi�/��w��8��r}|�d��G%��)��.f�c��h
a��4[��A������^�-�z.|�Tr��5��B��Q�_qp�|���^J�f�d#�4�j=r,��ZE����\;��ֻ�݌W�ޫ�Ucm�uWc
�pY�Q�����׏1�!rˮ��H�f��r���qƍ� r�suE1����W.�7�vh� �xW;�z�q�Fѥ��'VEd�w�� ��;QX�!�ݻ�:yT+�r;~��
�1��Ss�]�;�v�4uX����[���2���K�Ѿyi���9\t2�����W*j�R՗}z��5{��]�(���� ;8p��E%*�v��d���f��"��۸w$��l�ȯ��U�%��w���	�*v�\\��+�ꖵ��keg�u���ͷw��
�����`])���u�����/so�\F/�%,ս�5`]��~~���nU�(�zT4��j�������Wc�5�'����K���m�����<T*��O�g�Ņ�Q�B3W�� ,z#�^B��x�5�Ux�ؕ�m����7�u�&{/ͬ8�#%^��U쮈�nȯ�yN[���(7Y�g���Ŷ��ۺ_,]=�lnV��z^�!�4#E��^�<����(v礲���M�p'����ht.}��������4b��u۬�%�Zv�y����z��v������m�A�#<�6�v�����m���	׆n.{=nd.�1k�ol��a��@,�޸Ab�1z_nƭ��
=h^#��fuWm��^{�L�X�EI�t��7�:)k*�Ҭ�),�
��l��n�p�����g�]���G�79��ڛ:˹{Z�i�(��Ź�mgv���p=�,:v��ڣ�{=nc"�\ϖ��6Z�&��v�iUue�3��Xt���f�����5�k�!�c���zwh��F8���V��NL�ev-�6����Y�a�.qY�������m���Sbg���y���1�y^S/��g���t���lc���l�qn���%�:g���g���l,����n8*�nv��qgoj�ў�'��uqМ��f�n^�O�	�c�nj��m��t�ӮC��<��xۺ��iM��ַ&]8�w��x�\�n�D�^��8N5�1��i1ѹ�<OY��lsƜ�qj����g�X:�N=.��K���F�p���&s�9m�l�(6{�@p�5�:Cm�.c���6Ρ;B�Ý�H	���>sm��1jG&7lr������m��8��q��w.<�Br�ڇ��a�����q'ti9���B]�x���n�����'�����C�2�Y��]�7a�Eݗۇ,ӻ���ݰc#u�Xݜ��M��u���h�]�i�99z�+�A�i�m���gm�%�ݙz=1HΊ��n�u��w��czGe^۫�K�n�j�kv:�`ǌc	�*�N1E�d61ŋݸ8���V���ױ�㸸9�Jr{]�W�&.�d�s��6�δ=����[��������cg�Tо���Y�
��˷oREr�[�w\��T�{G[q�J��\u�g����6�V�/'討���nuc��j�s��-ǅ:Ƹv��7���|p\I�2��v ;���k��0�\�%��	ɞ���e��-�-�A�=o7;qw<w9��i;�%��zp�;�7k��ok���6�퇖�eیXs����Q�l�+�cE��Xqm��ݷ^M3v����;�:{u�s��n�F;uFWM����<��cٸӶ����v��Rc�t�����m��2`Y����ך���C�D��8�I
b8�
I�Q��ီA[�W���n�+:�rx9�Di/�i��-k���^�� �����Aݑ�zm!3'�Y���G�v�2�@�%Z�]e�̞�J{o��7�Xw1�Ƞ�y7J���y��Z�AY(���:���_%���2�v輗��~	��D�H8`��<3�'�hv�pP�W�m	�Q`�F6%�b�_WJ��Z�s��{��*��0eѻ1ȫ�6���������I!P��m�����Y��Б����n�������6��,Y�7g�C(of	_�����\���]��ڽ��ΗTM\��Ti.iHHB5	r��ҽ����EWbƇ\�h����ܷ���,����}_eg�v��{p��=�V��2�eogL#S�,��ݱ���ۜq�$��	�t��0����N1��Fm쑎��sA�
-���\~��W,�v�ENrV|ˇ��1'�ʆ�|�z��\u��+-���/���TX~�[�{�WyY�m�T"7m.�5a����V��S&Y�f�u����篟Z7��]���PĤ�˫��,R�����>��e��ta�� ��q;|7�����JS�f��A�ip���]�<}A=��bN���+2:�O�=Ղ��Eu�"��B�L�gp��P�ԑ��{%t�wDxI���yO<����9���if����VC���9�^3=9�BU7¼��2꼮�]Y�cP#�qYnюLXfJ�Y���=[x���3� �w�6������-��}�IV(�W��b����d�-x��\n��4{��r�쒁	\ǰڮ�5};x��p���<6��=�eqIVN�t�WKO4���^V�kc��]�[bl��2z�ʼ&��LH,��`ѐ�����b��4�E�Q�4���tG����L��P����$���~1�C~��Φw��<a]1T�uR�{�jw�zX��OlZp!��O:�l���87���/EI@��I�c�����}�x�ｑ�Jƍ밯�H�����Τ��;U�۴_�/�׋����{����f�o#�W�14�@���P���Z2�܇��3{i5&���^v.��\�Y �����g(`ʖ�칪��sU^�˱f�g�S��K�{��&�Z_*�B���e�֎��c� "V�]�8:�vS�c�.$gi�z��<��v1�yP�}y:Zx�a��^젍�B��A��p^v���e���z�����W/rk�g��}\�4{^���*f��c[�|�E;k�M�Ӳ�6�FFɂ��T5��Y¯��X��T=�(���G�v�t�i������{�N^�U�b��y�z��,��){�������F�u�`�R߈�c	k�K]����\������Rx�qu���n-g����aܵg2���Ԓ��@��D逸�,�ܖGsu���%M�:��ly�ӽsҋ�~��UՍB�|I1��F�y�z��Hx@���,uy�_E.m:g����'������*q�iKD�>�n@ƶ���<k�V^y�Y�:F
L����EePYӜ��w��*��;UfK��ۺ,1����6��"Ry*+����^tŞܺg��M�.��f�ƗF��" ��� ��׾e�t�����%����]1g��
yzr��������]#)5̷�y�G�V�B�&�ł�%�;(vn.�r�N����z�F�L�q�7x��r7�G��kp��_r|e�}\DOO2�՗��SA��X�bG�F[�Ȝ�i��WH���T~~X���W���wq	/���70w�^�J����~��W=b+����6��^��e�Yy�8�ֵ͛���i�xh��8�ES�n;^��Б��n���n���Rq��v�^����V�!�b[�ީiۼ4wt��ݫ����j�\
�g`;�a�
�.�܄��*wU�u�BT�p{E���FK�E %I.|�;Kq]�<�Ҷ�^��+\^9���3�oR��3��̚��w��O�粝̺YռwmJu~Y�>�F:��TVrrZ��G�%9N���eA�K+�^�`��n_8:�s�&����#�V2���.'[���IG	vh�`�p:=-�Ҙ�?$Z���z��)籯��ɵّ<{���ߦ��YS�b��&Cݞ��L�[O��L�[�=�XCʰ��9��A"�Фr�n�^3G�{��VV��t��8ޮ�Z�^��V��K�u�g&�W ڝRd.�b�Dy%/{$��->ynEע7[���׹.�0Z��Ñ^�C�U�k��;����R6�2er�B'��|���$T�+�T�M%`���E�?n��㝵��l.t>K�ַ!\q��y�7�y<�f�=��Cj���kCtv`?��~�彷O'J�=���a;i�箃FP�+��;2۱Ƕ���,�p\�榻r����ֶ�k$ۑ�۰���HSƍ���0a�l�Q��Ɠ��)6�2������N� /[�Kg]�\�]n�e��]�4Q����vx�ݶ��v�G(;���\�˞4��p�[S4ۧ���BѶ6ps��wk����}i5���?7��w^�t���ժKYv�MyK����VUo]�4��}WYW2�s��id�Tz�+�v.��3C)f�!gK�	��\��v�{�-긨��N��/=��un��f��%�Kg�nE=g�~b�Gyv��ם\��&�^�I��lh0(!M�1H���RB���qK�s��E>7��Vy�T�U�+~�0��p�n^J��Q�����R3�U��\p�	��ơ��E^I|[زz5o�dɫ��x,��D�^��=�\o�*�e��ե���T���A
i�_p��#F8NC��*�3�*��'V��+9�_z�A��7��f&'�(i�"�2�"�v�'=�b׏�z�׆iy��oĽ:ǹzYb�yU�ޠֶFo��`��6'��kə:Sw����]�m��c�-�,�1|9`��Q�}cN��W�%d^��V��*k]p��a�W�g��f���\����\���:z&�(Z�X�ǆ�*��ó�����	�<�>��=��i�gwؐ�e]��+�\�ɲ"҃�i7[X}e��w�v���`��IM�
��_�\y[���)�#l��X�D>Wf�H�㔝�rB��~���`��W"jח�7[2� n_��Ly��)��瞋�=�1��%Q�����3/�2�6&��W.w�����D�,��+3��H����뷏x)z�jܽ��z5w��=�)��o��H�!�@�Q7��S}�☼G2]{K,n�M�vp{8u�=�+�r��)�"T���$�������snA=��M�E��q�30%�S��y>��~�R���fC�3�����g��z�Y}�pW)k����w��WIB��[�|}��n�ڎoG<��s�[lK�2+��]5ͬ�wW���s۱��`ڎ����"N�Ӳ�9N'��i\^�j�]{9����������z�?-��h�b��PWS����+e�P�1l�w�-�¶�Cm��27#�j~A��	�]j��k���o:<zvwU\ݡ��`��?Ay*G�&,�����N�׫�f��3|\\�9�ra�^��e $)�m,c��[��0�7��h���bp+-�e�t�o��W��������/�h���b�u�xr��9�ݠTE|��D�7���h��Վ��u�q�љ�2L�-�W�����&S���+t�~��QQ���U3��GB�W�H�@�`R��'��.�*�$�QE�����H�g9.{f�7
�����r��х���#��1Æ+p���^w���Y�u�d�ھM��������(�9�&��Ycw{=޸�j[��i������X�]OO\n�v:�x�|�Iqϝ��Gq��]��m��9y6:��q��n�@"�w��2�_5�a�z�)�����)8ӡ��>Y=��#��~��}\M�3E�ƅgnLeӛ�-BAኁ�
��Xb c����^��(Z|	KW����C�e�^^�h;c,�~Ww��3hf���⽆���L>�����Lr�����/��ĩ��XӐA˺tC�Yw���[�q2��&�W�<�6���c���{�/ ,�NIRK�~��>�*G[�n�P�o��ü�[�T�������Cʦ죓��ܝ�^�..�R�q�9&�4�&�W�%��yBf^c�wWCQ��̋N� 5X��ԛ�6ܨ��t�pj[\f��];i��ƴ�p,�>o�m��x��6�8��.��H`�//32�ʭ%�תn��A��ڂ�7~��r��\�K��X����=�o�������-z� �p���f�Ph�˄��(Hۭ:�l/^:̻d:�g[�C�ӓ��\��.�f���DA)�u�b���}x30�ͩ+���nj� ��~3k����~y?l+��f\�i�Ͻ�V7�eO�1�d!7���n1�����%t����I��T�v:�}WXz����E��a>��YȮ�S^����at�ځZn@B-�	ȯ�x�=��R���eAAz����|��+��K7˴���aLwє���Ww�F�t�ޣ� ÿ�1�NL����	����������a��ʨdwUa��_��Ƴx8 c�A�}(��
��mzg�2i��y�?B�%Ɣ
0�pײ��9�f�^����K賍���V��Oʺz�]�^g��RV*c�{���4ȡ�{�v)޵�I*cý�$ģ�U����>��4�a4qU���.���X�-�C���[�wۄ�G4S-���1�ڮmް�*X��vռ��Zu��U#U�	���v��ֱ��z��g<clmv�tj����Z��Ivz�9{��x�&�xl<F��ͼ�uWlN�L���m�y�6��NT1��Ӑ��ۄ��3�B�����xT\u��f���"g^���>׷��'�n�:nw�gJ���nS]� ���. ��[��uŻs��;�\��pGg�����'>��E�����E�8�:0�v�g��Vph�5=���Ϲ�iX69ݴǼd'���lޓE�~�Uݚ�������ak&����myʙ,��(�Q�mmau�Z}��L�S~W1_�6�p@�i����G�l��0w��^�uԞ.�3æ�u�=jvx��T� <ûTq��IB�����Xڨgk��a��a�^�X����6�eXƜ�U�=��4^_o��˂�Zˌ������o�|�=��\��+Ơ������Z�3�Q�ĠZ�A$Ȥ����׳���h4�vei�]g�����s� �s�"sԚ�N�}X)T;%2��9l�Ю[�s��@�jT�)U���{�@�^���ݐ��;�mA�YS�n{�+n��yfw��l��3;`hWW�JQ���=	K��Ӈv`�O6�N����s6�6�`n9���Ύ&��S��h��o��Y�30aO�鞥���,�%=Y:�zT(��;�v���wM��đ�b
��W��Y�[�"��!���)0�	�g�4�fӔ3ޒ�b���æ���H��n)��*� �I�+\��@�%,��FC��j��Aj���#˙jb+xݑX��IZ��wWt�L���>^�=*�HT��{��}�c}�kUҜ-:Η=���8�:��W����aX`p�Z0(QR3M;�ނt��y�4�r�W�2=�]S�aD�=�xmɡ�	��N����z�赃�w��NA���V��ٙ��qJ���������BlK�n���'�v<z�����]��V��]����ys�'+��Q5�k�P]����7��"E	�H����]g��Y�B6�7D;�v=/�f�����\�[ЛuwL���=������)���;# �$H�Z(Ěx3<� ��csU���`.�%�P�������7=��
q4��㒫�h��Eu\�$��g�d��`�=�s���wM멑��G��)���x��,(�&�Xó�R�z�q�nJ�����nx �-i�
\�շP��G1G�����]�0�_���G��6_��(3������\/+����?J��G{�Z��|��gnsÞ�s2˜cWfi�ٚ!V)�7��^�(.k<"�W����ň����}-���rᥝ��
Z�����tzM�c��m��Ɖ���Ω�]�U/rc���o��ܽ.O�gr�e�ki:�i{3��h���w�Z���J�i81;�]z+�K�/���n�N�S,��h�:L5)�~��'[c%Oͽ�>�brX5�myV�,��Z��\v×Sc��mväK�w�c.]m�y�~LLշr��B���8z�X�0��T�i�������E��7N�a�6�
p��[������������x�7��G�k|vߞ��G
^��6�%t�@�x>�έ*#n�G_
�#�C�iIMЉ�/hy��-�Dߕ p٨���J�%��f�FSu��C �Y�9waT�Z����+V��<��\�;˸� ���93	x�5�c#g������l�3n����.�E
����..�s�G,�:�]�����!��W�v���3Qݥ�Ƶvf��������\Z�e`��p�-Pj����sm���ݚ*�@f>�r��2�H����!h^�����
F�HV�7���!��k!JǪLU��Z:F���*q+����^��c6�>�,�;�(�N�e�C]yZ��gM��#O\ɛ�<�tW����!����{S��ovb�Zp�N���]��	�6��(_s�s3-�t�=���%)t�FM�t�������%K�6V�e:�f�'��VtW7���4�ئY��X��v�m�/Xw�+��u�s��wbR*Y�1�2�83d�.�r��������F��+չ����{f�����}�פ�� 1�^���G��V{	���(���h��eI	�=o�:5�����_��:��*�MZБu�x����R�1-�f,��F����%{Z����{������u5$�R޽���6�I�YM��Ή3��^.ɺE������d��=�-fz�۳�9W�з�&�f;�致ϡ�n�u�"�Ξm�,�7���4������jؘ��	];����o�����y��B��_��)U�������7��r��Y�Z�3/q�u��-䘁R��୩��<uK�rh�X�V�Evg��_�ć��7�=w�@���v����c����w7��h�JhF�q�s@������G����[�T���۽��V�]�+~�T@���@hoA��w5�N��[Ncr�3]b�5Vd�W���=q���Iv�<�Y]J�=�v�_��C�H���{�r9oi	�0���F��	�
(�$��Ϙ3���fڨh��eҼ��J�^�O(;斧���)3�}|�u��Yd����=��5�Z���ol�4�� HU`�AC#���Q['�-��[�a\�2n<�pq�[�B�p��.C�σ~ͥ|��9��]�q_<2�jW���z{h�Ɛ���<�����J��txZ���*�ɔ-�HFJIx�U��v��KźXTݠ�v�Skh��gY�e�rd���5����3����4�$�ʖJ��m'�	QC6ӌ6�Ǐ ��-ъ�¹��z3�}A �>:�ԝ֛Ѻ�/;so���
v��\O��/)}����&B�QT'PZqq�U�Z�׹wƏ&��3I��Q\N�Q�|u�}�mu�3o/S�4�ڼ����;k���4��!�����C
�� P(�^�)4}���R��\�!��57!��AȬ�;����k_,�>E��тAkH�K�B{�����rڍ��B<v��9��].M`�����kY~����{������eݫ�8�J���-An8�I�fw*,�3�;9<�;�r��8����pv�����4���?rZ���u����7KŅ����+^Kt*�,i��{'y�m�K�=^JN��훍ɷA�����C�/�r����Z�g/��˺�c��w'P��sC���V˴Z�E��λ^ݵ���;n}��*���^�k8��9&W�v.���d��v�3����V��m*ݢ�r4����t���۶y6�w7b��Z�>%;ED>}h��鳜���%[��J>kv��+q=k� ��M��hW=N��?~~��}���.>�wAÚ2������-]-}h�{���*�9��$���I֥���@�bBb@\���K�r�zf9G���
��j\Y�u�g_����W��̹v�_IsqJ�<�m�vÌ䭴�X��P��"w�EF�RJM�o�^��{Ҧ=�b�6����P!\{zǱh�W��u�+uy��#0�$	��/+��r��-@�P�R<��Je�U�}N�24s���f��뫧��a���bޕی�ق<��~�A|�uǸ\�$�+g*w�α���,���⸣O���t���z�3#�7C��d커��u��"���:{rv��s�¾!���h���2�WC�E��vy�ݗ��� ax���.� ����sd㸻g�h��)!���0�$�����syK���VgCݦ֜�|��c���晥�x��	<��)7�^�^²�,�MM���}1�U�L�U����U~��˭�w؄��-]��:��Hya{X�nr��}2��o��H�fR�l�+uT��4f>$Ůn�[��>�-X|�����X�(L�޷��^g������8U;�ZM��58��e.�!�wM��hR6�̻圖`"б��+0�s�dk�R}��g���GC#Ǵ�-C�V������z9��N�r�j���}|�]ӹzk�T8zQ�����m�3\"��#���ǒo�n+�E��o�����3I8��{0.̻E�\:+Yy����効h��wx��9�Q��TNI��'�����{��N+�:cV�Z�Gz?q[�Un�g�{6ֆ�Z��O%�2�̱��nV���Y������g;`�׳��N|����<���]&:XC���G+\s5h����#e����!eS��;M�ͨ���K�T�s��뼛ƨ���f�OwK�S�" �������D��i��jI�ӳ��%L���-�U�.]�b=�M��}�'�a�|A]4]���3����M��D_L�_�B���.�//�b��.k}�?G�����93�i*F�����&�ߣ��#�oSĳC-ʼ4�cr>R�]�B�V�X<b��<8��.�7q�t�Q6k��+�c��P�\�#�OF)9�ޯj�䗕(���H[|B�H�"0�r;V�X:)�k�mv���{�}[�F{3ָ{�>���g�U��*�pIU�*�&[�^���,d��{Q\I
��5p�6�o����_O�wE]d�^�P\��㔖��0S=�kv�x!^D�-x�gZ��gm4.`�z���k�r@�X뭕8Չ��tv�7�M�\��;bz��]sѠ�OM�|�{�u�i��Q�B�����dl��w��t,����ݝ�~�j���q�Q����{%q��'L�~Z����Q�	�"N-��J��s���Y�n��L�x<�b{��o���2-E��N�b��:��#��{z�7���Ih�!��Y�����][��k2\������1y��7|��.�!�G��ӾĦg�'�珘�l�ֱˮ�J�PF'$Z�d�K��)C�5f��B%A����ka��ɑ��wG��i�`���;2S�,w�U����糌�:8y�A~�9�E��5����*}ʟ5o�7����ņ��m�s��ٷ��l�������6ؔwa����R �m��|��XQ�%6�ge\��o���H��L7=������;
���NW��qo�k:ucxuv�zǲ1n&Q�������:��oB)�5h�U�D���=�7�;����C�9�<�n8m���l�5��#&�D4r��TQ2���bu�	�rP�?Er�k�3!'<��5��;�.��ǳ��=z�hQQ�畖�+h��-�}�FEQx?\�F��[����F��n;0N�B*\�=���N]�!Ǹgi�@�;S��^�5$H�D����ϕJ���}Y}X�yzㄩ]oH���X�L^ýس��sG!����l���CU��m�r$�R
���I�17�^�?w��r�ɘ�����s�\ֺ�o�=9�=�Ť"�~����F��7�c���!�Sq�p�{�'7EQ���/F#�����1G���.|�޶]3��򨃝|�+���f�����%�������� exźL�W���ß�/g��Y�gEk�[�qҏV�ż}���J�j[�s1��@��lj�2&HU ��v�#�ik�tk�I��s���v$vۭ�`t�>��������p�y���v��J��N�G���g�u.��j���]슋Ӂ(Z��n�R\�#eTl�ݼn��]�0h�-�(�\΁m�v��Ʈ���8]۴Zv�7,m#�ܒ=�哳G.�.���q�T�$�\tx���:ݨ^e�����ч�n��xp[wjܽ�+�$P�v����7'��M��D�F�=k[!�LV��s���&HA�c��m~����+��y����8�b��ި����]���C�o�ܹ�-d�;v��w�@��v(����ؤ}��<u��{b7�r�W76VBh�C�Q���vx���=Vz+�~��(�w�d�+��nGӒ����7]����#:��mh���lG��ݗO9�V�ݝ�ķ7�[���>'�դ�9��Q�Xq�}iw@�jBI����~^�����e�'Zʝ��_�l�c��K]΅r�}1���ߪAb"mCUoS��,�g�G��Z&9)el���w;���Y��7�Ao���13@Y�{��yx�}	�wԱ�~��o��a,^�`
˵'6��̊�*j�
�A���R�8M�PU��n�b=E�]n�o�;�ǭ#bVp���\ɼY�K���(^���*���<{�g��O{�
�]}����70��Y��]{ު��6<��
�ȥo�ə/6��2���u�A�w�2�c[$���K�͈�m׭m����\��R�vP��]B��MZ�\���n�
ū-�r�K��1%V!~ܙ����x�a�opwHny�:<�ހ1����s3��m�B��D��Q�]C������7aWJ��5[f>�f_�����zO�u��W3�����^e�t��iQA����Ԓ���ӥ75��Kb�|j{3�3化����1	�"�J���6�
�IEQ߬[�s^u�빔ez���tQ����$��[�-�v.�ٖ�$ݜ��p̡�wxkߧ�5狕_����VdO�=34����/k�xF_��VWt�t��~��Bk�g�BlO&���	�V���ֲ%n\u�u���չ�F�]�������	]�/�O��~u��r�P�t^�b��8�آ�����0Б\�AN�+$镊V���q��6܋/A P��R���Lܣd�����L�qy��nO,N
8n�J��{�۷~����`�8<�Ր�����$�$����ʽ�n�f�0U���<������w%�(=���<�FA�#v�"��v�\�/q����.wtB�fV���m��]����e��A�&��s<�YZ!ݎ�oĶ-��L��΀��U�����۱�n�1���06B��"%H�����מ��o��vn�>��X�&��^�k��NTR�;��z���L�����|��˾[l=�E��!m��5�=&��3ν�R�V��Y���7L���Uu����~�ǆ5������X�F��\��s�{��Z�! HHZ�%a!
��&�!��`����Ļ��l�S��<�C��⁅92AV��p�ۮV�J��M�y��}f�f{3�6��ӊ����a����mtޢo����)����P&�0B�M��/D�몛��1�f��dM�����5}X�uU�,8��|�.�qk'�΄�=�t����O�$;dk�#fHTMHo2(�F+��7�`��Xd������r�]��&YG��������6@7�t�OXb�\wn��F-4Qo�(�q8���u�B�aU3.ۧ�Q����U�h)��OnF�z��|�;�(�^�	��Ŕ){I�8�[���n�8A�Ws�u�#�8�Q��}�q��]��8�6�@�/[����wx�ɩ:���M�V����m��K�Ǿcx�6�w�J��	����X���[}j��g����0c��V2�h�w��㶼�7���
^�n�2�]�iy�FH;�e^A5-'Y.-ܡn�X5WG3ǈ��y�^{�'c���\-�9T����]��8�1Z�x�M>#�(�-�wt�zK�ԅ�u`����|ޢ�[R���z�*Bʂ$�N�U�7�3i]K���.1��G�W�RS7�u�	��zm��;����U�y*k;E����1g>(��i¤V.��^9Vt�x��F�t�V+:���?	I��*w����_�N������&z�t�T�f��c�|�n'���+:�빌:���U"�}Oe����z�0rX�=��/;R����{T{.c�=Y��;�j�'&Uz�^*�(�Tu�YV���|wٞ�����<+��Z�eX8���z �8w��B�n�n�����ݪR�N��T�{-,�u�4�dWE�u�v���6��1�ܧ)���,9R�����.�����`˺j]uI��0��>���Ϣ�����T��,G��XLYt��+��[��%gd�ʺ�r]N)S���8�qk�vR;����f����ו�[�E��w���7y��cw�Ul� �M���K3n�̈́�<�OhY�+L�Y�Juj��A�rt����4�v�@�k0�&�,j\��ܭ�B~�l\Xw&m)�������`�}�R��g+�W��mⵕ�7t��^qfc�R�9,���΢�__�L�3����W>o��Oֻ��‬ԻkRȨ�Mݾ3�s2<�Ѐa��>!=�*߰���T��Ʈyd��4o�}�,Κ��c淽k0_P���b>��#=��I��]�lnl��u��$�N
}۽������c��W��*㡆�9��4�`��k4��d۱�;3X�����$�p;�S[�3����.���u?v�+�˱��/�+w��@��K�w������Nd�єS����r�bxnej�Ë(+(�����y�XX���y�/;�X�T^��{:�o%�c���&�+y��<c`�9��pw;ꭝR���n���K#q4ǧn�j~�h���=3�W3���Bcc��c�R��64�ס��ola3�*�`��tH�v��6�`4.wư��U��1�k�w���K4�vm�ʲ�o!��ݲ�sy�p!�o��xe���-��j�&l�M��bLA3�����*Ԓ0���k�sѝ�:O[�E�5�<�������������m3�Cv�֭���e�u�1ڑ�ù���Ȯ��Օ���e{cZ�<�:$�O��k�gXu�yN���Q�Ӳb�魝`f����nĈnG��,�Í���m�֋�xMnŧ�[;�Q�ݹ�\/YⷌR�v���ţ�՝ӥ���';���{6l�N0�7�����s�v�3�62�m�]��r�tk+�M�(��gγ�����v��n�l���S���q��T��7l.n�wN�c�K[�X�\M�v��nbm�E�vvpQ���]�yv�v93�9�����7#�r��`��f�z��X���v{�wF������n�;;lOp,���q�G-gX�V�s؞�r7'ZӺ�we�nci�̡�c�����;ﾗ���r]��g}��Ψ �o\^���ZۍC��n{]��� �S����VW��#]�5���{KX�۷mv8���B�=�����βp�t��&�A�70>��;�9w��'s���������>�綑:�u����j��!: R�y�*��	�G՞B�V%�8؞j�;R*��8���q��Ś�X)xɶ��歎M�8]lo��wܧ��{1��#��#G��c�N�gK���N�9�Yձۋ�l�V��gl�$�L:�*��N�Gl�'Lix�a��t	����]���ڵ'[��V���;۷���yͺ%�܆�k]���kPC��t;W��u�Β��;�'k��n�m���s�����:�ܝ5��Oj��絅�-�:�V\�ρ�h�z�p��w=t!�A�7�s�^�nC�n]��L�c]����vd����Q�%|�m�����n}c��NQ�kqة��˺I8{Fˇ���<r��r�'n���)��.�����0$g��۲�]�Ma��7@lvǶ�r����z�yz��i�/B���N�cl��yY�è{���d����4-�3��Z펆�H��{�
��F	�c�{gK��5�z���^]��v��fv�9�ɽvrv����F���gZ�y�Ɠ	VA�p�] �WN��cq�FN��p����ֻLu�6�nP���rv�{<��s�ƞ##ۮ�'��=f̙6�;�U�x�H㝸�^N�S�ixb�u�����x��\�l��3ɴ�9�6^�qp�gvi�]��ݽ��sN�X�{Q�c��f.Kn�n-�\'�8;Gcnz.sglu�/l�[�D��Lq�F6ԇ	�O�����琧�Uv`|���Y�mu�Zgӽ'��_��yK���z�=�@�C���j5!����ۡ����XuY��^ui���ه6����F�߯�Y�X�iu���dGi,~?`'}Y���c�_��Ɛ��Ru"�^c��Z�&�z��? Wv�t�~�T�䣦>\����7ⷂ�ԥ��3���~��|\�!'�8��/=j]��_Lt�d�^�m,?\L㻓�R�F�I�mw��GLF�W-���C$�u��bG\~��&�ZI��X14p���T���0E�Ϯ�x�^s�	'��9��35������;�ex�����R_q7ṽ�����(Fڮ����k�tU��u�n�M�ٷ=g\vNrx��f���yn�rR�RM�Y���5�n>̅������aͽe�uOz�1��Es����OYY/������t�o�R���*F����^f����J�k��s��¡�՗u[���dw[������g���3^����]�le�̘$JϚߍ'�~ѹ��gw�C�q��%�gt��\e�ʼ����Ctj����6./=�Ty̪��<�%��{6)�NɄ��0�	qH��,�o���0�\�&�7S��@�/�����Y�՝�-<�Y�.��e�d�-���7�@����[�K/EмS�N6�����ɍ�Zs�4\[����o��铋,;uGd^pu&�f<ʤD\,[� �g���	���*:��b����Ӓ�^Y���ɫxJ�_GOϹ�5i��f���3�\�3W�-2����>�qtOm}s���n���snn�L��e�{�s��`�<�MFO;��"�ַ0�:��]��w�ߵw_z`7Ż~��soܟ�x�>y�%ܲ�&�J��f?s��z�[R�Ƀ"�.24o2�2$,�K��WO^��rT�Z����:��y�S��:�T�.��\C꺞�ffٝ9�Y��^�E��oPT����9m��V�*�u�=t��}r�uO)��2�Q�)�_SW�"ʆ����9�WPj��D/���}���w�6V����Y����ʏvn��3n���Q�\�9V��"�-ܩ��!@F԰���y�ŵ������S���r�C��Պ2�mw�+jX�%���Iݯh��oU�>�"���k����ĕaX���K��O��*I�V�����Y�~g����M�9E���H�5]�@����&Oo\����1�/�]�yVs�}��`fG�*�G�gwB���������&��4��a'o�/7�m���{{G&u�� �����*�^�9�s��8��<Ӑ�c����ח�{3��ܺ+s�Sz�=g۩hC0l��2Iפ���uy\oܲkxg
�q$��XPDF8�ET�l����;~�l�(ۥ3�55��v��iw\	z�)���D�ٕ}LӶ�	d��
d�-��=M�*S�����X�b~ǘh���fh�n���{��>�=�-�l��g���ڍ�57a	��AHI�%#����[p�u����7ޭ�3�$�Ej�&��c+6�_>UX"
���
���,xT�_e��U� ۸Á�O2˥�(�V[���k~x!���wqS̬v)v��d�t��1u҆v%�� L�^j�Y�����A�B	lā�vƾ����O^��ʻ/�ą]�*�>d�nV�E8�PyJ�:���'��;��Mx�/4ەyY�����ϝ���z�<<n�q�m`.������� r����8Ǭ�;��-݇�ŕ�?����`{Ϟ�se���/l6��y;�f�٬/�3��vo/R�>;5��fy����������{�2;�g=����5(�7���}�zH�^�Ǫ;�T~��IY=��?��E�C0W������v�=���ek�Eƌd��f&��ɇ�Jv?��	���򱉝�=�]��%��PlA�P��p�M/2�{�^Io�<��)�&|��d�����/�+#o�]��َ�_t�vmy�X�ʆ�!��ʳ�˗����S�h�}^�͟_a�N�+*�Я����_Fq�Q��wW`5w�����o��km���R�e���r�o�H)��:�a��$�3���o�/��]�^'��n�sAOQ�br�`���eY�1F�_JA��Mb�]�x����Xs	����MNw�A�pu8��oy���"�؁���
O�o��ۤ������nme�.ۜ�z�a�P;�^�j#�[��+�����]�ק��	2FX�X��rZ���\v+#�3|=�s͉���˽�d9��ڝ�y�W���n6݌sā��滗�c$�܀�X��ݏL�ؙ-�̰�7k�:��3��=��q�ڼ�c��筷0�nw9��Ƿ'<5����c����s��v��t����׎u^�^�'G:�i�'�����]r�5�`�����[/������]�d;��1J���y��4��ʕ�f�׎��YaV�-����_������%5�h]��o"]v�ge(i�S��L�]�3�gR���zQ�\�6�h�u2�=�p�'8`��Tg{vT���Y���*��9��CW�lv��c,��^)^R.ݤ��\wms�y�Vx#r�Q�ڐ�9C��Ǔ�^��Sh<�/.��WHk�Ux]8�ߣ���dg���h��M1�~����^Y�N,��8�.A��ïN�v�9T���|b���]��V<�nt�rH.�OV���}oT�}c/�D�����t����&���ݎ����{7<�v3tY�K�wl��T�ɸn�L�9:�}���8to��m�{o�{�odU�43sv�C�q�?wzV��L=�+��b�*U7c�_+�=(�|:����Xr �r7W���������[j;�z�!�d��hp�]��)��m&n��pc��4	70M�}���-j\{�(,�(��ڱ�s�8}Uv)�X�f�u���ޮ�����Ɏ�(�s�w��mJ7q�	���=��]�ħ��nn��9�y���~a��08CP�'x�'��g�gf<��U���꼄�w�����P��UU��I�lc�UG�s�-�3�Hm�&D�Q0����U��;nw�Xd-���$~��IC��Y�GiV,��a�[��� 4t���NC��j���X�IO7�;9��_��-�r�V[}��v�Ʋu'E�ʪ�ʒ�%Zy/�\u~��e{�k��C{R��g��=��rgV�LY���M��hB��O��7n�͛��:�����qU�	e(�øD�Aey>ʂ{����j��^��A����t֋=ޅ�^� �*���3r."]�޿�4<�F��.B�q��P�wz�K!۝����Y�\e�n�i��ڭ�8x�����+��}��o�~r����jl{����<$���0��B0Dr38ZfGC��:w��O\��ÞQXbF�'<��jƷge���D��(� H��"�=FQ�u�bs��b��l�tm� �\���4�x�\�������{z���31ܻ��y��=��X�!q���F�.Ż\�/�Nl�i]�U����rٹi߻C�����p���:�_/B�"���[A��B��~�������x5r"B�Bm�B����w1�roӤ�x�vt��%�=^E�9rǤ�k1}d�:
�d�`���4z�&�$!嘣n���Lo���}�j�+3 � z.��ĵŵs实�ݻy4Ӯy:y�]�p=���
���H3$F6ܝ�n���}�S�EH�H��Qn������w��%�ou��ǈ�;R�@ޛ�� ���׍0��l-eV4���vL8�a�8z�Z]U�^o�^�����L��xwUL�|�qd똓l�X��S��xÎ2)���x�jr���
�F!jI�ܽ)�	���Y���J��o�ZT�U�J�w�u�.ov�T������V�n)�u#*}f8�rA6�3oV�]�X��w}�Ƕm�Ǉ����ݕ���L{k���3l�@�C���O���0d��Y��Vf�.�"J�JH�:m9W|�m���Ռ{�Z���R� ��(ʷK��Q9��]��w��ex�*Ρ�_u���v���6P,D�e"�b��v.�ҐK��Drn�aN=@�q^�5']�k��-���d��9�6�k�Q�$�_�m�)D�!�8-�v蝹�:;�Q0J;����I�/�ŷ۴�����#&7 ��Һ��u�NrO�������,]exz{�7'<�w{+�m	9���/���Ӹ{���H�E��-�y���������fy�Q�ʘ�c<��=��if����J��t��Ny}��N�]f�C�_�{D�`qHC���&����;�zЋ+]�PI���>���iHKw$����.�-�g��x;[$��ܯ�\���P O���2E�v�*�OG���;���Ӻnj�^C��]Z�,���M��ں���	)�rq�xȢ/*�{r
���o8a5�����(�IV�9<d�C�R/z���Ծ}V���V�$��O<�<L^/6�yK��G�g�gI�Hf׀�x��d�3w٫����3Bc�Ac�W`�ڵ����?��i�6�#�7<���bf~ڞ�A�;�g՞�/S|�5�i���Yb4V-ܪl_'�ޫ&6��>}]��7Viq�>73ͭ��AϨ�u�Y0��}��H�p\g�6ܸyy��_�����y&�.�d�Im�μ��mq�]��ѻ�Rx}5����9�>�Q�6�cu��6�6�6�qv���k�h�㍃��=Om��ł�v���v��k���=��fw�u�X�{m)����Ns�y�����y�s�� 6�^��ֻG8l�h���\���R��M� WI�u�r���s�J�֒҇7�bC)�K���l�������^J�a�:���X��?��Y��\ӽ�5^[|e{@�$�!� ��E\�׌�N�ZX�X_��Xtp*-�uח6Y�e)E���=�jIw��;�;�*&b��a�B��{�H&�R�F�X^��"����6�'�^�|�g��ݱ�|����ْjɡ��)��Ux>�~�9>|�f�B��BT������[��5�!+�쬑f��n�û4�����OMv/z''����(�t�
�y�v)^���:���G��Nd��-W=\:�٥�\�ne![�gjj�&fG�͗��㕹~�\�^.Ϩ�]ʦY�U]���w��l<�{e�L�HMd�k�WM�;�ms������Ѝ[��L(䘎'�mK�@��D؀���s�ɞ�S�O)��=t�M�ˣ�x��A�9������nV�׉�U�U�Z��QH�H�QFI��[u��of����[���'�%,�9�V=c]AS�&(���\ /s53Dٚ,��c4<���i�KZ?v�����N3�m������O>幒��X�����e�4�D'+����g��ڪ��'{0�쳊���
�io���S!�����^�ޣ��1�P���I�~Y�F��ݯL��E�V�\�����VdTj`�[���	�:���
�`!\m�`a��%� øՊ��5P�t����=�����{=m�zE3/�ݪ��Okv�����^Q��P��S��ꭐR��M�Q�R�sM�-�-��w�$kj�^ƼSG<�2f��_����%�ڰR�ooױ� yB���hU�e֕�*Ǹ$���|�מ�պ��F�����5;�q&I=e)�����v�o�7�х���mO��p����V��TnY���;�2դ�E��].�Oq��]���䀤��j�y{��}W���+�4^��$I	�Ȥe!�0C~=��b���z߶J�<�_���ʝ�n�-�:�3E�SW��;ޚO/{�H����n��jGR:Gf"�A��'�Ъ�|lA$III�B�:u�4�B��ޔ��0S%�X���\��l8~�}�Q9"$�ۜ�oR!;�x]���	�Ⱥ��N��Vù�εO�3�oQ`d԰���� �L�	�N��f1�\��NXY�4��w4��8�5ܺ�y3Unr�t�v:�g4�s@���	��_�l��݁VP�)|w�m]l��dֳ�����l��L�e��f�N{1��7��2��Y��Q��9�b��4:��w!V1�1
xX���/%V� xVX����J�^m1�Kw��ҧ�*�c��fZW<��w%�8�PU��
;�/�켚n��N�K���:�OU��{wy�+�`0U�sf+����W�F��%:J�r��r���2����4U�(x<�����	 Ѽn^�Id���j3+M�:��;�оcc%�Nwl�BP9����ݮ۳�
={Ih��.b��
]�1�M�_j��[��٫��mf_$[칽\��Y�9G�Ko G*/�Q�ŹPU�^�2��5Y�����b-�ѡ�u[�{�yK覹Y��i��d��x6<��A�]{���g���O.�t��ot��f�\"}���_CZQd'\-��Ò֙8��W6��㽵�.*݋��3T�X1�]�E����5j�_�ăߡ}���%����=X��\�{�M�)�#n�����)w���Tr[�w�ُ�ǚ�1OU���j0{�5�1mdY~ю$�+��ƁWH�n�;��.��R-�Xr�1�mZ9��Fa��sWkYn��|��":�����ԑ�*���Q�9mP�st^]C�����8l�躼*��C�L�VI�����]qu�iG�����ɷ�QhT7��a�F�G���ϖ��)c�5�bȢN5���Y�t~��Z�U;����r���������w�ޣ�u,`��-�ya���b�ț,#$��b�;#m��g1�o�tU��(�u���Q�ݕ3�U��������L���J���b�?=�����?B�0w��X�������kob�؜JP��"t�+@���9�k��nm���ֽJ��E76�F���"x�����aj��)��C�<I�}R�8Yn�͞υ5���4w.�*��w.�o~�|z�p���*��`Л*��6��˓����#�YX[V��Hω�K�E���b�T�}�}��ɗ�A+U��u1 �;���;�;&�^}NF�Pw܅{��O<��t��7��.�]�	r���p��!d	�b�ŭ���(�XB��7��_u�}�@���N,�ܯzg{%s?o ����pi�'�l�d�����TB���UE*�B$�K��N�6�L��^��O߮��N�P�4��(�ݽfƜ#�O�Si��(��/�Jr�3�z���4a$O �M GBȳ�_�?Ks����!��h���*�����*�c����@ۇ3`�뢂y{�+�2ŅO�{^�EI��z8jmX�Z��q�[��i8mN����jp.]�{�n��ߗ�*���ܭ[|�G�r�r�tϻ�6͊�~����Q�yM]��Ìx��[i���T��j�w��iY���~�|UW���s�{��:W�*�m�:�;��ɿ6ffH�?�!�g�_�'��YD��D#���K3�7߯��^M����w��/����ҳZ���?�Q�=T�'����.���ьx�8���?3g���f'nG#DL�/ԭ��yS�;�dګ�מ4�V���cpi�pW��2��0��wU��7��a�
]�+��U��W�k~��}T��ˡ�q�V�A���1��{�h��Q>�M�j�_ߪ�iJ�aY��έ��h;;���g���b��U�w�KJWݫ��S�o�٭��N���c�A4�6���ܡ^_����}$P����m���:�ƚ��m��jD�a���w3�$��N+>��˅y�G9�����_��~�<~�z�衘��S�F.5�hZ�߹���j�@�a�ݤ>,�?^��Ǧ�	��#��/ɜ�P=�� ����h*4��"��!!-w��vS>[{���H�I��?Dh��~d������!��\�����ӧ�~縛9�-l��?w�K}�U����&�J "yej�I��\4mG�)�S��ѷ�X�诪�y{pC���eh�}�_��E:Q���V�zci�m�ο+mv߉*��~:��1 ����K_�W�v�?b�����g���Ό�?T��;�6���/㟽�p~��*h�X��У���w߿}�ڨ�^'�>��a��W�I���_���F�~I����]�_k�����D��R�~��.��*$�	�`RIΡƓ9��v�M�ݺCv�����Ϙ��%�U*�~��2~Oݮ�G�5�}�7��|�������V����V觉S*�wQu����6q_Q^O&:}U6�_U9F������5����)���Z�S���^���pҞyeu~ܱ��M��	z"2PO1ূ�4�5]JU���%�Kwe�ծx/�m�WdW��Y5`�p��D�M�ZA�?B�ɷZ�8qv7GY�=X�5��u��i�8N3/R�9��嫭%ا��Ѹ�<y�n�a�"������=W;�j��������G�q�}�r�z�q�RuM����,u�v��:�2��j��{�i��+�;]���v�L-���n�=q�q�ӆ���j��ܛ�s{�ɫ;�lq����&9�5�7Z�e�I9^���v��e�y�nic����`�Q�2k��<��L)�E�@�婶�;X�v���Z�f���G���+O6�q��Ri)��?�����S1����	�-��㋢�y��y�a��݈�eJVҵJc������E���]����|�] �v0�#֝����"�xݤA$�����,�PF��8��I��'��ױ󟄗袶�t36m8�������.�>�ӎ�*���f��i��}߯��$R^�p�E�qE[�w�nm]��Ƙ�Њ�{��t'��⣕J����~�!���n��oP�k��#�Z�~?����{~HY�p؉���4o�7" ь�]��:�w_Y��I�U���4��}���S�T��)�ڼTG�Ѷk7�Y�a���"]{����4O#�'�����~͛L�3�J�t����[a���|�	L/+�^n��Uʷ���|~�z��AH1�f�>��������{Ӻ�љ�D"7���V���=Mg�ٴr�C��Y���:�o������q'�Hxߕ-�8��~@]��7џQ]�X�tT�z�T��_�s������»O(��څqT��_ I=O�"����"�ȍ���O�JF"�(\��u<�8�4�Wu_TGtW�w��OO[���GH���vv1�� �}����p��meء���B���?�9=i�ͳ�����	����n�G��UIꯞ%������S��ƕRK^����AQ l��އ~��Ô�j˺q. �d,u��#r"��L%7+qȼ��i�;x��W�۷dݟ Z�;�nv��8�^W�C�j��v�̮����M2�k�?s��^=hq�]Ԩ���U��|���4~�ϳJ�����2�����v�ۯʬ�W��.�|~&��Hj0�X��	�W���ַ����k�D6Eo�3����x��o*�l°n�ϟ/h]s�y/�
�}hO�\a�u.� �����C쉙V��ZGf*؅��-d�/��B���2�.��M3ׯ{1�u��bՔJ�դ�Y;N�qy�f���9}�?�ڕ\����˫}�F�W���~�]'����q7�-C3��V��}��k_���Ҕ��r���k�y��?aA�����S����?���(NC ;�>��2DÌFN}B�JT�Pm�T+*�?��U��AoQ�tЇ�z��F"r����kE��\q��ȼ�z5ɉ����I	��/�׽�(y1�QLu����m�6e���n�U:����!��i�Ѵ�i�m�];yQ�"q��q�c�IB=�Y�@�k��]Qw��!���ڵw�B���ɶmL������2���Q�r�6��ᨑ��?�B	��f�x~����/��% ����ޚ�W��7˻�I3���[U��ҫ,�]�=uU�z����8`�a����]�raI��ө��~{�ߵ~7v��yE3]�2i�E�o��Y~�<W��<Ew_4@�򵆉L�h�?~������2�����E��|��R_�������U��Ys�Q�4�|������mO�˛��ꖖ��(��!K<j��V���i8zp�Ƽ>V�N鵺=s�y�`Ս�f~DW�<�8��R;�v�iJ�+_�z��[N���V��m)R�����s_�_'�]*���C�<h����۾VCgǣ?�b���AW��Ҙ锛�ʎ�z�h�8�"�������{P���?�?��2��5'�4��_��A<@ۧ^o���~~��N������U���u�V�#��G��{�_�)^�.�\��V���-�%���-����S�h��Q�������Z�q�)FEB��/a3q�4���U_��!U�ĄL��)}̼]�(�֏�\�e7U*"	M���X!��u�5����b���U��
?C�/����BŇԅ��m���"uh2�m�>��`�)��d�����/�#�<��	��K�����)\!�g�,��ً|w�c���/o����F�k�D��@e����؀4���������_S�L�VQ�֙|(ۦ/?_-�&"n�%w�+��kM.���ر���&/�'r����yo~ xοn��x�!D����s��j���&B���U����>f�<z�M�m��s�&~���_�'mq�D�u����;[閖Y�ޮ�b5��?Y;�]őE�NN'��Z���[�7�S����s\�CHX����kL��j��iiꦵr��~�/���ϽU��]�<F��,�0�!9�
�~��q�mǭ��F�v��=|f�\���(���Lq�t��{N��&�S��g±1Z��%��|�읋ngu7F���SÁ�\q�;����Un4I��n�H����5�We �V�T���@U�#�q���͖��I�߮W¦~0��$�<�ҍ���s���r�;�>��3�߬�_q�) �\��~�w�b�����ߜ��!�D,P�0�#��?��L�ȍ�������o*&����6@�7��%i����h�r��a���	?Qֿ~L��]����"}�����~>0�H�G�WIDzf[��*�r�;�_�C_;4�<�����W�k��u:�Oki�}���3���T-��w�0�"H�q��p�������oڨg�aǇw��7�'��1�<��� B1�>�`�X ���H���{��B9�F�dx�q=���_�v�?������'Q}������u���7��3����_L�:<�$��#�ݐ<�QBc)1w����n��e��ߵ��:�r����n�b��%j���ܳ&��3L1wAo��A�j��-6��k�a��tL�t��D�Q(/�£A�u����nB�pSR�"m7I�,ʲ)�B���1��Ujڣ9����x���6��$�u��ѝ�]yw���DB4�W���06�8��4�����Կ#��㤭�=�Q��ͩV�F��_�A�����d��ө��A���w�k�����9�)ףl�}�:�G�u����7T��f0����N4��P�T�4S)=�񉷭O3W�����i�@(0q�h�!\tF�	:��U貽W���;�]�y;axq����2�
���~O?��16��\��S�rY��_óέm N#s"*a������Z@ܭ�����-7�����g��k���^"�w���߿T�|�v��8�u����e��
���t���V?���	�DIIb�`�[�-��[�[i��4���~u�Q���^����p�|�������]�Pv���U����+��	���	�{���i�B��Z��/�~��*�>̺��|��w����Ea�>q1S��l��uw�+�54�=�4�Y����ŝ&~�+�ځM�:La�V�}F���:���&<��i��0p�C�'�C*G��f��4��&��ٛg�VϽ[e'��4w�<�8�e�3�ь������M��V]e5Eӄe��3PgٌD�i?˻.4�z�bm��=������l:��{ws>˅�����j��u�g�"�r�+M�zg�_�j�!����QG���O߁ۥ��֯��_{H���CŐ;q�(��� #����㍘�j8�I"0��@��v�����S��j�:�n�'���~�n눢C��xE��d�_V�?B4��v�wk�?~�������C3��o�5�|��|[�N��U�|4I�h�@���3��'V4���`r���mC�Q8��]c�����+U]K��A��ܞj�:� �bX\^1&���
s�`��,=�ڷ\&ɵ��e���sN�x�;��ۜύ�n�I�g���4k�n�#�w&\�.��s�Ĳ�A96-�9��cdq��n"^ֶ��V{c�	=���m��u�0�Gs�.�+�H��>a'�t�݁խ��X�E��&�u=b��hް��.��t�#����sۥi�{e��v�Ov�3���������vB���{[���v�d�7 �ʦ�Ωׂ�qٓ&��jׇdn}��N뎸�:sS�nK�.���Z&TR��r�2�OQ^���Q�x�������m�ߪ�L4�e��ɻ���h�|�),q�7�+*,/�����ƻ�b~���߾�y-����o���Xs7Ͼ��gYO^ޯS����5A���gA���T7yW�n���=����f'��~��xאiS����w����}��D	��m�/ެ�k�
f��Z�=��褪���+���R�������BZ��!ڗ�|"*���4��9�#O��><�.}M30���js�m�����u����6S7���Kf���������~��9Ts�>Nv������w]��w�Z��ǽk�^t�;M&���W�P�پ���G�.�e?��R0����ˡ�"m� iĤR+��ۅ
(����v%���?zt���u��~���y9ʛa�k�b~g��[4~b{��&�G+�4�w��(3���2/�����do�������`/�N����ݢ�����?*P�����7�f�n�*��*�ʬ��������;j��4����5r��m��B�^�E�g7����b<����_m�c+�Ry�����4�X[��xgޫz�7��Z<�=B�骝L�O?���)���~��ݛ��ٯ�)ݕG��VE�h�fq�y���g�OB\���v0NwS�q�r-�::�!G�?o���1�x��r�)u��_�ez��돫VR|�)-���;�)%�_���4x���{ߍ[T�/�O#2[�u��^�5�V��n�{��)U�k�)~�|ʟ&إ�O�g���6-�b��a�u�Kk��i�)�F�l�V@�'����q:�=JB6.�2�y�K�j�~m���kj�)��7v٨u�T�^#:ʦ�ᕥV9|���Ub�1Q�a�{��v#}@���y]_���S3۹�i8�;W���}�����6�{�l�i�/w����[�:��A�,���`�)6���!�j�[�9־��"V"ŝ#���
�?-h.���i�.97����äC�V���ex�o���*�~�&���m]|/�1�?���hY�����������~��u�O�z��K�ր����]M'Xc����VZ_�}�э���[��L�/�6Zi����j�ٙ�����E9�g���H*@i�Y����\��3�E4��U鏽¾?~#�GSi�>��ᠷ1�s!�>��[��`~���?x�i!��01װ���v��t��w�P���`�إ��k���k+�����F��+3>B�anr��g�5��;V�m-7��4�s�~{��+���u�("'*y�}dw��:G��_gJ�VG�����-|0��s{��yS��i���*�`�N���_|�R�=S�Ϣ�lW%��5�2�����'c�Ȇ^�x�+�,���W�sq�������{tw�a�}�ٮ�b򏙦�g�o���|��(�����f5���f�ԜӾ�<��wU!�Ոh�m(g9z٬v��l���\�c�yF!������I��*���̭y���{U
��YE���O*�ec���:d�ߑ��ny��#?w����������L1>gկ�5�'��i�Lv�����u<h�y�/P�M�l���O��F�ƒe2RRF������͐Hk�ٳG��f�M0����I������������ó���e׆����G_^��o��s��wP�^�|�����M����7-J]��437-��d��{F�h�Q��{չ���=�4R�x��G��8��{<ý�?s6S���ha�V�i�:�64���ә�6Yn
����N+�𣽞u~�s���g�z�g��E��
��C[�q���g�X�_Y'P��Z�B�����6�6@�Gҝ4F���p�>���>q�7�͚1��P���q��a��>��m����������q[an;f'�����q]�>ʅ����Ӵ��EZ�Ҳ���3��WY�wTm�<g�S��ۢ��\~��@����{�X�9t����2?F�AG��,2O��Cm
;�����l��!r���n��y���v�B��ݶ^�'$��-�EXTZ�
�[_��}�PW�:�8�מ�~c��g��-���w%����_u6��n)�w�cl�=��[�~�������x�?qؾ�D8�k^�hSN��8��f�g�cuNĭ�jF�
!I�-�?@#��;��$a�+W�j�F��՟�~H���ek��;��Z~�N���i�v�SoS��[���8��?w4��:��N>v�g�l3��f��T9���/�Us�l���nڗ�p��m������&0��u1�~�/�����]�eq�M?Y�H�Q���|+����|��,^T6�W��z--۱�z��C��4�g+:)�C�<o�!�Q�)���Ó�"\�B���|0��#�o}�����6D#H�oݷʃ,��,����0�}��G�\���5SO�al����E���G��0���{w����n��hg�}�ɗ��ͺۛ�[�y֔��y�8㹓l�H��Kt������u57�aq�o��#d����p�?k�x��͢sC	B���\����]8��˪�1);T��V���CT.0���ZV��z�7��|��}ҁ0�?{x�?eT�@// Q����r���٠�ǩ������/�:������/�+��Q����L*0�on��6����r��+��xw�nܦYH�i�!�RR[N|��}�
��c�*߻.�F��f��@�C֮�P}�?Q^!F��@��㽢����#ꮓ��O׈^�bh�.os���=������C6h�A����m��,2ZE9�Ǭ-����&'7���>񭳯�ߵ��������ͯ�!R��+|0��.�Sk/ɏ���z�S�Ѥ��Q�fg^X����4���8�xЕ�ζOo]�YF&6�E�%W�.��q����'���1�������u9�Y�i>e��s[��r�����K��j��s�P׍�(�@m 2+=��~̯�h>z®�3O�0�}��j���ԑ���١
*�`o��zGd՞ȣ����!el�dix�����j�������q���h�8��3� �iڽ�������]Uo�3ϝ��3}h��W���]10�ʎ-e��C͹u�i�V�L>�_sP�v�[�J�q�{�bz�2���ʆ�R�b[{�`.�D�P/Y�w0�^���U�XRJ�c&��3U� BO��!$�r ��� �T !	'��!$�� �$�� BI��I?� BI�p �$�� ��� !$� ���I6@�P �$�� !	'� BI��B i$�$���I?� !	%����d�Me����~�Ad����v@�����!|t8@        
     �   �                      @   �0�Y1z��Ng;IVl�T�n���m����ݺT�dP�7A�wuQu���m�����        `    �@�:�`Iv h�� =�r  ��9 �{� x4 p     9�P;��� h@ �ݽ�28i]�@;�r;7m.��4u��-t��j�eu�m  �AM�J�:��ri�!K���-n�$��V�fQjA7nkI�;�  n     �[9�W7N�sw��K6��i��Yٕ���j�iH�1
`�$���  R�s��J�:�dgf��ۧgwTꫀ6U.�ڕ#-K�����v�      wjW{:��{�i��UN��� l'Wn��m�&sV�[1�]��Ӫ�ݗ@ ��Wu�� �Tfӣ.]t�3QL�*,��l`;�ȥ�]�9�j  8     .�Z���]�:m:�A;��S�-N��.�sa#m@Z�N� Z�7s�K��  ����ru�N��+�QKv���X��9��@ H}TT"")�BmU�       �~BR����2h 41 2 MT��4�m	�L���4�G����UH$��h      �~�ЙU%F� ɀ��I�D�I%<�I�)��4h�0�����~���?���?�2�|�}���I1�B�������s�S��Bγ���! @�V���F��I	 @�	$	!?x��|�"��,e�~�?�4�2

Ed�	H��$�
 �Ԥ��@��x�'��7�Y��j�!@��?���O�������C��)���/R!�?�΋N����U}Cf�}���6��u�m�2H�	��ٹ���+�̷kP��z�9J�0^3���YƎ\.bͬ����)j<�@^�;��i�okTA֛,Jƪ�-�>�Éؽ�t+kL#g\�JA����Щ����fˡV�]��b���9�F�=���l�`����.^�B�w{M\�g����l��a
�rN�Ep�CVy#�4����»:�M�{���;u:�|؆V�[�lC]��A�k4�]����/-�N���,t@�k�P�4�����2�X�n�F�5���\2�|�v-۷�d�w��mk����3v�+�����H�y��5���?Mķ^u#���η;z�4J#�wI�\*}{k,�N+��8.X����gRJR���.��{ٝ��C��3��]��V~���4�<URJj���^v9����~2�
��&�i�\�5�wIU�$�u�V���ܛ��s��9m�NWSk��Mk5HU��W23�W:9�oGÊ�R���S"�*��,�g�f���qn��)���4Q�>*��H%��~7�����ؤ��Q�:C��oqku�qpg"���u+,Ps�R�2���kE9*4�ut�ʻ��������kE[��v�V5������w̃NKZ��t�n�TJk˪�6�Х�^Df�h[ c���L��)Z�ݼ.]�8�ӻz��*4���j�az��D�M��@-��wh�0&��ăt�Z�ŭ�a�3%�֚�>ͬ܂�^�g�o(]j"�M3ỻt�,R�+���1;���/Z�����I=ڽ���a�$��%M�T�]M�%LD*Y��2L�)�o�Y˵E�[W�fQ0�u�0Y�9/C�r��v|�E;��j=[)Yn�h��f�eeY�TQe3ώ�H�V:�ZZ��IY0f�6A�Ta��Y�����D��I4���[WX�ѐ��q�9�ӻWJVe:�il���ӈ��q���+�B�so!Ku�7��K�kJ�
����x7Uܬ�7�t�l^uUxa����`�e��ɣ5�Z���#&�:h�{t^Bev� D��� kk-�݆d[�2����P��N����� �����&Z�;����`��
ۺGli�%N�Mj��j��
0
6ZD�A��ђ�uu�n�h{*&�v�bƩ,l��q��&�>6�v�`�����݊��e�i���$u��ا	^K��U��q��+2�E��x[{E$&]�E
��f�m:'fm�n�96^V����T��ޘ6�3�I��P���O*m�9Jc�kh����\�f��b�n�����Z�w%�a�pU�j�p�E[�OXūH�u>�
��[N��W ��n�6��|%��5�Xd����Z/eM CA%N��&�E|��M�Y���j
���@���.�^|Љ�lCK\x�'Je��k�Em:�%�#��[�4E���=8�;t�5�%�^��/�(�$V��q`;��v�2���q���+�sP��m�����[$������J�Ч"�:�6��vL�(̆�ʹZ���y,(�������5��u�j#{�em�b"nˢ��su�usv^�t��\���E,BS����ja̗�z��"۸Fcg
hf��N��兠ޚ�0d�ř�Un�i����Y���
�^{��Ƃ��ΣY�դɛviVޤ�����1X��ň\�5��aj�T͛���`ɵ�[��%a�nB6�"]�Ct�\�PF�e,�E�J�i�c�d ��U36���Ay�{fn]4��[(��Mj�e��s5������ ��y{q��k.ȩXN�/.i�{��//n±��[F�l�W�n�$��+߲�^
R����o���[�%K��\=F�`��w�b4����i�W�U��opVH�_ly�N$6�|�860>�Hl�M_�-��nZ�����`�ѫ��<�����9:W�$R��1�����y[�M����h�q���XiWG�k^7yni�n���Z���m�H�:]���WV�'��KY��!�PܨM�G]����o 5��ɕ�E��ک��Ӻ�e�P��'p��ߞ▧�O��V�H�pe���Y��E�����ۨ���X��{%�ڏh�3{Wp���J��=ɕ6��s�snB-�vn�T�ы]jnGʮ��"����P�Id|�M�kMM�1U¯^���ݩi�jҸ&���T�tι�j��]��UX]Tm`CnV�,X	F��i_�Q�[)�Mn��8½�3k�-�wFX|�����v1X��׮�M��2�zWp�t#0[�,�M;�]�c	���حWS,m] �8�K�Y�����ܷ�$m���y_ٔH�[��՜ٳb
b�i-F�I�wsӪ���]Hwse	F�R�0K�r�����Va3��L*x�:,2IW�v�"�6�ĳV�Q�2���B�u�{�hŐ�nl{u-�"�4��v��7��I�/q3�2n���n���BP�WȌw�X�n��Ɇ�^At˔]	y�|MOpO(e�X�]".�|&`���bK>������*��Y��^��B�;����sHBf�*ն�tu�록�G��pwR�%l�v5&�.�\���y!ǫ*�[���Y�u���B���R7�oiͺ�4M���l�mGV���$C��L���dtEG������yIZ���2�]K-b����^�wr�=�-��-��m�컬x�e+t�r��Z��e@(�x+D�Z�2�7!���XV3Mఞ(��X���4]Xh��df�n���8jV�%ܨp�������ǹ�kQE���nI�/oYp��)�2� ҫϡ�g
y��b�;�wQ�����л|��g�E����D�t�;��5��M�� �L��)���^��-[hʻ�"�R`�;��n:WB��ʽ�5y�k�y����B�e�Bb��Y0fX��(��ֽ�X�B��^��3	�j��F�4��n����B�3��c3V�VS�&^��6�:!|�IR:1�J��q��ո:x0�w5F�]�V+�n�����+h*�X�Nـ<[Ndn��̽��.�.�жY��U��QQ��Ա��O.���^��Yԫў����jҝX}��1�pSk,՘�S'P�Qv�M-���t��kj;�C��K5��V�K6�5��/;pWb�@>�9�"j��;{���9s���P���]������ T��;Z�Y�ח����@*�t^N��s`��v�.U�����YITW��!�WvY7���e�Le;��襈[�pZ�KR�Xw�z���[��y�6Ƒ�\�Rsw�n��"���ЖC�*������c�.ՂݖZ�ش$� �P8��u�C1�4ԥ3ʖ^�K�jU�����.���
��m;ӌA�t�i�se��eo}���fw|e3�sKd�P�����̂[�ea�޻��2G$�ξ���nh�t����]_pU�BF��: ���F�[1�t��w���Ė�F�< ��e�AcVI!�ڣ��6�|{;m仺9P޻�ZCz�a�Y@3���ݨ8���=��T���p��]V�<���+@������Ks��)�/�w�5��l즞u��%1;�{ESj˳�uq�i�{dP�k%B��:���N��K+�Q�ޝ;�7O�ŝ�3��Cr���I���A�諭�o��}��$D�Yd��2� ���J�����_��F�A@BE�e��t�@*�US��0 W*�T�����т�]�J��!oPeLe����U�tlQu1�R��1�uCu��q�w\F���gEYNz�U[�J�QU@UUmm+��UU�h�y��'��Uc��v�������������������������������������������������������������������������������������������������������U�SUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUz��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUN^�ՋHs�jC��!6��7����WP��<��j����-n&�w8���56�jk��K�U������C��P�֩�=��F��i0���p�ܮ8���J�����5�Gh�kqf�ԩ��Շxyw6�*q�[��.5��n2�ay:�YMYWN�0�v������u
�|��n�u��0gQ��m�{U�n�͑�b�B���r�Lׂ�nsv�>�!d��e֫]�we$˴�K�c��d��6��F�܊*Av��w9�b�����X� KDm�h��I��{i�0/��5v�ms{qƹ0��7Xp�ݙz2nv�md�^�'�[��ɻ�����ۭ��m�*c�g�Y,ʞ{�=c�C]�[%�9�a��/>����z=c�5�����cu�&yp�ͺ5vm��=T+�{< S��>��*�`X\���<�����M�t-Iƣ��q��lF�aeɲ�B��e��d��Ot��<b�w`�x9��Glnmn����w1�"]Ν�����r�sg�����o-�j[f����x�o\����������!�ݓ�NNS��67w[�λX�#�A�2���n-�1���ۡ[��NxGJs���:Oƽ`m���rƪ1���b�:�W�ݞˍ�1���P�cû��-��9f���ힲ��7�d(�۲��J��gqDj�-ې;��8�k��m���[���n�{Gi]�.����u�1�z��G$v��1O���5�0�4rݻK�l�n8�7l3��^�r�.7�7=�:��k��P��i[k��f{wG��\n]/�����}m���[�v�\�b�۰��K����wk�ۄ��$�6��fz����o'#q�f5��:,\I�8��[�]KT��������e���AyL�M��d��Q��`l�c�D�lx���o6]�W�w�{���jw��(q�4u�s���IG�����W#��l]u���r�M�p���Μ'3���p�d:ȉq���v9x?�~d����]��d�k��8�˵��oW5մ�m5�v�9�g��{ndױT�K���;5�;s c����,tՄt�R���(Zpթ܊�KK۷a�KY��׵�c[<sM�;u=v��Ip�:��X�lN�/��q��V��5��U�:�ɼd^����k����q�� v��q��6S��N��Wj.�v<�l�������u۶���CŻ=��œy�2]����c���l\Z�7pFXg]�Ź���%��9y�����e`��;�K��n{r�\x��c��`�ܨ9�kF�mcg��sf�˸9n4�`��÷t��;�>5���g�;S��EU�(%�mn�s6����=rs[u�I,������/|<�nS�ob�{r���;�K�nhr�װ��@x�7j����8��f�#�ݳ�g<��;��_�_36�cl`�s��px��q�.��� ֻv�(�q�p��b��<r<��Gl�����#q�1m�S.���8����A�i5#��\��kf|<���6n���,��2��u�{=����<>��\�^��};s�wnې��s���ѻ��|zu�b�݋����&���8QՐ�����m�Z��s��|��ήKg�	v��ݵۇ��u��X;sc���8y����Z���n���zv�v.����p��g3�vG�����:�(�
��9��P'��7g�2���d;����4���gf.�l���nt����q���i�cɸ�Z�xF��xk��3^,)����:�!1X���/g��B3.���&��l�x6�uړ�	:=��(5b��zm��v�s�ۯ^��#�q3M��rv=�U����ͻi�Eׇ��{<��G[��j�v���-k�����'78x�����q�khGs��+�rQhc�����<vG�ruƸ�\�to^�F��VD�;6z�l*r�G1��]#��jj��ɸ�U1֗��i_Sp�A�p�fy۵�6$ݚ.w$��gۃJ��v�~���ñ�d�J�M��2Mm�v����ٝ�����2ې��eTCk��`zmvbG �ӍV��^�ǃ<�z����܎�뱨�n�6�)±�Wmp=������E:�&ʂls��ƌ8j5�cTn=�w;�e������z�M��:.޷f�ב6�=�V.��v��`��
��ꝃl��lrZ�:9<u�H�nrin+h��\dcsh{oOn ���vJ盳gf��Fݦ��nܙ��X��M�������-���[��}�Vm؜��g�[F��`�\�7l�㮹��8ř<����잸u�9�6�P��Y��j�0v��y�<�f������Wu��r�۹�ݜ��n�n�|u��ַ�^LD�8��moj��r�]����O;	;)Խ��푷&����˄v�B���:ۃ�����tV�n�E��-n68�gc����{=q�m�z��jG��i&-d�.'�;;�,<vg��'�3���@P��;o;{<�[��cs��ymZT��*�E�����[�_�@��@׬����ǋ�~��(��O�����T���
E�LT�ԁ$�O��wߗw��wT�r�T��`��N��j�V��nV���������������������������j�����������������������O��ӑU.����=���Ns"n��.Ц��t�Cُ"(s�5�2��na�2�<i�zِ�ӴVܡyIV'�[�l�,x��z���g3�L�Qy�8;z����=i��V��j@�q��t��%�ַC��외w��8��Ss���]��[��ۤxQ��W������6�F������c��v��Ƣw�WFN�N�s��G�a;/)��Z��J��W&�gnr���֋�wm=����hի ���>%�q��kn�wl�<���y�ƻE����l��=z��=zۢ�-�n����,E�sm�gt�s���c:���ź��67k�a��v;[nix�x��#o<�K�	�k��E&ֹ�B�퓢,���Q:\;��=v���U�R��:�nyz��2�O��_]��:��'�Aݮ�oiMțSuE<�Vӳl<�r;]k�q�p;yq[�\�^�W���-�mSL42�8���;nu�S��'&�Tv}t�ɠΌuC�yo Z�?~�		�I  ,E�q���.����gjF�����Z����.�#�FW��gqԇ%��r<]мn�4cu�X�qo*=�{�^1�9�G�z���ݍn.�i&3�tmQ���g���]i}�E2��'[vk�ײw{���W�`������9r8�y~t2�����A��O����N��,������������w�b��'�]�h����^�Z#f^�{d�|m���;ۃ��c �u��V��%�a�~���o������=Yi�YW���t*L: +�3���q͜R�u�s��q_rp�8�m��3�0�᪦l�(�����A��޻�o]�%;>EY�%�{r<�z+���*+�U��}���tr�gN��kbo`�:�2�_3������X~�=���X`�6a�q������3�w��4�FĞ\�����@ͯ��n�a�lj1?�����1�˷�J��g�[瀪r�cQ'�˻�]��Bk�;ҷ�sR�m�w�i�\G��k}ܚ�:_�-�4��׵5���͒Ni��5EgL�����[���x�L����9�;�],���X_9{��ۧ͒��D{��ʬ>����տ4)���(nb��t4nӐa��|H
%��i���;���F]�NJ���'X��yNr�P�n�%��MJt��׬Ԯ루��d'�K��n��U��8W�{
��g�(c~��a�F���b��H�` ~�q����8t:W�^ڳ�՗n�عۥV�U���H��//��f��8�%s;J_
�n������b���w�*���G�LxoVu��uY�]Y�I@�ԹM�e�v�zu���~��U��ylE`����WǃQ+u�P�e%����ǰ��#6���A�������=�ݘ������Q�c[�o��S��Cs���v(��m��P&iK����V���p�=8�S�8�R�IS&]�d��M��T!Hg�E�&>�D����T�;ox��z6�贑$w�(Ei�4�['��A6�*Cm�!���>�6������r��7�t�V�C^����z�9�7;�k��φÝ�+A2t��&�H�z�Gmw�ۢ��у�����/���?�羕��K��U3�sz �(C컰/��I ��h���t~;�,t~С^X���`@-��PI��Xӵ���R��{r��+�+G6@/h�\�v����k�6�ʿz�ٵ�|�d�# �$܅�c��يJ4���6YQE7ط� O��e0��*+�`6^B�˥�^Yf�{9�V�@����ge^d���d��m"�4e����ɦ,�}1J�^����\%aAQ/-P�+��K�c�ݫ#7��Z�fn�'%<4�AgI� '1���$�!�rUUUUUUUUUPV�%̖|]�|~t�e�u�ugm:�t���9�<�m�آX��ovۇ��ذ/l稺�vQ���#ezze�[�e��_@W n3 �=��l{u֮�P�Dm�A���l\��8M2eB������J���;�i�GO���E~O��ӈ���x@��&!��6���X�b˾%q�(�I���c�Zy=x���p����w�^4�����v�
��_`M�:xfQ���]Tg���X都�ݛ
Ij�8u=Q ����Ju��*mV�l9v�ܶ^멃;�RD��!���f���FSx�>6�0�l v��s��Rqs���.)��ֹ�|�Z�[l2*��I��X�vu�fm�m ��,��p�֝��c<�����{}�C�[��tZ|�o�<�.�4^m�Tm��U
�뾎��P�]�dڳn�y��]�!����#T��=�H��Ui�����0�:Ͳc�rDPT/oO����,��a�-ý|�/���F�'g�N�K?��C�s�z�#[�y�<�k�BF��'4̪�l��'D.��	TI��Sܬi �Gz�j)d��W�ä=ʺۯ3 ��X�a�
� CM�x�ϧ�t�����\��*�T�g4:��D{���S��V�>�=�T	�͋�W�W[&S��T{w�.�z=H��Q��tՊ�_Z/���E晽���	�i0ּ��qF�\r�԰B���I;�-��՘�x;�ݼT,Rt1m�Q�m��
}�4|��|[���Q��@)L���x��{m�������:�w�w��R���IVh��������m���t��WyL3�K��\�&M��)��2��!!	��S��q����[��9�[1^�վD�,q�����N�c�w�b5��>Ķw����:n��4~���y�w|�v�Ì�i��sS���lP��ڤ�(���=��������s{7��=���L:͌�7��PM����w<r�������u��n�Ӝ:�u��R�E�ݽ>lCO7�Û�I�1gU�X5"�}��S-�>t�׺�4Zd*$��'K���q2�goE�6�c��Y�Rd��@��h�GmL]�xh�uk�A�un��f�t�h6N9F��V�슝�/�K�6Fy�;�*��R����@����~/(a�;8,~���&滥w��=){���(�Ϧ����[�o]^���f�i<�;urKρt
��F�鸫{E{��Uj=x�@�2sǆԐ�)瑼�v�{Xj�26�l�����W�oְ]�3����{$D#Y�|tOc!]�r��J�Mx�ܪ�m^����0�V������抵��|#��I8��I��4Kn����Wʪ����7gu�4p���ݣWK����d���9�sA�D\z�]�l9�j���R�t.�z���t�vH��vl�=i����H�����&�8��&�����,�k�RYx)T���U��|*���:��Q�����ERi"�N�m�Z>��?���܈C�B�|N2�pԞw�|���j�N,�%rdAv���w��hJڋ�����?f�tM�*n�:a��I"vj�W ]��{j7�E�![�=с�(���$�L����&�p��
�`A	�U1L��]�V���=F�4�$���н�~��2�9�;��m�\E�>���
�����_6����� �m`ll�Ds�nŰ[�8��ڇ0�^]����T�S�^���>%J>�ܠ��t^Eu�����H�~eT�t0R1xv���kk����/g]5J�I�H1�9��y��Mޡ������c�(H��n<�熏rc�@�\	��;�E?ӈ�E���e���W�SV����R�d:t��W�VtS}5U=9���������5��8���57�k��*t��wf�m�u���:�g<k�w����B�LZ*6萁-�(wiǵ�q+����7:(Rl0�Eb�9� J��{�8M�.u,���J�C��(�'O]B
`&�9Zup�HCqK��0+��t鰞k=_z�:Ola㽲��8q,�a'��W��|9�p�}��D~b�?V;�$�o�����g���T������٬fo�m���B-��Jںλ�(u�����v��ܣ�����+��֕N�<,8�����&/ڻ� ��b4���um9���ͺ vV��o��;O����ͭ�f0��3��ō�ۡ��t��ӑ���єv�Nv��.w�W>��}zMӵ�X.֪seD6Z���pQKt4h��~���v�ի#���v�^�'xQ�Ջ4�ۋ�i�D&#b[]�/c9�������{����W��Z�XU1���Y�VvՓ�&3�����Za���w@;o6wN����2�ڍ�}u��;6���-�X)ٚy�EX�!
�ufg�1F�Vb��]^k��6�}�����V�2�k���u�[q
Y~�/n��kۇB�ެ�ͻ�:h7%p�͟��}�>5~���`��L�u��&�Mx�XC��<:���J;O�JM�B�Tլ�q����[���)	��ӄ �����.��A{��vRW�{�����[���Dn�"lw5�H}��i��	�E� ����\�V���<«��G���=D�m�_�=��Vzj�����m|k^���@�t�Z#8��`^�l����7��}�WBv�k��*�- '�s��t��\�y��Rl����Q�\kÙ�ߩYU:���`�X�#s�"����i��7ˮ�	��@�����&�w�-�5d���w؂_K�j����s�Ц���<w_{1��_lyP�eE�V�,7�ثcA3M���qY���|M����>/�+E`��������-�31�|����!��k$�T�*S�����TB�i)�� }���;�$�Q��BB�>m$"�%2J�ՀBIL�Y$<!- Oˠ�Q ��B��$��@w<9z7�ff^Z�tݵw����;#֝V�]C�HsNb�Yw_� ��
H)UR
AH)!�D��R�d�TR�$����) ����}�VAH) �7U0�m��
ACRAH) �*���RAH) �=ʴ��R��a ���\jZAH) ���tAH,1�2u��R
AH(JHj�<��
AH)
�� ����c������
AH) �7TAH)!uD��P=�E���R
AHf�Y����䔐R
AH,
i ���Q ��
z����R
AH,<�WD�H)!���Te�aw���
AH)!��
A`SI ���R
B��) �|��R
AH,?RCz�Z ���R
Af�]%$��ʢ
AH,�%$��R
AH]Q��$�j�^����
AH,�Ϯ�/��R
II!ʢ<�I�I��H) ���R
AH_2�) � n肐R
AH)� ���R
AH) �*�4��aI ���wņ�
C�D;TAH) ����ÙωĂ�R
AHUQ �����R
AH)�~[l������R
AH) �����I!�D��R
AdX���RTAH)�ݨZB�����R
CUD|�I�
H)3t�c%$l]R&2�
AC���.�)!y�� ���R
AH/�RTAH,;��k��[g!i�M$��R
I��M$���[`~%$��R� ���R
CUD��RTAH)
�䤂�R
AH)�k0��HRR��� ���R
CuD��R
AH)!�P��ʢ
AH)!z���^�+D��R
CuD���I ���R�]IU/�����$��R�$��R��0��R
Ad�) ��RTAH.��R
AH) �.���R
AHj��
)���)���Q ���$���X}څ����,3uH) ���R
C?=Y���R
AH)���AB�]� ����i�I �9����$.���R
AH^������!���
B�,�%$���D����HRAH*��Q ���R
AH)�����~f]�`��~ ����Q ���RTAH) ���R
AHUQ �[)�S1��7VAIHRACRCUD~j����R
AH) �@�YD��R
AH,�ֽ����ZAH)�0�j��) �2���R�$��R}P���R
AH)!�A�Jz��Je$��n�)����Lj�) ����Q ���R
A@�����R
AH,�d�wZ�
N!I ���R
AC�2肐R1��
AH) �.���R
AHk��?fUg�v�骆��k,7O9����e�h�v���F�D��j����������ܦ�ݹ�݈�k�M�E�	��emwL�\qg��ͻBg�˷<z�����%]c+.|\�v��{\x�f���`+�G9��v-U������}`��]����j�ٸe��h��i��9tt��6PT��3���S���Q ���D��R
Ai��Iڨ���R�R'L-�=`k�Y�i) ���l� ��)
II�II ��񱓌�aI �5TA`y���RݖAH)6�$M���m$4�R�R�T- �7TAH) �$���R
B�=Y�`RAH)��;����R
AH)�!�
AH)H)!��4���Q �aIե�Rst�R
CuD�
H) � ����� ��)!Ĵ�$��R
C=�q���̺���)UR
A
A`y���ʢ
AH) � ��������RUAH~e�AH)!��� �(��I � ���RTAH) �"�R!L��+2O�I �Mj�� ���Q� ���D��R
AH]PW���AH,����,��Y�JG�$7TAH) �!��a ���R&�I � �|�H)�~V�AI�RAH)H) �>��[��WDd��*�B��v����a6��B����~U��6����yRba˭��ލ�e��f�*ì��!O�*,�í�ۨ,y���ʻk.�~d��E��Qy���9������}���'�@Rc��VB��Q��މ1��+�6ͻa�i��i�}y�k̟n��2Z[�N>�t�����r�Z^.e�q7B��W���V�ʲ���M���s��&��d��^�)>a���<���0���9r����k���~����32��ol��v���C��G7F5yY����-���%+ԅ0�Q-<ɴ��yڸyv�B)�q��\*��N�Hi2��Y���Hy�{�[����<Kz���]�O�-��/�}_�~70���?,�u�e:.��t���,˾8__*\�p|�U����i�%��+�8�aWAIl��w*ͣ�\�V�4��bz��\ݷ�&�S��kw�X�mejO�kTc�8���'}GSI��H� m�|�d2�S)�=���߾��@�z�O��S��\g/WVwu�8Ϙy1�-��}ms�-&�<�m��0����3�)���g]��ZM%�������q�cI6�j���i�O�$��Iˢ,����ݽe�V^SU���(i礼��\�!n�ǥ�׏�����Iۢ���P�h�d|���Uj�>�}j���\�hr�[�Oaj��9��u���k���}Y7Z|��n%��Tg���ow�m���e�7�U�,�&�T�Cn��%3���;�Z��Ԕ�a��=�:�Hb�f�y_V��U�W��Jd�R��}]������/�8ϐ�j�3�7��dJd-���%�i�6ϨFUU1�f��+���Uc�"L<�����Q6�N2[ۢ�U��T���W�g�C]��\�y϶Q�_�}�O8%CGM�ƥ,�2�":���~�R�~VCI)��|��?f%���[!ݝ*��VU%�h!L6�Ϛ�S4�WP�kH�cL�T;�v�L���[��z��V��6�1
ٮ���d���h-�P���*���̩�m�)�Z�Հ�JC��﷩��&��gS�d�T~��"��{�>�JK�1��/�'�ץ!k 1��D�ڇI0��v2Du�F���n4�Yuc��ӕ�eKa䔆����4�E��2�ڲ�i)
CB
�:C�j>ټ�׿����y%oUp�h����i�|��.�UZ0�̶�~|��\)�~@Ɲ��d>+�ۚb�d�Y�T뉺����g�L�������L�ۯk3gs�o�!��ׯyx]�c�Z�Ħ�ZA�{m;C�8��1�^�\�!I��7��^(�w��O!H>�+����ܠ��#Tǽ<���[�5�Hj�����B�� )���=f+-)%�CW]e�^�HSBDB������CG����)�_��_�_�~K�����R�K��Kl�kgm�1p���h�}�k�U���ϟ܇=F<�4�Bۺ��9���g�̬n���F8�0ZO�suM���R�U��߳~���s���)�e��Ex�M]؜g�gޫ����Q�����{6R!.m�
�QW`����[��Ե�[t��̶��s.��s��;uyup�Ŕ��M�]Փz��2bZC泵a^��;}=�I��!m�b�>�C��9�i�{���тVV�h|�1!�ӯQ1:��Ve�i��+��L�
z�ީ18�(1�@����
v���/E��ii�u�e<.�̧(�|�KH��d���
CiI�_��5�m��]�m���^ou��N]VLm��L���m�5\��2�r���Ɗ�UZ�
��WRbu�wAl��U�Ȥ��ĞOj�T۹-��O��9�׹�묜�U�0���������*�a�f�.��T����8��l4��W�%�7{���n��>aϨ�#\�<�)��S��������㷅�;W��`޴�Zy��	R��[��oV���dvجn����PN��l\�UUUUUUUUU��k�)��h�&q��
���-�g�%��P6���\�����w&��nz��'g�Ék����ˎ�t��`\�磷+���nѬ��o(�����N���c�|_�X3q�Q�q�v챗��=g��y���8�H{tb���1����N'��>���g�R�~���뼩�-6�x�|c5�T�y֮m����HA���}�x�u'�R��n�wW�L3������1��Ɍ�����g:v��A|o�M>e�t�L�P��*MV�+;W �HS����0���3M�u1�~�c9���ūʬn�a�[&!HX稞{��@�ϻS5uzUJd_'��t}����i�z�g�d�
O��6^0��ڹ0�����^[�yV���~z�-�Wy{��q�ek�0'R��^�t���CMꡈi>�1�m13��z���6��}�4��}���RK����=�W����U�Ԕ���و�u����ʲ~m�8�����>Ih[6��Rޫ!���>�Q+�������ؠ�A,J]��v����͢�nn��mʼm���ϓ[�N3nou`o��(��S���N]I�Q���Vy}���%��$ӌ�9�&'��<�s�H֏�ݔ�Uu��IH|R��j��Y�1�w�^'����۷w�������Fl.��7l���T�_t���9���!W��:�j�8�N6�v������Ki����r;=�� �{�ݮW��s�I�$�L�f�up�c�c;U�-��h�ʁ�w}�Fٌ<��ϷW&!�ԧs�i��3l�AO�[L����Y�+u�>e2o��7������i�jɤ�i:��W꾳l��/�sU>f�e�^o^��[������l%7�k�����j����[i�T�Lo�U�AIN2��7̝���dAߪ�P)��S-->��NS[�i>h�{z3��_�c��6��{[�n�N:s��t�� s(>�t������q4��6�v��n�e'�y�3�USnӬ��K�P��x뻠�%o��yq~�bM}�����m1�!�1
�U�������N�Um6�E1�7F!�n�i�l����]u���i��m�����C+��G~�"�r���=���a�e.V��m:�&��o}�M3����R�yW �e]�4�ݷV�*�@�%%��7=��y� ������#n�M���U4a�Ԗ�`r�e{�r
�F����,N�L3_h�b��!_�&W�>�}V2��Uv��^T2��Շ*�14�ߪ�Uϫ�q>�N3L>f&�c&�퍮�cuWZ��Qhb3*�A�i>`]ѫ�w������g's�3N'�i*���P�)
d}W���:�1?]�esZ�U��UA�Z9f�q<x���C�v�M(lZ;rn����~2
u�Iz�\�
��Ii-%&z��D��p7��`V�V|u/�s�|�Ӯ$����,1'{��e����V�ZSl���8��LJ���5�]i������\)%2L;�6� �2��3��C�L�Ug��so�^�RL��QW�i�h��C��-<�xɚ�XE�q�[;aj��6W���JLީ��%?$)6̪<��~q�3��9�����Me�h>d�M�[�+��I�Ri�{�{tR37�\��U ��?Q��}�����~[�2�����'6Y�:4`<�˰�]�&~xat���K:u�Q?g�V'c��i9�a�W�tN��������86j�D�K�ȓ���E��|o��7�Mr����&%�-��Vu�Oۦُ��6��r�R���L��>R6ہ��"̛n�'�9y�!��Xچ��yZ��[i�PhCN�mj�Y��lU��K�U�*�d�nz���)�SXwt��2�:�_}W!��-
C{�Uۺ0��m�k(*La]�X��'~�2,��ݿ3�3u9�жeP}���"�T8��T�QI���pE׫�_J�QI�ZGLp�$���
dS���k����SAc���m%3���h�b|�cD�M�2оԜ޵�ь
`i���\�7nVcfRM3�@/�״��^�l�e� cM��]YS��IY��1�|���L�Վ�&!��X�~KI�#��X�8SuZ�N�l�8�q�f�۠�o�4��L����{��7o���)-RR]R��lӽԂ�ƾ�X�P9u&�<La���������C���������ś�w��i#'mh �wr!�f�x�D޷w��qQec.Vj�}���ɧ�"��Ֆ	��3�U��͒�#� �ۈ�M��L��sEnĞsͪ(�}��Tv`Sb����\^�bM�lHC�3iT��C��.���3��ΰ��;Hv��8�ـ.�_R��oN>E�ZQI_#����wݝ|�6�b��y1��=��|vU��Y[���"��r���E�Fr�vˣ����:������k�4�L�}:'�2�؏�c�	i�>yr[5yy���ܫ6����^ӽ�*x5�ݜO 2l�U���뷭*�nn���v3���ҭh��ց�.>�����^����i�G�z���۫/��]��3�j�{*��HI��vR��v�jul`U����8���������������������������������������������������������}��u��[���q�"��5f0m��ϕ�b�9�G�vK]�<8��8���<�#v�m��oQ+��'*��$��7D�p�����n�����c� փ��a�ї��l[��s�:��b��Ӯ0���pnwը�v�eS0�ۣO�қ�Ϟ��U9��֬�N����ݜ�zͥ<[u{p��n�[r��	��pom�wW]|u���w<������LZ��v)�v�u���7m'4�U��%z۫>�/9t�joF�ݏ7��뉺�����`�O�6����W%=�8�j��۱Y�V���oK�;�z���uჷV�jv��I�O����������]GU�=S��vz�8:݌1�,�m�ݹ�\]9�6�{�����vJ��6�/l��B�����[�	�v�Q:�p�v�5\cx��)�����8��%�h����3��pv��D�=�'^z�,ػ8{+�u��.�t�m��'=Y@�b	�;Qv���������^ݚ������������!�v�w.n���'&cA�9^.��̌��p��L�L�C���"'Z��nѫs���)ƅ\m�8��[���<�y�Z�v9��z�wg��(���vz��V]�=�f���;j�8��Etug�\�D6��������_���Ua�~�D]�ϝ$�TJHc����ϻ���=�!�s�5]��i��lد
zi���h:�i��7�S!���|n���+��otr���������[:��2��#u�PRZ��1��i.�������/d�9��q��X�^Uܥ�_��g����m
x�`򉫠��Ę���{}vq)����ut�S��$�*-R*���3b��V+���F�)Ц��KCHUW�e��-��T�<�S �ڸs�dP6�I^�-�����z7��T���a�ֲ�l4���o�m�aZR���>C�P�1�3���!I�E)*�w}>�����C����1�Mj�G>�d-���)'ީǉ�͸�CQ�����XL�̈A�(9=�Gx��{]Z���Mر���p4��������4��)��i7v�Agܨ|�4�=Pj���m�u��7R�V]e��U'�SS�l9������^e�u&�%�8�u�"�|.�V+������/�O�rhY.��5�H�Vt�@E���^�7o"�tEY�G����g�m1��qb�
i�q�<��VR�S�,���E�^���V>B�Y��gU����W�{#�xe�U�u��:��2Sl�i�<�f$�P�i~���
z��gh�/�"�>I����<�~f�/]����C��-�O{�Y���S�ǌ�U{��)���C�Ɋ��)>O��z���$V�M!_r��v�E�&3Z]}�[|�N�RZ�u:��s]��e�ݙ�U�4���h��QN�Kgޠ�c$��*No�ٴϵ���R�a���W��ɶ-%5��K�U�I�!���c��'�H�m��H�F��'燷:ʗzt��YX�Y��yTM��8�J`+�a�y��d���4�}����l�r�>�����������`��ZL��l1%% /9��x���:6�d�M8�C��fP�ϫ�od���B�B��\�ǽ����S���9���g��b{Ur�i�������Vs�W{kf���q)Jd�c~���)4��s�O�՟;C���5����z����*SP	Ӫo������]��������Ls�pĔ��P�m��n�*~~T��=U8�w���r��.�PX[O~�k����:��?4��?5E�*��P��g9Vm�
��q�ޡ�L��`RZQx�9��I� �]�B��������*��l�ǈ�YTRI�E�^�ת��eg괅3����>������?!媘�B,���u_|mKʿfaIw�j�MZ�ck�K�ts�5�J��ƭʮH}U
K�Ն$�h�"b���S�*c�3z�Ci7��Jx�?v��e�r���R��+j�C_n�}P=��R6������V��xYUA��/��-����<�0��|�|ww�J`�Rw()�Tj�y��3;W �i��j�멤���8�r�{낯X�R�����*�y�d�O��&���Y���>i�jq'{���UeXE��}��6O'�g��ӽ��
Co��'{z�l�2ޤ�*����u^�9�8^Uϐ� �����~!�ʸ[5���!IHgh��i�1�S-�~��*�TM>O���9y��ܽ����a>�+f^�{)��+�g�����o�Ɇ�
f����
C�P�gYT�(�F�7ߕk���ν�Hc��[Ʈ���E��r�]�i��~�����/�co�:a ���	'A�*��KQ��qq�`��i����'N�9��~wd�1�?úLW�����e��K�h���;�D�ږb���S�C���8��\�2�)��km�+�s�-4!g�R�q�P��26��l��V9�ҫ+r��a�T�#sa��
'�5��h�im�)�[��$L��js��7&��oU�M��|H�2~C�'�v�:��Oh}n�g��h�I��B1��bjwQ��vu-WgZ�o��"�9n�O�M�ȋ��R�"�rvÔ6z�+��4�/��s6>U��a���h��'E0� ��n��������ml<g�����3�X<�8�Ɲ��ޟp�l{t���:����,���i��ǘVx0�^�<�q�����)��4�N�<�+]DC#n]�Ѻ�Z��]�]u�i3l�UmöD�vmX ��"Y��Z>��U������N�=gV��+�@"�E�<�ԡB�)�6�nŶC�q�L�k���J�{�YY̳�ci[��5$g�y��m^�G)�i��Tұha8�tMY�Y%+*�*���_�|Xx���WM������sf�?�\��̷b�o=��S�F�gwm���2Z'���zd1��V�N��q|�kE��[G��TF���n�ތ\���O-t	���	�oj���n�v�ͳ�i��&^�Bh��Qm�@6�=�Yeu���*��W���o��"�f:��۽g���l��!�` ���f�(z𥳐�igO�����&��3Յ�joD��_H~�p� �/T��r��T9�����Vb�w�ɉ�猯��4b��SF���j��e��D��HP�yi�%�}�6�4t^�6�c�̅
�=���{#�q��,Lb�x�.�|K�!Ŋk��p��7e���>B��\\lAj��䗩2�i�λ�~�p�!�^[�6�ta0M���X&A��p<�Vz�[(f������¿�V��y����c�i��I��!V��|~��B��ֿ�e��H�;f���AXݸ�L�3�(����m�/ބ��utQ�8
�+�u�f�w�����Å���L��|�^Mo�%de_��ᕩ�'�|9�[M���H�6'8%�O%�U��K�]�u�M�.��Z���������G�����2v�=��~�.�G?vK�F/�O��T� :�J8���W��R���t{��l:�k��:A\�0���^+(��B���E�ԕ�[*�Xa=��5��nF���]�RƖs�&�����i6ۧJ�z9[�nsv�֞�{t�SH�D$C��6�Fd�_#�3ݖ�Y���[�t�Y��U��T�^���U��?x�N�n�d:o[�Nc!����J��&-S-_v��a�bY	�Ǉ��8ae%^�F��8���t���7;�0���Y���Yg��!V׮�e�QF�����/w}�vl\��.7���Z���n3wD�i��i����+Q�Ԕ����{���[\�$��=��K`���{��=3�ue��Ҁ��Vh���BH��g���r׌�(�%���U�d�����w��?s�5\𦭸l��X	L��� Muφ�$�t�2�K��pN�@�]%w�N]-V��s�=/�l�d���D�hV��T������M�1ꓒ�K����ֲ�����*�Y�a̽;zPw�Ԥ�����kMw��	'̭V�Û[=���ky�o�#q�>Ѫ2t����P
h�8�K���~g���o��-�>s��s{w�6�^�'ό�V��N�d���ԕZ��b(6�Mޘ�>���9��=�[m��kQ�10�������N��D�R����y��gu�lk�|aj<���|��Y��v�UUUUUUUUUI�Z�E֞	�i�a��fͰW�v1г�g\]����&q�[���y� p�ֆ�[�[>]����ٻM�y�wgL{͸2�I���� Dm�<n��V9��+��}|��W�OHW\�]��Oh۝�h\��eWN�M�i���ٍ��drm�a�k֑�wqb�����<�kp�QwQ��t���^rXWt����.g_i�)�%��2s})ڄ���s˲3B?Q�6�vn'�ſ��ʿʹE�t�&߽v�ҟ��!G4�y��p@����Dț+ �/)���t_2{��_i.�>��^*^�^�K�E+�[B����Z�4�Gwlw��7A�}y��+�׊�cJ���_ƌ�yw�FN�D�m�`RM"i�t�����KXF���=s��;:$W?sh��z���g&(N��Lw���zf�Ҩ�\T(��~,z��t��m(�J{�G���S�`+�����т謃��v?P���u�[R����'=_�P�[6��d�u5Se�Y���]H4�3k�HV]�.�Yl-U�/H��f\����<m�Ԣ�1Ei�paJ����
L�N��i�lmʼ�]ꖟHq�=`�I��).ڜ'�{ٺ\,F�۾�]F"�&�2Ό`�n2�D�i�JWva�x�Tp�]#|���+�W^���k��y�M*}���'�w�;�\���gE�΋e�h�)�f�Zh���0��J�e�����H���N�����b�Q�0��XWQ)2�ͅ*��n�=���7��*�N���HVƕ���j7�O^pHj���B�A�h^�4	=e"wc�e��jߪ��ٔ�%����ɵ���u���M33*�8�8ݭ+emu\��BS���[c���3�9�/3��V�,'���|�B.y��j�P=xl]�j��;3{4w]�����' �F+�Q�oC�]x��egM�S�2�\ɸ�1�q�,��5��:�"!`�n�a��ȷ�ַj֕{m��d�V9]e9NI؅�e;��
����/��4�l\�o1m+�Y�Z���Z��^��W6�`��b�n�+`����geop��jY�޶���n�@
zј��b�z�K����kvb���l��ݤ@U3/��m�� @ݞՊX���mv��)��{�	����C�ѷh���W/nQ�p�e����O��c�:�l-T�[���S�f�4Shs�{c�s9*N�
+dA��޾���8�zl�K�l�?z��nQ�C���=쾷*�3Ki�	�x��δk�x�x�VE"|���6p-x�oyԨ�MΫ <O�ГM&�D�r��W���z'"c{��N�4|I����\�����U]m=�޵���.�S����H��M��N�D�{��`j��͊p��z�
j���J�-ݕD���+z�h2:�����]�r�G*����G�:w��f�����S��}��.)�N�Gh[Fk�X�����]����;�ަ�^�R��q'q�47����j�GJ�?��g瞥]t�Fnϝ������������gsN_e;�ų��xn�|�����l�������_�{�婃���e������;v����=�o��:~Y�L����mh�ٖ�
#F_������~\��Vx�=7f�b��%�KӪ���`�� �).x/�Ey��fm樂H�(N��F�%�1OJM�m���mH^QT�z\�E�S��u�}
V��:�rT�3Y�z){�(i�+�Dt���
x�� g��o���^������K��`.�6þ�m&�M2%A�9W��m�6���i�Ût�5Juۑ�{�[�ݶN�n�#+�(��Q���@Ⱟ��5� �{�o3�U�L�B�y^��p+�X"������$���ړ-L��Yb���:r��ƢnΥ8�wf�����������Q�8,���Z��MnӶ�mR[������N+�!]s��5z�����{����U�cQ��hx��5����4/)��g�l"��(��&Wy�Amg��!ћ����Yr��<ܗZ<��hϓ�]n��Ա���p>�ݸ̳���E^\Z�¯)�7�=�yB�uu~��Y���<.������i�!!�Ь �u�^��zA��6�'(ʧ|6�����>�t�����'�u����A� �ޗ�s(�$�����{'�-�i�N����׵���#�'ba�S�	>����K�b���3�/*�FʖH'WT\��X���%��:�`*����<�����]fK����N$�`��@�t�z�z4طd�Vųm�p�ہ��6���;�:��	�/U'�;}��%�J�{� >}�-��'9�`c�*�,ߎ�,C)`���5W�)�}÷2�����B�[�n�ŷF�=��
Wm�C� ��圆�[Im
Z�.�eS��v��*9L\(a�4�v��yٻ�&���臉S;�T�$���d�^/Yת8�ou|MQ�3�θjm��7\�@�Y��{�ᯬ�h!�O���{�pX�IU��<Ea��Ю)R'�쬑�H?��� �	|�"�%�S�Z`���ul��VY�����V-��/�^r�6���)�
�U.�׉A����4g�h]�|�����Ep�
�Ub����M�����na��՝���JU7�۸X����g��б{Sn���:>{0f�:ݴ�]��B:�&iȎ�b�AvC�|��{s��G�*�T�!�:�l!�H�����-����b2T,�~��|���j�W\�t:��X.���%�ی���'2���&9�M��E-'�Z�
�w��Z��(Ujs���{zj'�����`�9��uC����'bv�M\pF��q�\�����۟�o����Z�R�i��Ef�[7�
�4�!�o�N�2P�R�hSy���"��>�W��>˥f��.HU�����J�R*�x����)�H紭��q�����\O��]�7���j���Oy�4�LG�V��5����	VT�_k^�4e�6F�o�nv��B�߮
��}��oe./�]W]ә~�C�fBw�lη7�b�7y��[���U�]�X�w��t�N��Za�l2J�%�sk���1��+�]���Ns��H
���:,�l�'��n���h�`�	���x��_4�-��*�b�>�<P���)�O4vR��bК;�M#�T��
�����f�%4BQ�
���eM2oL���3[��N���T{
y�q�x��:�D�T�&�q��3�@0�m�6�L���d����B��P���0U4.e���QM��i4��9&�/mn'ug���.�uN��I�����5�<t�������s��b�f@�S��ug�䛽���m�`���n��K��}�9K(�U�)M��eP��E�M�mU�k]2u�P�����H4�)���)�Zm��UUUUUUUu�<�v72�'b��&NΥ8��<]��Z�m��!�f�۴�'V�]T3&Z1rA�7c''�쮛a��i�Rv�:.�`���7m��u�p�BY����yvf�LsvՅz ؖ�˓�m�I��O.�Y�z����"A��"�����f�S �ʀ�߫�s;Ʃ>6ˣ���`��.ܤmK̲���ޕo�	��-�����5�[�a����C���5;��<�tQ;I�YH�^�2
"�#���nХ~4���5.՝i��灿�p�{��AS�AZFL�:��>�ފ%��㪥�k�ta4��O��[�Gc�Sm�Jh
�J���^�W��v�9��J))��r��^PF�Z��3��c�W��R,�+m�PT�.�ke��ط��h��H���I0Z7޴}F(J�	S��։�]gT��w�����˼-�MJ&�h�h��,`��!�ѯo�fo��:��f�x�C����Ӕ���o��M+�~^#~�PX��@��dϺ3ի�<�I/�t\�͖aXz�
����.�~�7TO�ZQyAV�!]�C�'�vj�����?RW�s��uM5Vx2i��Ί}"un=Wxj����ޝ����E<�
��RH��^���AT	��>��OL�8�n�3
�[�O+�#���(�|�U��y�6:l���`pڠ�N�����H:�]މ��Mv�}k���-�9G�ý�p��f�$3<�f���!��f�>kl�N#��~�r@3��:��z���u|�n�n�,��"��I{|��BгɡO�U���]��`��"\��YAR������*��wޮ���T�.�g����r��e��]1��m��9��+ݍ�W&f�ĩ�1�ܠ�ҹ�4~��b�]E&���(�M����o�܎���1G^��g��?Y-J���?\v�Km��(\ȏ6:�i��ѐnSH����4.�#d�"�g�T�mCnې����1^�����������.�J�^���i�Q��� �#K��Gf]!� �I,� �ǎ�\�$O����S���3c	���4���Q�Z�"�Iuf��:�]dg�ᥓ:�^T�3�{�wx��G7kv�-��׎l���]6���xll[-�l����G���/�c��)� 1�;��.�&����G��;�<|$(�E����&�*�{.�;��~��j��Dv���ӳ�\��v�^�υ�lurIl�������]�x�m��]5EK���u9f�mz�¼&��'��p_���M$���@P>)�Ƅ�(k���v�Ŭvڠ�C���뺥 �FwpW��{�-4�VP'�<�j{x���%�6�fqR�N���P�ƴ���8����yQ�ѿ1>��"}�}��=���TT��5:���۷���%;)$�,�fP�_����~_~f�~�'u-�^���
<|K���QUU��C��O�(�i��uY�w_��66��է��s�{ԸX�{+o��t�q1�nd�����&ލ�d9ognN,<���O�w������WvV�J��&Q�6��op�֗@e�
`X��9vJ7�ʱҲ�ح����YK�JTCo0d� �ϝ]�+��"�"o��eҔ�*�a�7O(7�:;�ʃ��&���F�T��4��h
'[��V��WB�j��*�bte�ˢ:#��l��:�L�eo+�.ڶm����זh�/]�7wgl�����|sLV���x6���o�2�	���뗅���m���Y�`Ԭ˼���Vc�����Lܓ���E��vXZ�e�����Q��+30�{jnf��I�w5�+Iѝ]+/_��H�iu��f��2%K�w�	\/] �l	�6 ��'( @�P,��$�!M�5UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU$rZ�`�\�Q$P���5ɶ�r���x����N���	�e,�\�[uܚ�ǂ�6�n�niլ�]]��;�EvŹ�ܥ�[�X\�vN�����yڽ�wlt���I�>m%�E��K�vzўyZ�ɱ�#[�U�'\$O>2���'\��ŗs�q��b���x.1��޲�n�8�z�XKs)���q=��Т�k���8�\hؽ���{-$lؚ��{Ok������m#��vp�mx꺲���^.4Ucٸ9��jSe�����9\dGn�ɸ��ݑ����vɝ��G��m��:�y�������N�v�˻Z6�r曷I��.c���h�9�ͻmsGmS�mi���v8��ɻ��o��t���K�7\�6;x�Zpns8��'��ӊ˺�n����fݵ���ȨC
{2��s+HK��F�&7O1����ɘ��f��6Ԧ����2g������'$\hb��r��B���\\<Ri��gb�ю˽���<u�`��wo��������������������ӷ.�]���zh��c��$�{se9���g'FGj�tu�vݝ��1�ʽlH8�iN];v�z�Լv,'cg�.ƅC���۝[�in��l���<t�C]��Ur�aN�#�cj5`�����=�]7B��VΟ�4�.���y�,�T��._�t���V�9��}����>���`~%B\���nFilp���!|�����U��{��4H��th�!O�o2�ʃ)r1�gu��������s;:ۯ48(�zS�;�!	K�	��SN�Ż��]���� �a"m�
��%1u��<R j�=��N�a^h0�*��������o��+�lʷ�]x���$݊S���U�6��ǎa������*����-�"�v��o��o��.���6�iX�:Ӈ��m�~!�Y�Q����-�n�y��Y�/c[�T�Wcc0�D�ԅ�O��'U*Z�c�1Q��f��n��B�.(j����ɹ�:�����s���VNT�E~F�w캕Ɲ��֎tz�s���~
�b���)�i�Q���u�Y�t��t^]o(������
UR��e��{������ٳ(�J� C���i�ϓ�(�_f�O]����]�l�Ov��ި��ȡoA�b�Ē�LW.�ѷlǵ\-�t&	ɸ��'����?��[d��tL�.Q�Cy���[����uIv�i~�UcB�@X�&~��([��>I�!�S|�?jf���+�g�oywPxRE6.� u:d0�$���p*gBT�����X�bȉ��6m�ű��'~��7g�R� �X�i'4��:r��Y�T���^��sK����a�|k�zk,\4j�/|��a�}�i��먭 D�:�T
"�8��dl�������!K�3s�I(zC�(p�*J?:��h��
 �U����OhM�zM��Q������6�N�������ؚ��.�{�>k�?~�3����ߊ�+KZ��t��=�;�o����@V�%���.~��R��Sen�%��n��W� kk7��ʑ� 
��.�b��R��b��	�� d򷥢�ePu>�h��Z��ڗ2��)��2yh��xjL�*�_�l�(%��JQgtӹx���� b��n��]r#Du���i���e{r�۽�Ѳ��4����:��Z��_��_<�V����Ji��$a_��5꫺j���d�Mވ �m�i�@W��=���]������'�Wk]���\v�#u��c�^�#o�4K ��J��A�Y��hԘ�i>ҷ/$��}ޏ#�o� T�����Ħ^�W��zӐ���,�a��Y���6�F�̟bqo[���/�L&��U�B�=
�#�>N��X4���t�^�A�u�t/���·��9Q�"*���^�X��m�q�ߜF�K�I�3=�CH�[/(�����M�K���\�i,�1�.�B��F���5��;=٘�Ÿ�6\G���b�A���Vj��Y�(��\�#@|�I7UUUUUUUUU=���o7ml���n'�n��9��7n4]gc�um��Nۯ<�)ݫ�5D�N��]w<����	�����;s�f��3���u;7n�7v79���K�N���n��Z��n�λ�]�kWV�/��=*Ip��;��ɾ����|��Ye�<({t�̉)^R�'UIo��x
;�G٣��ȅi[�{è�G�
���WN���w]8��ܝ��M[���l�}�}K_=~�꼐k���R~jϣm��J~E�ed�~d�$BH'�BnWksM^�̥%��y])9���,v*��z�Z�>��ʱ\6	�]/��9��z�Yyv �zL,w%��v��������
��4��0*���=����p�5n����F��u'g�;��^>__�~ /�l4��]A����װ
Z�y����<S��+�f���0E5ߗ�?��w�!���p�:>��mMDb������G��ƶi��U|,�-���)��:V�*#N�Zf����	gU=H&����Jchv��{�.tB%���ā�$��g��Gį��]X���F�*mMQt��>nAw�æo�����T��r���V_zK��Q�{�^�-=��+���F���&�I�6NE��4%{W�z�=��_4���Pm��ur�0!#Y�׺���鹞m���#N��aCS�J`�^,ݮ��Z����Lu�!��\yx�� ���O����,�Q�?a�W�d c��M6W��B���ƙ��i�1�寫*����� �D����St�4}{� �I������&~�B�&/d�}���v[n�ƒa\P�5����/��^�>��uJ6*��<�۽�ߠ�O���T ��p���,��`V�l�ƇY` |���ͽ]xG�m�E�:���1Vw")���,��M��U`o����y��ɻ5R��Q�%�X���P{��Tۨ�X�)~���e���*-n�ܼd�,�덖�L�K��%Th�T5���6>g�W�-ey��#%V$�K<�E�[���Z�SL#�
�S�m.[�>��4�]������i�U��Α����@�������ߙ�@���\��ݩ�j�b.�T�-��f�|B��x�E�$����p\�U-|�_i�)��x,�w����ėi�~�c��'d�\,�8:�Y¦��m��ܱ��]��e{��-�Z2��!T+ߍ*r��}=&e��|ny_�Kj��h�>�����V�lR���
k6���)ŝkvun� �;[�g�exVe�E҇j�, �����&Ķ����KQW�w-F!^Z�H32��a.��m����'%ҲA�)>EVx��t�%#�5���β�?۰�Y�B�b��b��Ц��t�f��b���/hQ����E�Cy%�t	_�i�[�N�S!�J P4��z���0��*+褩�l�&���	�h3PF�>�o�^y�ѽ[@"�=ʬPg���^�Mm+44��$�c������~m�מ{�kr���k�M�2dlե��-��i��������������j�L=v�pz����(vܦ�vJ�u��g�v;���!&�n*��關v����^70a��F9���r�͞:�q�-����䕰n�mֺ��q����^հ5Y(������-f��=���B\��?��Ϗ���xX�R����UJ�W�G3H�n��N�AUgv
�CbA�n&Q�G�����`�o7_+���_��qm����Uw�;��}�>a�=�g�q��fB���f�z�H*!�j�ε~�wR��ѸB�a NU4��n�p�6��2��B>���]:X�(w�ʀ��j��/�zU�X����K|��ȶ���z�A�Xi[d9��H�Ӯ�h�i�BTIF�P`5wH�.�#yi��� ��HR�	�(в8��NN��,���'���a��'��g��K�b]Q���~�e:tR(-ǻwMZ��Z)�?���{ؿ_�F[�����ΙG�n v���z�#�n	�ڋ���7^�l���B�I�C��6��yA
�)3y�ж�-�z��G��ݠ��A��օ
���U.4B'D,�7�VP\�\^��x��?������

�V����d>p�{
��K�\����+�z���d�ON��ne;j�M�݉V)�a�)1g��r޿��j��߿>�s���Ö��/���M�(8�nsǵ��2�j�Xs��l�Kۼ�ӡ��y��;�Qİ���^�zϫ{�ˏ��nz�3���$��GI�95��+4��W�Tp�=2e)���q���v���W�0Cڶ��e�B�׻�(���zl`5�e:w����}��u��������fe��~:�+#b�ui�ZO+|�*f�ÝYl*���2 ���[��K�����lh��� f^��е��&�ΛϠx^�Ռ���r������̳ʎf�m�"oL��ڇ2iD�ӡt9Iw{�BfTu%e�3el�����na8��Ek	�)�o���
�1����m@2V��Z�\^�dܥ����ɐ�7�DfE��v��=)�MK�����J��w ��>��o��ފk�L�GVP�yO(ٱ��vq�.���J�U������բ�]�ʇ:�aU�7F^���S�58a��Ļ|��^����ӳ�����l��y�u�'+.�-����+���wX�wr���o7��,omku�(�/��o6�v��xFuɋ�Gf�z�^6�D�����f4�{�ۜm����.ܔi_޻��)��?W�4~���)=�����y2R���utQ��`=Gގ]��-��������I�8����X���Z����Z�mʋv��J�� ٕ����!�Mz��F�D�|���><��ie�|���e������F:�ӑ�֭`M:��>������5�{W{���5�EРď_������i��,�ŝ��H�n��m�T�`Щ�X�r��3G��g�����[���!ƭd��dzGj��V=��Ą�S ���yv_�ڨbWf��˳Q�����Xr�7��Q�j�H�G�OT��l�nJ-�f1���O��aG�lڶ�9�,�S������]�$�5��!c2�P�@�\���![T_KW���eƅ1f�y z�%�#L%���:*ᖺ����U�7V|�z5��2q�E`��6��ע2/6�M�0q�����Mm������E�	�@
T
�I��	/dUܒ��؞*����zeU��ct�Q��]�E�G?W�=��.�(���xP�R���ث�D�L^�U���\�<�Sm���O�<WŪB��u��������
S
 Ey-�^n��G}>�N�*@�MY���gb�lԮ���Y<dDֽ�.|���x��龴+!RN�S���w��#�Tr��Vb�)nGVxp���Z�Aw.��{w|��:(Q���쩰�Then���m�Ӊ�.�"�n�=�۝A���?�����q�v�������������#�/mN�Ӝێ��睁��cgs3Z��m����]��. 7l��{r;��c^�7&�q�����N�j&�O$4uOoZ ��m����@����s6.(�ⲍU���������q�b���v'@vE��4IxU(���;U�kw%@�:T��h=��ߵ���:�,,E(�rMG�m�(��iؙ�:�0��ʉT����T�=�%1���?c�T�M^�@�T@]e�>j��蟱T�
���Df�
��S�
�$,!@-��R�)�H;�m7�������՚72�lC����;|����N�տ�ݿ�m�,�L���B��;������0��:�]f�+�:]P�����G��>��l�:���,�m��ͮ�=��R%��1e��tFm:�d�C~G���ݕ1T��n�U�IpmP���K�'Y��oU8�=�3k/^i�����?�'1�75^𶓩��1���	���4^�.����*�WL����7y$\<�GHC�*�PeM>�V��yy|2u:�Yw^��:_Bk@Hd�]ƪ>̆�*YI�	3�wݶ5��.���4�������-��U�㔶+Ou�W�RD��}��ҡU�͟��:���x{,�3l�-��z��5oO��"�^(�m�B�o�4Hy��ٺT��݂��m��
ll:i���WW���S(�V���=�vr�)SVA)e���a�/+D�G^ec�3 ��tV0��Z-�H|N�*��[ܪ]a�Y��Բ�,�E���I�_�6�3�:7����J��?*ڽ��Pm�s���p��լ&H��cl���_�ؕ�h�"�c�fz�t����{�:��U�Jt��6��W��/�|(	�/X���ڼ��c�T-�@4���ǵJ�ӽ���YǞt�9KWT�3����i��V�γeU��X����ͅA�@��i* �:g�=#t�+�Yy�J(\L-���G�~�#�����p+�c�?i������/5�������G�UڞW�i��R�1�[)J�e��>M4�FC��g|Ov�W�v��,E,a��a=��M�j�EJE��F�Y���ޤ6��j��#,ӻPo�Uho���m�_z��/�ws�[�x��K#�XT:�j���b�`�6�����$�ttΚa�>L� vG��#<O�0ޛ���۱a�z�֗�	���J��P]+�FX,�m�Bc���6�'�F��1���������ҳ�d�Q?�Z�Ӻ��&��!��tK��l�:�ݟX�ǟI�5W�(��E&Rv�e"�~	�W6^V`q몪�	!�����y�W̯�t��9����A R2��d
�n���Ђ���m�A�\�M7B����Z��}��A���T��I:3*#�B���W����gݏ[6k���כ��x�@�
��_�@���|��~qLES�>�mt�v�m�U�t�+5�����v�
�9)"�-���MՎS̄^p���SO�����as��V�~__!�� ��UUUUUUUUV��`��k۠��һ'�{iG�pkuQ4�qڳ��ݧC�eҮ��6�g���� |�W�`�.p���n�e{u]U'm�g�n�����`\Z��֜��]lU]�㔭r-cѵ�u O�[�L��@���^ת�XZ0��xLRǗ�d�����.� G�^��<�j�
�a��]���^˺ᦂ&��m�>4�~����i�87�z�\����񎙡E�*i����t��;�rWv��
�$'�[Z�0^T�A�h�E�m��ց���x�����(<?!Af�DX���M����B*5��kk��� �&���p�gFN���P���lN��s�oxz�D���*X^���_n �z�)y�B�Il�p�n��F���&[Fg�(�E:�#��m~��j[��=�n���yن��ۥp��NX�z�Tiy�t �Vo��v�	{��Vsܻ�U������.k���\�V=����&��;=�m�<�����8�X�Xr�,T�����2����E N�A����<��b�V�.�jw�p݃֮�J��Mvzo[]������5��B��uA� \�~e�k�XR��KX���Q�zY�%A��l�J����3o�����T�Z,!Ye��1�/�ճHQ�$m�V�|����Gi7� �Mڦ�69u�����Z�
�ۮs����ǋ�}�O��v�-s�9U��*��x�Y!�w�P��e0���4{����=�
G�+��b�϶�_��O�>�B�ד5�(뾝6r�n�~�X�>�:���T;���	�/�l��z�}��8�q�Q;{w�e��f��'�S�T��Q�vrAj�C�{�k�����l�B��k:�J�`wQa�y�{ ��x�4c���?��R%|��!�X}K��d;��P1�����Hg��ݦ�YdY��ߝ��?��sv�@�l^ݵ�d��`^��t�:]����]��*��Qd��{G��WvHV�fP�Us0e����l �i�D,��
���2��ܬ%h#oW�L*�g�.�+�B�^��.	7A0JFG{�.��1t�[��:o+0<C.ٔ���&��E�09X�����e��^����(�[��Z�?
 �]
g�/������(�}0z������gf�֛��!^>�RY��hJi�/8deuCR�����ln	�D��,G�?k�?;�����y����=��!���&�E���=�����Ǜq*b�d����÷�4���ڛ�m��2�x�T7��]�����{��$=��Ma4ͷlb�t��`��UzM$����-��|�]#y^1;��b=�V�,����e��˽�h�H�=�2��]̃�$]hUF@{�����ȫ�a$���I����
�6;.!\�Q_����;���^�&/oe�z��e�;�����Cn�Da�����\>�M`�Z���$M"Z�������(z��r�E��e�)�\��x��+�:��tUތ�:i.$��n�L�u����\��2�ٶ�%��BZ���'z���K��.�cE���+����{�5�v��[�8�h�o.n���h�"R���]�L*��T�3���M�q�Z?f�έ��خ�h���Cf��J����7$���p{P��ha�l�x����d�޼�&L�u	V;�N��B����+Q�ՙE��K�m�4*�B�]{r���5��f:`a�m��n>�|�-��4-w�s:���̥������جH�:u���ȥє̢_-�x�m�����ټR���8qwu�f��F�X�kU�;��1V�4�&�Џ{�%ql'*��;`ގ�qRr�ͶjV.�d�g!�s��wz�:�S��ۚƍ��H��)��	Km]+iVd%� �R�[;�����������������������������������������������������r�h�Z�^d#�O]��M��U��烨�;��;=\��4C3�gG� ����v��Q��s��1ͦ�g�q�#-��^�pk��cO<g�[nt\�ܷp�}#��$��[]&)�Eب�f�枭���;n9�����^��'��7�=G�y�3���>n5aq�yw���km�s�s�S��ZL�[��tS�.3��]l+�gd�z�F<�Nڈ͕;s	�;n�p�	�ђ�w8�+va|�<�ç\Z�۷\^I��[���\��۲jۮ�i�O�v&�ެۀ;Y�����]z�o�ޝͦ����h4G����r�m����I�nw:h��X��q/1:�����kv���m��ʊ��ױlǎw�ť�^�-�q����][\˷N�!Yy���l��rp��X�
*��	ҍ���a9�0�v���'��n���5uN�[���7�N��sSXr<l ���j�4$�0��P�m\T�u֦]�-Ӯw&��{��ø�{�����_2v3��UUUUUUUUU\"���l�v{\s�����6�׶��:��c����j9r��WP[u=��!�in1�gt�۱��wi9ß-���u���G3�u��ڻ����-������qd�Fa��j�î<.�c�I��݊�"�\!��B��~��]� ��7�Y���Kh���^�P�*�$p� T�e7�v�v��uU���E$v�7�D���w3g�ߑ9��;�����x����Bt���Ѕ}�Y�?f�o��ڳ�!�Pq֓�7���Y|=G��T�\47�Xp����kO/(�w]S�4�o.�G\_X��iJ<]slM"�e���N�}��=���>D����b����D��t�U� ���kN
+`�wF�6��7n��n�4NTG-���0V��D�_(��9}�DDE9yk�פ�y����/H٢@T�lJ'�]�r5��Z�B.��b�Պ5����i'��q9w6�� 7����fP��b���-U�������e:W�y|r�UU�'7S{��b�}cU�8轫�L��7��ֆ��� #,���C"��<�5�������ۺI.gz�����g�E�b���=B��>��T�to��h��8�\@�M������i�k��'℺!)l�kH����s�|�Y�m�PM��vw�u�<۩ĝAp�����A�H�*đ���4��N���:�ru�V�p��_�[�c�`IQ.��I�����A�3��^���@ ������&"|T�h���5/Z@�]�Z��>.��ܥ(wM��?z�T�F�N�u�q��OY�*'�-�ȪO=��ݠ��B�Q'(��;$6�0(���pq-���@�U�{'"�[�"��o*��6F6�.��Q5v�
�$+ε�'a�m��ޛǪ';l�/�ɄV\���,2ӣd*8"�]D��n�l�ڤ���@��綄�Ã ]�r�E�x�tt����7Lm+�۽jwN�i��K�n�=�!�:��ʩӭ�,�P�ʱP|�2���N���̊���B��K^�� �/���|9le6�����I�Z����f"�S��:y�N�[�ǎXoGH��L>B�;<S�}�WN�m�3�ʴ{qB���7/���
�=�p��DWV�;޽Ї�$��
X}��u;������y�B/U�
� \�'U{XS�W��|�S(��q�,G���βv۩j�$�v!U�tL�Sm6Ɇ��R�ڔ��v���]�����b�q8e��w�U���sr��q5�Ù0;�w����P�����/�1=R12C��)�<�v���oۓ�נ

>KVҸ��Qz̔�^��Ut�@���!Q����v[�B��|(h����
]�u�M!u���ػ��_#���;Q�e�p�Z�Q�0,�G��ØVŬw�^B��ʛӢ��Z�_QD�_�e�h�Nd�f��wzr�(��{Kl��;�۠�7�{��[]���m��6�:7�S:L�.T��<�~�v����~�Ԅ��*�����������;�����z6[v�W`v�:6\�4۶,�eD��G�Şzh���&]�QN�ў4�<4�มL9%���j�v�c&:�s����n����:F-j�ێmŐ%�8�<����c�,n�;��N��$J��4��k|���Y��ុ
��匩�.ʽ�3s�ҷY�.���� �g$t_���_XO��W�\��㴰j��w3�1��;=�[T�l"��.ƞ�5�����5�,Hhл;���J&U���<�4�	�SH�q>�Ve8�;�>�+��u��ހ�mz�%_g):�<[<@nhX�B�B���S!
�U�w�٧��V2Ū�p�׸ȵ�2�2�m�CI�H�jԆ��ý��6KA=�	I�D���Є(S�ZT������Э�*	_no�R>D��a�m��ɕ�xä���a�.�ߡ�}�WaN��0�=�}d�j�3PFbw����=�7�<�5]�S[�iտC��
����}yG4������y���3��շC6��ڙ��;^Vԟu��񡬛CU��.�*�x�Nv��	:!�m�~��9�
��v_�Z���v�~7''����d�F��x��.R��^�Bb�����Q�kb���sh�a��6�ww�.]ހz6�|�C=�P��X9�&u�١0Rta6�&�K�vẤxY.�'����|ȼ���E)3E��$y��]3A$kx=j�7�>��Q݇��@.:����}���e�����gV��� ����=�\RRL̩�Z��̿������gnɽ����K�#��LF���{����b&�y��u���5)|����p �s��b��<'dz�Y�&;�����l��o,�	T�9mI�ғ>&�|��eІ"�'9O���\�d)�z���������[����WV�W�Q���۰��:�'�w�ʍ���zeg�����LuI]�a7w�x�lN�M���0h6��^L:-�s�؉f�%����K�/z��T�'I�G	��j������mQ��xZ��l�{�,����{���wd������[��=�F����m��N�Kwl'
�7t�d̀�ͅA��P�kս��'=�l@$[�W݆�bN��oa�ُ�\�`�g՝��b�]�ۊ-H�)Ch?H�<��޻�k�K�9� P>*��oh/���)��cm�Ce�k��U�K��O<{V: �$�(:(&j#G���j�t�]�|m��P�y��Hy�������ʃ1)��&��GGO/*7'*#2+Ok��xMT�FWP�v�6-�=ȎAQ��H�D�
vL���p�����TT�|i&��T)�^�&6�4G���s���P���nu󮮞�����5�If�pm2�Hi��L;<�*��7��:��<�p�oZ!��b����5�����Ly6�u �Yv9:�
ىr'�a5���??S��_�lm�UUUUUUUUUG!�mã����k`��cnP���q!���mu���n'�c�_�~|>|�����	����vՆa-���x4Y�6�8Bώy7��Wm�-�
kwDk��6��]=U���������ϙ9�ى�N��w�n�V�	��C�#N�o�C�W<��՗���|�֢�Ă&�l-��	t�Q���dۑe�έ���:x)�	���y�Q+�C/3�}��$��R)��J��/��*H�Op����u:F~F��hW��tLN%��8��NT�@��I,�>�����tU��z��r�a��6�lO�\c��RhQ���=���B�OTq� m��t�f�ڔQ��$�X�N�`�:�ʩ����n�c�Pz(�R��C�ⷖ��|.?`�l*σ�w������Xd�^��E���+�s��,�N�oi�.T<�C[ >��v@�8l��Ě#���q8%\�*��,mYL���D�#�ps��oQ���-w�R��!0A� Y����1f�m����$w�>/ug��t�`�y��+��+6�3?#���z�=&�Y��[�-Ֆ¾��,l�g��R�n�z���E�)�jdV��c��[�]/ ���^.��a�yG�u`*g�3נTt��m��ݘ�.���z��^҈��Ɇ)����BCgy��s!V�T$;=�k���f\�G݃4�NE�V�
��R� )�P��c�m�j5\�}�`�m^Ƹ�ND��Pɻ��ҏq��`i	���sʍ���'�q�S�5�~�LK?Z3����c�;� .���ɚ*d�����[�k�'���^���[�b�T����ۚG��/5u��1�U�U��E[���ސ�@>'�h�:�-��eK�Ի�֠�-t(�ӻ��c�ж�Mu��"�*��"���i��x{ve��b���t%\Y"򰻻�7�]�b���wr�@J���]�kl=緄n�<�Ix�b��X(/o��}�{�����K�����mebǛ�z�un�偶�=�]�s#c:L��;-k��p0U�3��es��P�sEK��W[��/[˟j���7ՏD�:G��*d�$���}�Cu��v�3p��`���j���]��k��W�F[wN��q�G˸d�IJ7"]�-ͧ4r��4��)��&��9��!�S��J���得7���	�� |5J�-��LP�(we�I�n��0���)���J����}�/�ߺr����3�2���"x���J8�U�x�$����6�".0#Q���:;Gl�h�n�����p�;4c�_��"��v:E��ǿ]`�{���8Ө~��媻)v�$
_��������$VNM�u��\�:O�/G1�{|P����b�t
t	Y�����;(缷�ޭ���Oh��w�f��5)��&�,�h����f��9<����~���[&!=9��9�K�w���)��fN�h����3EB��<=ר��]�q\1aXJ�X�MS��=4\�o�������b���+{���Eu�=Wy�a�ۗ	�r�-99��X���a���֚m�%�������;FR�v�![1�Z<c��p@=��à�G�կoi�ST�m���9����X뇧	��	C.G~�H;�Ub��N��u��H>t�;��I��P�z-o�V6��������<��
i�M:O�h�ǻ�p1�Hy� �bwC��B�(�~��&�,��i�@�X�-U�����,{����8���F;�{u�	i^�q� V��.�PR�nnٟ\��.tpm��goh��	ށ�Hw���o��F�����������x2�v�>5	=Ԝgu:��r<�nvG��a�Gy�TWZ�{vz�ۑVݞS!k9K۷+�Ev�wطl�qņ����"ɭqh�e��/��y�v�6�Z�Tn�=\����젖�b��=u���l=s���~����X�K7�z�ĪǛxz��N����8}(�D
A��G&$OZbMݿ�@ϡ���
��L�>�6�VOF_o���� =������UdK|���6����S׬֋��|�z����ƞ*ih��®zrO̾絑�Z���m0Z���)l��>�����o�p0J��[Z�g^����6��ˍR�@H�����{{�ooW�^�Z��U����Kg��5�͑ݏ-�!¹3Wi�P���?lu_�<[`���E�!S�Y�|���x�Vj��4��:i�F�%x�f�=q��wf��^<��Z�z�n#D���`�V���"�UA҆W��&��X�(��w�6Y!�.'�p��e紗���YT,��'R�c��f�u��8m���l�����$�q5�֤�Oz�:-�A�l�E��֌�<MXӧ�w����0�$w@ �*^Ovf��B�
��
�@�	E�\�7m��~<x��T���j��k�=N�ߍ֕���\9����������Qn^�nv\=�ݣ���u�k�~��?O�}mwB�■AB��;�������T!҂Aw��>��%J"�[����;Ĥ��ud��X��p����#h*i�`���3�f����q{Y%��n]�x�f�v�#���/���F�x����Oy�K�P�����ڤxB!�e��?n�ޔ2��<��E�'l�`�`Z����K��?��iN1`�wzs��m9D�1���k���,.�R������8W�==-�ն-�v�a�mׯ\қU�?;��������ݟ�ŅN!Q�~͞l�k�C�����V�ff�A�n�@�J���/=
�wu���~���t��u�+���^R�n�I�'��G�oA��l�Y��,�vλo.S�m�2��QФ�7g8�fzv�jW��üX�W���V��!U��wC��]�7��F�Ѿ�84#(�[�cڥ 'P���Jtn�$�>4!Y����+�wn�H\����߿}�e�Ur�D�;�u:G]C]'��[]��:�:߯������sλff�|���i�y����m�j�oA��-�ɷ��
V��&�Z��~�T�����ʺ��}�F�����Ze�g?���k{-��}:�h�u�3�'u;B��MNU[��WdMM��j�ہ |���W@cOݗpV�.��{j
�v��AӤU�^x�E���m��<�',�n�E�F����uug�4��Ft�n�G����@��\�.�>���T��m	�Al�I�w��A�媪����������yk=f����k{���f���T<��<����*�Z�M\�
�,�;sbp�8��R���ЧnܻI6��tcuu��1��͢ ���og�x��MTC�7�뵝��%����O!q�i1��f��qG���k�wN��7��թ���%P:��(M���BI�/�P��z������Z�����`-�I7��~�P�l�A%m5\5����]�d�oW���BO;�t��U������eS' �`� � hLK�U�(!H��h�~�r�"�lL�5��vMm.';�س
;��\��W���1�U<ں�G���� PM6��r��v�:Mt]�ۛ����-�{� ��Dx�&���&qt���}=qu:�wQ�;���%��bǫ�r�����}��Wh�GT��xp�Éw��Q��g���S�6� �����뫕A�@ݒ<�*j�j��^ɽ�T�D�t餓�b(�Q
�E 1X���� �g7o{���%�2�:a���
TV������ïlb�V�}��}=ۧ�ҫ9�f��I�4WC f���)�2�T���%�o	G�݇{ń�6�M1$�D&z��1�z۪gۚ��$�
��mͿ���[<I����q,���j3���+`��`��ͳ�:F���ծf��R�X\��_@v+y�se��S
�H�wi#}c���.�b�M���_P����ϲ��Է�{�E�Jɒ�{���-G�N�Z]e��
����?��:yIҠnP������4����.�zV	Ɵ{���+Ee�w��6�N��c��yt�Z5���Iw�[��C�#����M.��C�,0uwYۿV@"��$U")�a��H��M�|�:q��;q��KLk������.K���&���u��=����Jz�7qa�b��>ATA��Fo��3�����m��]K���!媫���wH����� �O�}���MWY�7ֽۏ
}�R<oƭ\r��==��������6�\�:���;�= ��d
��[�P�]b晓p��ڔ�ff%��\Z���,���Y�·��M�H�l�,�M�e��Y��ՎF��T�w��;���o����~}S��9�������X�>�ccs�5��z݅�����<�J7�>�e��V�)��}���i��K?K��IJM�}܉��:�N�y[aW���e!G7|����+Y�f�[_�Z��(n�تO����|lxGRN�:�񃄆]>pJ�G���O%���)QO���ϩL�GK(t>�Ϧ�-tt�|��x"�e��U��&��^-����罷����U1�p�q+��x2c���r'L"1$���ґT��
ټ��ִg+6����mgWfⵧ5\KB2��]�t���l�_�_��'�.�@��֥���'Q�^��|:2'L�f���':�R��i��$����B���e���y6*�t3�)���&`�\��,)	�����)��4���Gpуpf�ܬ��t�.��e!�R�y��u,c4-��v ���cV��m��$� "�lw�J�]�OS�=���h��5�U���CT�����ۺ.��ގU�Ҵ>W��a6��y��wm�J��W���푫.�����-n��u�&7�n��Fѻ�Us�vP�
�����$�μ.���yM�ӡ�
Yy�WV$�'r�D�H3w*��ue�f���s�� ��ǔ [m�e��c ��Ɲ�hbMA�9�	����������������������������������������������������[[u�@�m�;�N�x%w/n�N<�SY�u�[��G�ص�{%q��1�u�9��۵��˸�c����Y�^B��h{9c��^ծ����-���iz�6���q��15��:�^X�^�a�Z7:1�uW:z}��s�����'��fƦݤ��F#�lϙ�ݎ�{���ɀx:���%�`5��hv�p�=���H�n�u��E�:�]=��e����j�kv�k�����u��I[c�-a�����c=q�r�6;Riv-�����E^��Vvg��[u��X�Xľ�Rw1���ֵ�g=���&�ې�H歬��[�y��
;�Z]�7�x3O"�Z�U�x����e�c<=�����9ǃT^{;���X��!瞚�s�3ېT�����yG5����]�FR;=#'5����\�����k�;r�˲��A�;v��n��K�9���F��X�4(���r'������7��9�[�f�ޑ�%�Sݍ�B�۬=o��|庌�+��t��j�[�����h
������������>�����k�������u,.��<���㇓��u����WkM�懬�Y1��uo9l[�^t�6m,!�q(�t��ٵn�d ��Hںʘ���K�^����N�����k���i�]غ��CH��j�?��~���y�mNS�Dl�%�x	��{�$~+U�&XT6Y(�O�?u�R�Af��xy� +�����	�)��x��(���OT��X��sV__cO�Պ��J��lx�����s�]���G�n:>���י����hG�!���(j����n�]�x%��)�]�tx�h�k=�,[rŤ"A����l�"wf�K��c����|u��e�_�6�$_�j��������W��k�~~�Du�^�c#a�f��"R��T�Ӟ	NWe
�Q	��/XJ�����z.uX�ڻ�ʾ�� �ʖ�U徒��m��ӎ��ʇG��ٌ�R�En�®@�ѦJ0pv侳�9�n����m>W/��
 �O��	���o4+��w���x�� ����ux�{<�*��vL�#�FfW�=�����[I��,�W�EH����w:{$(z�H֞^����u&cl
T���j��/�k6�.��p���L�xo�MGM�A��t�-gGE]��:>���s'M�n��!O}q�זP��bM�1�#���⠻Ic��ܑ�z�m��d�ځt
tN�ma�^;�yK��_Sޥ�S�Yu�vu��5�]�b��!��ep�"����3{w�r>�s�\��~©�Ӣ�m\��b����'���痞�HH#6w���(72w[pN����s��7�X:�+�N��ca�6�2���u���]mdZۢZ�U&��QgG6^�N\��Ma��m	M��&J6��W�e^D��&���bsx����<w��Cz�͙�6���ޅ��;�7���U�o�7� )��I����Ֆ�(p�K�
��{�,Q�P�q8�������V�LC�i�����t=	U�]1Bt�.��6�My���Jj�v�}��v�7�Q���Z�[�̹3&�Ի/�+W˥{���B�:uw�y����K=S��e@n���CT�zzJ�|m� F������إ7(��^͌Q[O^]�XבL���4�.�� \��>��k�/�����}˥	��,��b�0���[S�O��N{~�U���/�e��b=�<����B��I�Y��.�5��;��(w%|�j�gou݇ٽ|�L7I���7ݏ�[�CzkY"C�xH�{^���%'ζ��"�t�0�^��(q5�/����R�]�y&�{"�W,�����"��Z�χc���/o��1>�3:���S��_wT���4���hQ6�UUUUUUUUX�K��7j���7-<��u�[:7eϷ�C2�<����3Ӌú�r$�WP��ǎ�U��������|=�>I��[5%s盖�$r�����njQsccu�z�;�.�<�U0��=7[]vي�Bx�q��F��ϛ�"��?w���|�O0�g��(���{x
�n�Kq�Ȝ�L�E�{�����������������۷�뗏9�����2z�r͉J�:M#�D��FzJc}Nz���tDј��:<�-X��x�Ո�	+[�� /e�F��5g&x�xSq3��'�s�_Q�w�v�ܔ80���[��~��k��L��ݩ�C��;�x��<��k*-�5��wLѢ��!���Y�­ka�6+T�4�?�C�	K:)����I3|4--��c�w����QJz(�L�	���<��]d���α~��i��u~�+O�.��j�.�������:�{��R�]����u����fstb��@%["*m��i�d��ٴ��߉�1z]m|e��ف`�2�|�m ]E]�Q�+~P�h���ڸ�4+�`� Gg0���@�1A��}F4���Q��GR�������X��C�^=w_���3���(�UF�|Te;c����=��My� ��YE�{�D��������>
���Q����X�.�U1��+����Ӿ<(WMz�w��-Ǵ|BԷ�ikz���h��4���ѳ3�T/�ۿ<����w]�j`@]��9b��_ā��.'2�v�Õo���ͫ��d�C�����͠�T�k}���K�5��N^��W�FV���'�P�u��*va����m��R,�u>R��uO^�w�}�γ��[�Ǟ";w3�`���Ξ\���F8�{�0t�I��HQa$@-�X )޺z�m�%��[� �Jܤ���=�L��0$�Etz��U�}�*yh:�c#����ɴ(����*���Mψ�ä��RE%
�x��4��8W[D��|n��5�'���H�I�nyxI�M�;��$����a@����
H�[���2au�3q�ތ��n>X����j�2����V��+�?�!.3�y�a��5E��ts�P[�^G�|�^�sVx$U�U�#�\.�Urq��c��	��S��4���L�`�C�b2�����"�	���L����|�/9^�`�66�N���{�C�۹�A/L>��x��ٗ����w�H���ݜm�[{�Y�[�ޓ^���2c6��;�sֲ�彳=����;�/Pt��A��U	���X����7C��D<5���uM����q�$�Ⱥ�! ��(�d#��X��}6_���~����[cm7��q=ZXtr�����0b+��^�+$�~�����UUUUUUUUTc`� gg���Яq۷=e��ݬm��·��8Bw'>�n�n�mw'vN<��eS��[G��sl�!@D�qۚv��<�g��k \�x�=�ۧ�3�6��j�8aL��cXܹ�� \�Cŀz�e�����]��7Zt��I!�I�pu	�]��ƃ\P�.�Y&�ӫ��@�I��V�ҽ�]�j#�y���r�W%�6�REw�5�zc���9�+#��8��-��	c�л��&���M�W|������ڽ.�"�pß�����~���Up@�	��}���J9��8!�|]�A���v����O��M�=z�;>��|��[l�4���ЧM�1�Ft(A��CnP���)Щ_n�_���zd��7R�%��u��e@��=���>A$���E�qYE;C�uqC�$*�e�v�{Ҭ]��5>��%��b B�o�ѐҲ����3��g�"	x��H�~��'�ZĮ�v��έ��AUo�n���e.��`�^��YRH�<l�;[��}#;�]�v�����ݛ��f�5�u�7E:M�|IK����o���EI�/RF�X�es`��m�tH��4�M�ź�t=!�ل�v���4K&h��s#:(��!g���T[�]~m�no�Q.��_�g�Oò����=�X������xq�����R�x;OG��"�w�;����Gy_]�/��ܢ�u�J��%��W�.�{ �wvƫ�S ��M[{x��E�,=[�5j�R�{�][۫�tY��b76a|%Дxe	P"�2��_��{靯wN�\�����蕹6��&�N�f���X�:��C����V;3�Y�qT&��1J�{��쮬�gP�"kA�So�}�-�ӁD�ގck �{
��%�L k�{�Ȼ:_:��������f**�KaN1�C3��̠QD6��0!x4«'Y�͕�+���3&ݐ��+7�qf[�;<�ॗ[os0�Ұh����կ��j֊�
�;.�VN��TG����Y���L*�/�!}O�X��4��%����׭�=���p���N��V��2�5�<|_v��Z1S��v�M�6�[o�3s0Y���a#6����#K:�9�O�l�Yɞp�x��C���M��'�������>�J���2N�kΤ�:h(p�&j��l�Q��ڕ�F�H�<�^�J����D�(�M��H��My]&}��v������$�4��(�y^�r#��n�(7����w���|�=�s�m��h��VF��MwX�V�]��h��o��
\	iU�;K��L����}~*B^n��:���w3mk4��\���}����i��ݖ�wβ̱����OK�z��Զ6��uX��ы�m�ۦ-H��`vSp2��Qu"72R{c�{����.��L�?���֛�TA��/*�[�vMy�*���ڢ�]����D��p��q�ւ؊P���}���}���7��.v��P�r�Z�Ex���kT;=q$�S`��g�B��{:kU%.0V��B�67����sM�;#V$AM�
̣�:�b���x�x=�/ÉU?jS��ׄ&�&�F�n��w��K0TZ�\̬���}��ﮗ[c��T�4�e0���dk�CՑd�ɝN��؊L��]�����|�tƍ�y���z�:��0	��#��7�����µm�;�,|�a��m��m�ꪪ���m�k3�b����k�ԍf��V��9/��Cv+v}uFԓA���u���]:�&z��N6�gcuo:�S[�Z^�֑�D��U�jS�eꌭӔ��%��k�� �ܚY%���]�3��GX�gWd��a #�Bm4��M��#�Qx������.����m]-����GW�Ug�*�z�X	�u7�x���>#z/5w��Lo�kn��&���ABX�e�n�?=9����b��Yn�,�)���Is:-E�^�/~t�:E��O��XY��P�bYU��5|��G�廊߮P���)��F�
s���e�u�62{�����qH��o�v5�ͬ�����q��7J�x�{u����[Ả@�e�4l=4;J^�we�>�"e��R|��R��٤#)�XH v�I�ժsz�Q��;\����
��I�E�6����ws"���L�V,�&$ݻ�է�������R�!��X��i�������AB!|�s�u��x2�٬Z��š&�)�p�S����s�ӣ4�-N��ޏk���ۧ���Y��������-��^>�W^���<��Y����pl�q��h������5
h��˽*c�Z���3Dl!�՚���[����w-2l,;O<��]c;k6�n�  �E1�Q���w׶�v
K�h�A�{�+��y[���گN����ٛhZ�e����
�����vz���2��\xgʭ�7[�j�]��Q�*i�c���/�;ą�$l�)��;	�#��� %=�\(�r���Jz?K�e�K{���T� <OO�{[	��+]��E�75�) |g���o��m�PN�i��i�\����:�nm���9k�X4�ބ`xgc�[�⣨���3��;�g7qي�6g�H5A��7dC�LyZ��l����z�	`p{�����V�����&�����gz�����eu�eǍ�T�ot����:�1R��?���5�~Ϳ�{M{O��obT%K������*3����/v�݌�ʦ*Qg&���,���т�ٙz��q���7�ϛTS���˱�
�]��k��*�GS*�ץ��(��tve�4�j��b�3=nا�L�3ׁ����[�su��������A5��%Oy076>��D�<��3�'�M�C7HO��J��u<v�h��f��v�]���P�M����f����4�]ί��o�׹ٓ�Y�Hslm&�m�q���&iz��m�ƍ���vkNZg�vG�Z��a���<���/	�@鯮�{�q�ܲ'�TμhT��Y�曷ٔ�@-޲p-�\Kf���G���q�w���G�#�.V�UUUUUUUUUi�o ��N׻]��m�<��x���8i��u�mָ��u��G�q���l]Վ�������[/`�7�Q�8//�����3�&�<uk�p��1՜s˻]�k�N9�*�s���Jo;���$�&�6�ex5M&KVOܩ�64V�_߯E1Y�B�������KG�SFxF���
�����1W�ޓ˜� os�u�p�[Ts�a,�JtU��w��ͣ�oU�n<�lö���7ҡ��dL�cM�j�۞�C:����^� zN�>���(�4�\�!$������ �}����FiL�Eg֚�ex3^򄪭Dv{]�]�cCo7z��;qaz\֎"я�����6&���f�w��<�����b�p�J�l�Z���S�?�T;19����RGc��V�b�\�-ڜ6�� ���J�a1K��.�w�^��.��G}:���mG�0(X*��Lߍ!˕�����Վ=ק��Y�V!�|	T|��p���6+��?�zBwo[�E[�p�[B�J���,�ϸ���܉/π��2����0���T��?�O�U�mP�*-ɲv�PF��!�Τ��h��O��¨~� �Fc��6�$+�GU���-��rj˽8��h��D27�$��թ�g�f<�����D��a9%t��QT-�;�%�«�]E��8Gn�w4v�J�yݱ�
�\�m���,)3'WG��̑]ڪ�oU��I�E����;�ޏv/��g|@�v���*��tl����P-t!��^}c/�����G;ޭ�0�:�:b۰����~���r�u[>���#v"ƺ�g��h�A&n.�G�6��	���:)�qC{�:���� ���ci.�l���)$q��B!㷛>c���e��!G�]uΒ�JK?][t��7��+�X������z�wݑw'�q�z�BE:	���'��3k��a��;f�����Y�Mn�aev�] ��&��"�Bl�n���M3ol����=�:�)�0�6|@-�XH���_/�w#��Zk��i�mk7v�U�Ȯlm��)�g��.�uɵ=vx�tm
�h��}8{}~���S�1��v:pZ��+�L��m6 U��U�W|��\XU��Y�K��{�v�W]�X�|�6YJh�%#[��5�\Mn�h��@��4��YT�:#"���=Y�ݝ*�;�;�+��s�1�TK�!4���.'�J�㽻����4�jf���j�������ʊ(���!@��l����6�V%�]�J�wy����� I&���5��[��� @܅���IY@��X"���J K9A���T��L������@� q$����?{\�$��������j��Z�2�2��ݳL/���,�� nI¡����%+�zZ�7_]S��W9(�|� QJ�i�S�V{��l�X�Ŏ��پ\��u�V���lo�"Hd+D
	�'��w��A�d���S"����Z5��]^FXc�\,�32Q����7�?�O�HPD $�܄	H:��,?�$GZ�C����4�g����� H<~�4ɗ#{�[w}���\%����oZ����؇����O��������&�}N����>��g��n��RȴT��[��}%oR��im�zx]>oIjn%�M���c��.RӤ��M�1U�(R�K��R�ױ�SnMe��R@�C��aSf��� �I�BH1��'ą�?_�@��H(!{@�HoN�0	��%����oeו<Z!E+~�7z4��\�����\�_>;�y}�M5���	��2���9K��u��w��;�E+�t]^��%�+ag�|������Z�pܞI?i����"��tP�ID���$�9^k߿�Gb\�{&~�N�f%�q�:3�v'��9��ˎ�v�X/6�vz�FS�3��5�%���uY�TY�����p�VѴY�,��͕Z��;��~�_&B	�����.�p� �'�f