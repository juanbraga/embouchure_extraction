BZh91AY&SYl�V[ؖ߀`p���2� ����bF�q�O	}SM%�c"@&�4 ��@*�((�`��!@!��HP �U,�(� ���4 @ �
 
4 
U(B�Pm� 
4 �"(h�PQ��R@EU�>         ���"EJ���A@���־        ��\  AB� �j�ê�:m��uԬ�6�N�uU
P�*\�ȭV��ٻd���ΔN�
 [�F��Շ;m�{�^6�^���
u�vҴ���m;sj]��iZ� kD� (-�-CV��5�"�-Wv�ٳlQ j�HQ�Z6�M+*���V�V� �LP��E�hj���m�ԁKU�5� ԕI,5�Ң�(��Ci�5CB�P �����L�6Sf�Y�06��ښD�lCH��l�f��-�M��%-M���l��&��-2�ɖm4�d��1�`�ŭ`mhi��cKXmk6��QRITh@ U JZ�mY��2E-2�h���4�`%Kjֶ[m�!���� �l��Y��-Kb�-�cQ���R�cKm�i���j���X�`���($QZ������2m�i��Z-�Rb�����3�d�̢��if���f��AkV�m1m��Z�f���,i6�*��%hՕ �f[59��6����i{7� ��R��Bb��A��h��,�l��C��(�
����bki�-�Y�QiT�V�j�&�kV�*�̪�Q�9����Mۧa��4ta�m�Vʖ)mJ�mSj��ͫA�Z�����ڴ�!MF���m��Z�K%�3Z6��[�*6�m���Pfl�֐j�	�
�
( ����6���Y�j��-j�KM2`6Q[j�Ye���)-5����T���l���l@M�Ii��[M��ͨ�mV�eF���P �(U		���mf*�iZ`�f�i�
�A��h5�Uf��U��f�K-��ii�`��KV�mVm���T�kJ�h(Ti�$j֋Y�2�+5�+��5���ei�C-��E6���ɣE�1�j�)�-��iJ��36F25m��P�P  U�>�"��'��TA� �� S��$�*Q��   L5IA���О�Sɔ�=ڣMʞ��S����P� CF� I	��SI���@    �P�*��� �   �����[�p::�����1� ���5�y��Hؼi����Y��d�!In�:�jk��$9��!�I$5XyRI�u�I$6g�U��Co�$���O^l���d�����,%�c��H���� ��EdZ�`��;���#����bA��S4�1v��Mv�7�[�NܤJ5Y���5�=9ڀ��
�����6�Ή�ݩX���6��vmVn���arL��B�b��]�~�f1H��*�MqTJ�zэ�J�m[z�髗KRYom��Pt��?�iۚ���h�Q���UÏ���Z�h���p���Fu���d����4ɦE@��Y���r��M�R�z1���]��� ���U����Ջb�ɛ�����ÊF�l��n͋ú��e�U�m �]��eT�E����rZ��S.Ԉ�VM�&lQT��n�<���u�t "��6i��֮��%V���m��YpFJ`n�A`)lQ��Rj���,EF �v�����i;mn�p]���38^��WA�.�g\����$-��l�(RR`a1AB���P]����am���=���SN�E�i�"�Z�q�O�,*aW6Ne�/$[i3�����DEbV�#�A��w6�ZA2>����`M��7E+��-�I���x���A<f�O3{�|��Q[�v���8��yǸ2�:t���(w7V~CB٧Q	e��튁��MƑ8�h�2�x�JV+����
� 9Fl��V��K"K�D�ED���
j���Qr�,u�18�N2`7�Aa*��5R�d6��'c֕X��6�AQUN�
(��Èޜ�kFZ�[f\@n�k�f���wa��ӻhޒvJ���7��Jj�x�ȷ�wJ��Hm[�L_�w&LW��R��&�t�U���E�vFM�s0����Q��ʉRe��f~��Y��j�� _L��v�X^Z��![GB[*�.��Ȣ�.��Z�t�4#1�A�h	M��BR�U�
hU�h�f	 *��8��6Ҍ�8M�R�����"ʐ"�t],r�c*P�ؕ�Kn����˪t�ըm�%<�[(į/�2��蓕�b.����RTsPj��ⱙY��� I��L���6n�5��F=�2����qCWy�8.�9b�)����HTN"�/�Z�`+����^f�+���ej��un�uu�0�v�eĩ.�c����Sf�N^���,9�b�k���zo�"�d���j����E��SVP5WR��lV�c��s0����H�*�`���\U����M����[u�����mbU.6u�y�1۬�(����Q�+3C(�b*Bv�w+]杼:��&�QJ�F��f�K[�4����nǭa�$�f��te p�Z��Rd�Z����zv��J^��+sB���H�ڙ{1�N�0[���n���1,*��דC�E%�УKc7FI����:���嚎�w�7�-�l�bs��-���s!��i�����qm!�C���x������s��E�7�6�Z1�5�kKZ�5kf��D�+��2&���l����n�#�W0��a@��B����bE�Ƚw�� bDd�������;&��[��P4�{SI:��U�:��@Ӫ�l�$:��Ct����
J[��	&�&�Hj܃r���cKV詉⟶Zh�qj�gc%˶�sTf�Yb��L<��t!�n2j�L_Ң�x�p��)%"P`+�F����	ދnҷQ�d�a��-V~����HC������h��r�b�oN�w�yC�s���ea6��WF�^��]-iV�˚?a4��v�<�R��ѦK��)�63[.� ��-�G�3@�fX����:(mAea
�n�n~7���,��y��3u ��{ev��7Ku�;v��v��S6�,q���)fM; M
(;u���.V��"v�@��[��&f��/IM������Rm��`l��G#i�fX�b�yi�r^b�m�M����[�7P��C$'%f�ǲ2*2'��f��fYGn�S[�4]��⭥��텡Һ�ʻ�VVQ�1@w)�##m]��.^;�&c,��U���߄�4�dC_MXJ�ew�mRm���lڂ�г��o1EX�Ë%E��oB��hc��(�N�e�,��{z����xX�P��]-P�"�8tH,*T3Ch����¬R�n���U{s�A:6�v�P�l�������7!t�^�GD�EXVV"e�л���E��f��.�˫�&L#&�\��v�(��B�� j^-wK-�b��/6�8��V]�V-�W`�gZÐZ
"**8Cf��x�*��ڂ)R��,Ǌ��I{@ڬ��Ÿ�:��|�3y����/v��4J�;s���V"0Y���b�IUJ�Jj���S)�dU��@b,`�UA�I
R���!L)
IT���A���{�m��;���8��)3I���@)�vJ��/!��;�	�4P��&h�F�d����!Ґ��4�l�yJ�vb�r���V�kzX&��֣V�����c��e�ݦ�m�N�&cI^���j�v��D茋U������h��&ѻY�0���жr3���w&I3�4ʺz�f(�(�.�)F�S�{�[�{ �lӳ	0Cۻ[�E�!�)H��+sZ��3S�éiC^��PQ��bb���-<"� �V]�j��5���7&�6���r�ee,���lX�'E�mݵwr���CC1�	���BU����E
��]ք���
��$n�w��x��ǐ�\�u'%��K V"n��*�S�f�O.�0R��^m(<�����C��౩nfK
�����L�:n M�k̴aY�[c2a7*�g�7u�6X��0ۻ܋�NG������"@�M�&��X*�u��J2�eC�ɫLf��{X��V��#��J��a�'�naɖ+Na��b&ۥz!��HXP�t�J�m���e�PF~E���6�U�9��dJ�x��Yz(�[��/0[8�̱�0-�
����!	"��Y�75@�bW�SS]�r�D[*be�W��-�7p��m�V�Da%�הl:o-
˭�'Gp��hӠ�Me�M$�4Р���ţB���c[M��ƶ�GX�`�H��;Â�2��K�GQ��������0�
�	�YK(@�5�&��/\�xh˫�z���T�J%S�
�w[�+V���ub�ݹ%�&�� �w��%���Ve:����xU���I�[���B2�i0T]��B�0�V�
��\M�Z�Iҵm츖l�sq-
�%+I)�@���v�_9�=�y�֫}9fӐ��!���o��k��Y�[�)(�l�Ѭ���͜��\�k��Ry��EQ%w���R8fn��ۙP���^���{+�b�)X�왦:v�V03q��RV�.���0�=�e�N�%qb�N2�' .K�e�f���C�0/0��PӖ-�ZE��)~{�{��ԉ�2��4�HLlh1��k�w�Vs\{ޔ�aс�G�!z�R%�HbC��TVj�HUR�=e
ƪ�&4�N!B&�q4�@6��!I�bu� �/��T�����̻���+�nN�wl͈Zb��yhXlY�ڔ�*� �YQkD:�%)�cej;�������(tӽs�7��q��B�)$�L�\q���P��_w�����&i�w�	ÏjM2�l,0(�6IB��c�*j���]0m|�.�rl����M)t��#Tl%p�Cb��2tf��t��0��*�o*���#)�5ʔ#Vh�F@&�?��Ҁ�6E�+2T�$�܏���It��/7kh�=����o`xB�a�n�+kE�p�i�F'uv"ey*ӭ�Q#{��Õ�óx.�*VE�ܩeb�6���#^�;�}d���Zv�f�и�Bֱ������e7RakQ����gnR���6�el�(�y��
ͬ�u�U��Y�փ��O+!a�􈃕t��Q �n���̐���v���t�,h���,;��v=P�p���jⵙm���]e�+FY�{���L�68�w��9��ڽ
�`ł��×m�w*T F6�)F�J�R�1�� .��Y�`on�H����T�Pn+$ʰ�
,�]
�r�5J���)�$;�H�0�t�UP��92\02b�8!�c���c�䩵(�*�I���he^]�j�X��ejY�0��Jˌ�%�o���^d����ܕ��~b��QV��]IR�%�OAj�5S	�����ˢd6�fE��D���R���Kot����%��Z��*b��U���,چV�m���O��d�-��B1K5u��FȒTb�,�o/]��i���JX�.�RnX��7os%h����kS/\�kz���m//q�ú^(�7X� 0�&���B�M�v�U�2�h�źv��Ê	w�q`k��б�d֜��9`,�-rB�k,�
��*"���;��􃻌�nn��-W�9$�VSز��l)�㈷BKy%`�m��9���o*�M!AERIIH��)B�Kd�d�(0H�H��f�y��g;�xuZ֎R!dq�*���TȫLi[�,� :���+i�bׯ)�ůk%�$q�0�-��ҳx:�ӎ�M�q�5_�#�:a�e����0�o.Ղ�O� జѴnh,���S3u��n��W��XU��:2�Ѻ($��ʈ�fDvD�J�,��=gE�Swfս݋v�&]�9�Մe�����?f��Fb�
u�����`<x�c���\���
�3-�6Q)���_|b��,�����~k�x`����u���-`@'fܻ��z���l�L�t ��R�E�kD� �-̨r��
f�X겁��#.f�*E��"nB��8�H�O/&���+�r��Ȋ�Y�F�� �
V!���<�^��V�,�N�y5��a6��d,�V[����t��ڍ���z�e��,��$�+2V���%�K��B�P
�2E�X�*P�~��i�neL�+kA�,����� ��c�B��֤�u���4r�62���.�:��~��ܶ��i �-F�	���Z��n9X,��:��^8�䖝���-�:@h;.�6wpK���\��H�v�)���[�a�r��ʍ��sY��.��X����)��p�FR��CU'? t���/&iK��g.�dS�	�t(ێ�@��Q&[�����Lb�t�ǍȎ
�j��Q�eܫr𽙗M�åmy�-�2�	�sj.� É��¾���:k#܋J���&�]Dг�ޚ[/Xԁ�)��/o2�҅fJ;��̌�$b��کc�՘!���J���^����F�� y�@�k6kmԧC&f:;�h�L��j�Tfԭ�ld�p�TӃl
ˑ����b�����ۙ�����и�(��J��x����[v����2k��z��������)�B�f]��3.�T�f�����K��\��`~�13J�JS��?A���;��5�!�D���K�n���դ]U%��7
�y��n�j*���é:����2��u��K�ڱ�u�T҇H��M<��6gK���Uy�u{����]��I8Ȥ{�4n��5��w/{l�Lah���n�����NR�!��`ԩ3����
qt��lS��6�wyB���,%���G(��Lc*h��\J,��2�bXo
ĶIox�G��7�6wT���ja65q ʽ�l9Pe'�՘?md;�1N�]b�(i�di����0�T{��Ɖ�����N���)4^���f�݆���a%I#p!#���$S��V՜�	��]�6��"�嶘f�"ĺ�#������ �*���Eb�:����C�7r�ˉ��{N�@��8��&ح@&֯����B���YX2��LCR�խj��u�Jd��Ae����ڻB�Z;��[{�k(ۋ{�2Ƌ�7��N۲�f�����Su[�˘BE�����/(Yrj���S�:+Ph��q�m[�b������Y�D���fj-�e�Q��JW*0K
��#G-�"�6�&���ȉ���YKESU�Ux���N�!G��*���;�4�$e�0��S�5� �nM�h87.Q���xUDw\Z��h&5u*�zB�P���De�37*K��CkA/-7r)v+tX�n���W[R��F� =?�BnAL��[P�Ub�)�J�kc0�҆$ͥ�[�����g9��z����8��`}���fk/��W�4_�	�W3���s0��D�a.�
Rղ	B���I
L��Ybm�_Q��Ó��
�����㫠�YnA7@E�۵�SʉML�L�*S�s)[k1A0���Ea�CZ��^�p��m7�����!Kl�!�`��n)�e[�H˦]b�+��u��;�f��*k�mudm/�{��lm2�Ѭ���5Vt��J|F�7d�J^J���3�;����κ��YF�o~���YJ*�+S�/�vS�S���Z]컣*Nz��W�T��i�����j��so���u��.��X�vJx�1��b�{�^���{{���.���L��M]v�_b��gS[I�ޓ�:X��᠎p:6�;��npYOZe�v��Q�;�5�������� ��wJ2���D�3Ӧ5`�i��Wf^�V!\�V4W6X��oo�D*���A^V�ө��l����y��"b�0\t�NF�RT��F$�-��U�����W�[R��
���0	=\	=�ո�ͳy5���Z26���t`�;]�e��+��m�R�ϯ/)Z�t�C��Yc�A`���+�!+z�Ndฦ��L�*i�FQ"%�M�2�F��t�7�,�nҙ�e�@��2P�e�G([���l��o(ܭ�ˮH��	.j(a(�U�Q�M�i��0�!���v!�S;n����:6��fg"M#v����L�Ƴ����� �hF����Ucf�P2vXr���w)m��b��i��  c'H�oD[��5�hhT\7���tw2�4%e�8����mJF����්
'�.��ND��7���f�o���f�ؠ��#��r���^���%/�ryvss&�6�(��ƙUV.�	�u=�M���ڲ� �KG&�ǏtY�����/7e�5bv�%a;��x�4�j.��
d��Mţ`ݼTę����JA`�{�Y�.��s�R���҄Y�	9R!YL�ݹ�.�t��l�_���퇄��)�XFZ�YK%�F�_hD�Rݓyj��Ư�j�Ļ�fp���P�ƪ�+#c0��'
r�*I��.��Z�R�T�{3�VCٶt�W�\0�oM�or�}��Y�����G%u|Q[�bxj�g��\N��VWgAy�.s�����ؔ���&T[B+��^��J9�cV �͝aq�ԭ_E�8��ȷp3߶��E���bLإ����TBu�.�?�/��ý{A�ޚ��+�c��0)e�I�ػ�_\�$b�\]ǵ��'5X���P[N��r�A7���f��]� �.����&�p��E�V"�\��v���N�s���]m�"-Ɇ�]r۔�����F����j���Z�U*)	;� 65��t�f��Y�]C�K�o����ެ�Ws��F�vS������FB�Ī��T~�0�h\Ո����n�ݺe(�l�3 tiQJn�3s���k��MC�Ε�n\�NA�=�s���W�Ǉ�_^��.5�-�+�ݾy�u�zp���D���:�5r��U�̩��o9�=@�`���W8�~�2&�e���Y���x0�P麉V�����rS@��扽�Ι�lڳw;���9hph度��{�Opk\q�K�25��!��
r3֝���H�Zt�/!V1�h��36�`�w�U'����⺻�H�V�����H�)g.���륻;�e�B�4���4Z�����ݗ��<��սX7�w-L=Uw�5.��$u)&�*�ص��=��N<�VM`v� �)]���O(:]W���0�4��1��6�]`�s
�/x�Z\���SC�g!n�a��mu��W��|�Ɖ
p��ح�߆��/s�'�R/5�ӌ�=]׉�+�7kF���*�g3/��Jƶ�y���6�ӛ v]�=:o-���ѱ�E�v	f�E�˄<��rr8��/7H��sN%�(�cV/���ܻxi�m��ا�s�[gD��[� .aк�q���/6�P�ز� ����cⶲ�慨R���䯪�v�u����[�����C78�M�!�G��G�*�3��+9X�^�̼�x~K�_��^�4�	�9����w\�%F�a�F��40iՕEL)��Y���d��Q�9��nM`��s�w��6���1���)哸e��y�q]�����tr`!n7�������vۂ!F�f���թ�N�M��G���5�nH�r�S���;/�k,dC'%��A�R�=�98L���p �X��`��Q��7�U�;}3��[�vq��-�u�_ ��_>Z]=�Q`G��o9' ۺ�Y�,�Vj㝙�D�Y�9E���������eД�`a��eK�����uZZ̚e�����.�fv�I���y�f���0]��"�:�@�u�W����tW�&M)�&uzi����]&%��U�n�QQ�ЁuĀ�j{W�*U���H��p�3��y8�=t�H�3[����2���ǿ_��$�;��D�����z�3X� �#��']�^.w��pͭ�;.��j`&%k	�W���7FV�\�r��|ֱE+�2��f�p�u�u�*���e���;d�ػ2�w�0F�]��7�HJ��QT\��yo�N�Wx��)g��umIIR׹��fP����.3�%,���T�_lU���9Վ���\����+Ȋ�S��Wu5�d���d���}������vM��h�4NE;l�	����nR��;�qѽV�� G�N0���ԫ��S���4v�����'mC0��	�%�ś��^T@���M�y5}��Q޳�2J��K޵!�ډ��	2ڄ��ƞ7-aN >�5
ʗ�6�3����c]�\t��R�nMmo@K��� s��`����(-pN�cކp�x��5��/؂����w���=8Mnr�ݙ�b��Oi�d8�m�*�� e����5m�w�lS߉U��x�Ƙ,-�i���4X�s����{pc7Է�)�f�p��(�Q��e�w��	�DI��:�#94�C����V[��*�f-Ô�+m�G�l�Ty��	�r��$vfq�X�E�h���b����H9�n3R(�gv��M^������O���M���8�a��B��&'1�'��%Sƨj����ؘ�U�˾�������*"�1+�(�P~�$�� Hn\ڝw��z�й	.K�}Y�?]�'l#�`x
t��m�n������{���萷��T(��B�$�r�垥��E�hT��	��B>6�t�5�嫣��gk����/�[.�b�{n�~[R�s�]�^�be�n�fBs/�����tr�����P��*CRr�G6^�Ԗ`���IN<���de!&�*��X����c^TRX�
79jV+�oW���
ȨV�.�@�̡��N��4��e�#%�P��璸C�4�ޟ�/7��b�fV���,�o��ǡ�l��뼹�*&�Uy}�9fh�ը�"a�fJA��CڭS���(�1T�GV�f�f�mKƸ��G��Ke޳�Aww�1�.�j��u�54I9=�V�ܷ����#t�.;���R��{�-Z�O��҆`k����괘�Mm[�_�1y���t�(>��_
��y[�{.�âmcɧ#�X{s��Z�ZEi:���f���)�궳x^8�|
�#����M��˲G�S���Ǔot|�Ci��bƽ)�qwh�7�R��l˕�.���:��#[�&~�nث瀽�x[|�b*}�m)2<��⃓yY�̫�����ʧ-OF�њ�fV �-�+v�P�.oƹ�ڗ�ԇ:�TjjBwVb;�]���Xt\���.�g%��I���p۩���\���]���W<єT6)91&�p^���	�ɦ�v�*��qc7:j����Xi���Zٸ�}���t�f2�z�כI��u���ų]2ll�.~٬(@�ݛ�m��[:�����)�T�����S9f��L5��P,+��j]\��� f���X��G�P9r��KXSf��&�8�|�r����yd��Wq��^�ú��sGY7@�VKˣ���9��>p��e���2���1��*��6���~��·*6�v�]J�N��uo9ض]� �8��.�3U�W�t;Bd��z�E�bdή7�,���+:q�n���L��.��K
�%#�ڮ��-�ϩ�R�I{�%��A�i�/	i��(��Et��f+�u�N�^�����t��T�;F��u��]ot�&J,'��H�v��8�/�O����&���<�¦���V�of43*�1��c�{����|�W��_����3.�SE1�)�&�w�tn��=�z��xb�����+����a�N�qǴ��5ۏ�f���{��C[u5��{����p��Ҭ��[K7�÷8�q���q��H�*���y���.f�n� �иhSM�Z��lX�}C�s�S"�E���X���]�
��`V�Zu�"�-v�W�H�5�^~����
�]v�*���j��Tq���Q�f�<�6�(�B�qmJE[��SӴ��jnSa'7K��u�g�s�A�9crsW|.�<]$�.]���f@ޚl�u$��_]�k8v�oO�h_gP!��C3T��'��v弩6�j���
�SsF6+G<;|1t��{��n�	u9PW0��WM��ux���X�"�&v!S�������s�<k��=��C�t�䔖�Eɔ�r����X�_��{�:a�g��k��c�]ڲ��ֳ���3)���x,T�o&i�Hp�IvFb\�vA��{1�f�b�Z7p�B�� c�JP�K���yW`}�����aǩ�h��_7 �[�;��oJ	R���'����ﱋ�9�N�]s�[5�����$�7:�ި������ �Y�����e¸�t�N�����aB8���w��&�x(]:�Y�>�����j@�m,�:����7|'�J�r;Z��Z�_�C#����X:7\5W(�J��c"]'7�UeQ_֥�0�i�S,v�S�^}�腚�e�O�v�@��	 �r,��឵�=N"e�aj��]n բ�������s�
\͛.ͅ�NgL5����unΰy4w7&�s�Z��MFP�^�r�
Lȭ����D�., ���.��wq�,��%NF�Jُ6l��+y��o��-m�Yos��#�sz��`��'���Eu3��F~k�5R�usb�,���VwH���:t�����ӫʱ�q������{Qjy�Qsn�s�#����ƺ��s"w��.�٬���oL��O��%���f�}�r)�5^�-�a�vi��7���u���j��+u*�buʲ�:a���Zk��Y9j�fwU��fU�,����{�*�]cl��n\堾;���ǥe�V;���af�F��]CN;2dظ,Q��N:|�:]�Ǔ�k�q���2B�X���r��ͩf��Óv���]�b���W�����d����������:����QI�eo�C0<}�p�S�k���'sx Ghef����L����g4��G���b�Sס� (��Y����p�O
�Wq!oU�BC�v�m|�оw��,�2K�e����H��E+؎Z�<c J���t����]E�5̸����B��e`B'*����- �C]WF�WIL��xi�L��\����ѹڎ�|��pɪK�����K"�U���d��������#7Z����)\�b��m�8��oZ����ۥ;`6����wd� 8U�3j�pfc�$L��XۜcmӼ�p|:�lP�{6ƽq���U�ő��ϼ���s%��4��\���q��Q�5����ahG�y�ft��m����y?(nB��W���fvl��.a�w&��Cl5հ���r`9{�w8Wxa;:fU͊.f��[��Ty�eh=��5�Z�	W;M���՗
ZΗ��'�Q�u�yug���)�t��Z6cwk���+��nL��Ɠ���F�l^v๔���t9���)�}�X��h���Idj��(�Y�ͫ�㸸�=�69�&Pn�kp�u��YN�f,i؟_e��-<R�:v���)%�]���B�ً.��B�r��Y���㜨֌G 
h<t;�Aj�ř�7�E-S�
�7��9��`L���9�sy���J�bh�U�&o0��7u-X6��6��)jfdd�P�+�;��B�rH<��6��@N���x�J�6��	L�c���	���ݭ����8s�u��M�V&:{3��Fb�������s��~�A��V*���n��[yw���Ҁ"�i�n�Y�Y8��ɻ���2�u�N�JcVR.����eH��Ȳ��\,�Ĥɍf9�C����`x���]w܍�+6��nU�����@�PYi�늬Wd�J{�f��!�8<:	R%N=:d�8�x%���V�#�����z�!)]�A��9 b��!�`9�!��������{"�V�ڑ�!Y`�M4�ғ8l�z���6U��Z6�څ�"��h��s�~��Db�L-�
�Ĩ��}W�8�wW<C�Δ9��T�`U�aZ	s��oGvGt�����q3ya��s��O����U��9�dn��ī��������pn��M(Te����s�}OE�Wu�ԩ%���v����������7V�SZ��|�.�3�R����|]ɮB����E,�K�Z�K�i��;(D�/��ۊ�����[���{[��`}J)ח�4s��\�ES���r
*�5��Ǫ[�~Պ����0)��=!e��I�#,�a����-wM��H���7���v��P��u�"륆�C|m�(��\�� �u��G��]�Kq�M�I����;(���0�!�{8n����$�<�Ŗ�t-\���O,g7W���%x*߶���.�md�2�dY�i���Z`�'��N����A��D.W�F���f��,Yy��D����:%V�k��[vu�E�6��j�깮K�d�����A�؃�5d�ӵ�tV6�]�q�[WlY0�<+7AKf���h�eեo �����Mj]��'�w�͗ZݬȺt���	�����ԵWV���1*;N�,P��ʺ�N[A�^3*✙%��5��HB:��쐒;�V�(_��YeBWVES�W�m����Rۈ�b�v$�d���߄��I���� ��C!�I����I�
d%0��H0 1$$ JI4��!wP
a�5- �@��!L�'R(N!�I�`S!!�-O$��8�$�)L�$d�P��b
���0�T�i$����� R`B��L@XS	��ީ2.��Ia
�Bq	�C:ɉ-!ĐB1�2��W(-�3U$-�CH��j�m�7� �d�j�Ih� c!��@�v�&2o�I�Q$���&���b��a!L
Z0XO$�I�1$���)�Y$����O �����m$�� HZH��M���PI�6���1��8�̆2N3�	��8��4�2IL
J@�IL� �8�� )�l!�%�AI$��S!-���
AI!��$���i��Nn��S RI3�2u	2�L!��<�3;rKB������@���I!L4$��L)��<��'7P��q���!L%2DNC������'Y-$�m�`K�,���A@-�6��Pq'�"���B�$�!��M$"��@���Af�Ja8�4˺�L��@�I�`q`�ͤ	�uR���BL`�T��<��m$�aޔd)�6��d&$�HBy�<�$����)����Cl ���BHk��Dn�m�d\�Hu�%�j�r��g*CI����u�b�&2A�-�RS$-�(HLI1��I�C'�!۩"����f1B`�- ����-�KF褀S Đ��d8��VPM��!*�$�4��$6�Će@�q aII
�Xٶ��� �1	)��, � [I��Ij�l��Q�wP8ͱ�q��i4��$;���HS'�m��7u �����$���U	�՝@��$%�C̒�gY�w\�m�;ۓL�Hs(9U$:�תm����2��7P=�%�8�Y�vbH[:�2lLO$����m�RAd�i ,��}@t�y�%z����`R�)��*�9�e���QaL��0�z��%��M��8�Ho
��3i6�t��-�i�L:��Ka�q4��ՒVP)���H�)�Pq���&��БKd�u��E��-o�0�R
���-�JAHV��m�e�M��*M�,4�ߓy��r���Ja��j�r�����q�(a1&&в��}��0�ئ0�e�n�&"�y���9Eѕ�Ćө�xd�E��C]�I�
��1���g.���;o�<�I�bbw
�C�ˤ)'RNv�f��j�<�C������v���iyD�W4i�Q�����Wh�^�wwhc����i<�m���Bp�\�;B��n��*b�f��J�u�Y�4�-������S|���J|�}vLN'IJ!�#�""Ub0}��D7N�#,vU��q��D��1T.*KMv�]����8�C|�ӽi�k�ft��oB����i5&���" �B��7��_k�QY��!38m�J���_\��"Y�����x���D:�T�ZM��L�2�ն�L$E)Q���C�eQ@�j��Ŵ��r�@�+H7nL8P\71%�D0�f���8�Z3a��5�z�����V:KU�XU��Z�$�zfd�"�u����әW�3UcX�rW\�.�� ���fnV�9*�ln��M\��z�{E�5�s�0+�tR��]�w�n	i10��L�+9_@�bT�kUnV����4�]�x�d�ح�kzHq��&�'n��-R!���J�VV��x��-�a@���na;R�2N��,i��@���T�sz�Z�O�LYI�:�|�B��*�O4pep5�����AP����\7�d%u�9?n��eu��X\|(��tގGô�WS(*
�	x%M�0��p�y6�]�b���K�E�`�*/�!�"�%$366KĐ��nf���qJw���P(���+���?���ر�!ʗwwA�,�Ã(�4�5��c���Z+ilJ�,���9�+ 0�f*�7PAcK��  O��
�-���M�1�b���R%�:e�_H��6D�A��û[�9j�b�|��Kz�WO"�B���S[wS8p1Ee�I � *�n�����W��\�����v�-�9y����H���lii6�bI6�ہf�X2�˲�ʠ�B�]�qՌ��j��6��֐����*S�m�p�[���
�T!/.C���e�)V�nحf����_��[[I�֘ʰ�M��W[0�eէ6�\�����r��eY�j�ҽ��Yt7jXd�0鄯NSY6XIQm����jC�c���hk�P�r���kt^�R�X	dcf=���h:��h�j�|;�IM~����=��暺yv��fν���˖еۘ.�J�C�7L,�5V�[�s,3�oF�ͻ���W��v9d��w��r��Y���hE��yp���`ɜt�� �>��.@�I�4Z�u��n��*���`j�9:u���co5m6�ܻGy�yB@N�l㶳�*�Ћ*V��W�4�6t�}��y6���&Ӥ���*��j�j�8�LgjJ�@�೷^���u�����YմEH�2�c�Վ��cJ�lV�6�S�]#]��A�Y1w+��):
o̡-m�
�<i�\6p�,:k$hٷ�{p�|���)��=�֖�6����+�G0^�b���뻶K��Gpt��Vu��$+����pM���7R�4��:�{Jq�*+��b���h�X�p̊��u��.�Vr�s������Aк��;�ޑJ�z����l���1С��񵕭Ω�*ʗ�$�P�5zo�&,�/��J�mvK��ܕwL�w:�t�3\xJ��6/�X�a�׽���D������s�MC��8�9��kmUB�n���Ñ[)�E'k9�F5Ҡx���H����!��r��;7��Il�Fﴫ1�O����
�B�LY�:Hf�se+��D����4�m�|����P� �<r�~��;
�1�u-r�W��(	l�D7p.��P���%�f��
�̼�Ȏ��#��<��7`���(���˭���W�����ɍ:�rb55-�HH��5�����51%���M�3��=X�j��*|^L�7��굌U&4��;�������1��[�Ӽ��0��pG���_����L��O>��z.��	�y	�\�А4�����I'B2 9��:�	�H�!y�i߹��� �B�$-�	��$稒�y�����I!�y���ܶ`�Z�;ϳ�����{|����_}� �1b�Db���DTPT`�H*0QTXZR"���ʼ���AH�*>�F�DQQEUTQ"����eJU��FAb��d
�����*�E���2ҕ��,X��־�H�DAb������U���R�E|Ќ40S�WTQb��"��#b�DUc�L�EDR#�����j+�H���,Q��V"�4����X(��AH�YD�����H�TDPPU���"��XK"�QUTc�TAb�`�R�TAGVw&b��
�J`���X�,D`�UE ��\nਊRPТ�UN�I�X

�PT�
+�)�z���q���g��׳���zz��v}�L�(���*a���ڥ�U(�DfT�Uz��`��(��E��b��.��"�"Eb/��B��Agj��=x�AE�"�AAEE*���}븱PQEX���J�"��(.刢*)�AVV0�%�AV(��b���E��^�+UB�TD�P� ��uU�w~�DiDUQ�_UF*"�u�wE&�]4��U
��T^��������u��5߳~�o��Z����
��n��TL�d�PF6��TTQEDU/TZ"
�AA���\�3��QO�b,V(���j�D~޹��V��Jb(��F�fDDT��:iES5Q�h���AdNԔE�,�I��z1)��*��D]P[h'R��;*R�����,-TM4��fT�ꢪ���QU�Wy��[��W��Y�|���{��5�����uK	m(���bV�dH�(�T���@QD5����v�"��D������Xŗ\m"ǝ��*,�X�Sm�:Ԃ�X�>J��{�֔(*˪ԥPEY�*Z��jQUUF<����(��ԥ����dEM�ꥏ̥PPP�o���uT;xfz������7�)/�%�H0Uu���QuT�jj�(�1�Y����$���a�sX\c�M�
��Ҟ����TPU^��(�SU�(������uH5��b���DE����s����PD��k9�O�������/��Ş���@	(�����{0e[�Q�"�ʱTUQ�JR5F�S*���P��OYCv�()^{�b��um�QC�|f.�QV�g�?4AyUb�(���W���C�S415���*�Q�F*��g�(c4�!ƅ��w���]*���}�v���h<u�:�\kw�&/�� ��̺X�z����iHj�b�Ĥi
Vgk�J�21QM�/;�h`��!ĭ�]�\Q��5Mv�(����Ҫ�PDo]c��
QG�<]�H*,U�嘢J�fz�l��Z�������ݮ��\���>��ϊD�(TG̤k>��GM��G�E��x�AX��D~e*;q-k�w�QDYꪢ���g/�#T�YF��4h^�	�j��Z�R1�`�҅����v!�ya��Y� |�����d�[�z'�����z�{�����`�s~�;ö���k�S��b��v�}r����m)�1EU_]�����Sw+�Qm��b���\��e2�U��4Pi�.�J��b��S����wZb1��8��.��K�V��k;]m�[pBˮ�*j+.�Gu��������#F 3u��/��eO-�ؐΝ�;��oqzS��WJaǢ)l��}c�����L`�"2�NL&��y*�;��`��Eo]�}��OX_�b���]�Y��`<�k7W��������;J�v�`u4u)�Q��j�(��z���딊�)��_�Q���B�j��x�hSe���t�f����;t*�%��h�\����Bm�&*"�oW�j�(+U�����j�7��?w�����P���:���>Jz�"���9�)>J{E+�L���>x��0�S:��A�s49Y~�R�����+f�U���G�V�v��T���"�F*l�e"��N�00E�����t����ۮߏ������g{��,q)bS��}կ�������'�v���fLi>�"���w[����y_a�r�E<��(b(�ƹA��W��UO5�	Ƒ�ձ��#M|��WϬڳ�PD��Q����9�r}Z�]�����>�y��:���q�'��N�(�}�4>gQ��}�Z(���Sɤc��ު�U�UE�����SHu�W׻�
�*<;R����QQsUL��R������k>��Z�ds�U��@�@� d>݁k��Q4�,�
�}\������P}t��7�D7�[ڦ=�ֵ���Gꨏ���h.��W���7����B�X�����q��i-'��s�ɨ3IKEP�E�ڕ�U��ѳu,.��cn�i����0|�`�<�u��4�L�_5J�>���6��y�"eq-���K>~��}�ȱ�p�*-��״�s��h}T���;�W_6���wy�{�w
��U^�kt[@mo�|�p�A�J#�U_],~�ڜ(��>���J#^�F�WCAT>����ꩭ�}E(�ܻ8�5E
*��M0�5��
G�_h��eD�W)v��o[�qيZ��k�MC�����GùD(
Sˇu��Ĥ�jꪕ��]Ρ�m�˺K�La���ob�U���q5�%�;���kf���uB �^��i3��,QuT��{�{���=u�w�wz�g��>EQ5R��aI�(�O�E��O�G}�3���V�Ui`���U���s���բ��*�{v`��C�l�ﳾ;y�x�" & B6��(G�W;��51��$���7[�+8��?���?AP|]m�BՈ}EG+�~��T/�Q�[h�)S�B��Wj�Rz��5�uE �kWZ�E�Ϛ�i,���λ��"� ���|MF'	�wE�;`��<�|�P�-�R}ہͯH�_b��c���配fԌs[-�b�`Z�4C���oJ��]]<4����Q�W��m&}N��E�('g!�.,��ŭv����Ž��RͽWG�9�i\�������D�p�&���������;w�r�E#�)��)��P��Z�EO��)h�U2�L���1N4&Җ)��PZ���v��(uڵ����T<;�k0DE��[љQ �hu>%�6��U�إ�	<o]����������|q\Et��Hi�
\��p�QC�<�S���z�#u�l�S������B��`|1h��77.N����,�9~�4��?�@_=s���a���2���|%Gu�s�4��,���Vb1]��g7��Gee޷���絣��B�+_}���](��V�g͉��D!�ᇛ�+�i��9R(�.��_	�q�Ɖ���r��٬�U(E�Y��U�,N2��ę�u�}Y��E�;f
*�~�SNh�]5gs?R����`�5����lM]N���w�)��ύf����4h��1E>ʱ�}k3�V5֪���D������l�O�� q G���?�
�<�㝃��G��N��޻H��߷�ot&�_V���"���}�G�.J�AFQA[��� j0������4�z�To�kUB��쎠A�ps����N��鸠���w�Z�@���#�W7��#�O�LH:Q̦��=��W�����l�Ns���1�g/:a��-�]�/�V 0�.���Xa.F,&ԫ酌
�_�:�;}��5G��g���×W��(<ʆu"L( �F���Y��J�2��;y��8�7]��B�Uܩ�)Wpu^;����4�7���·%����>`�ٚEh���P�ǉO~��P��s !чj�D|����+�F�3��E���҇Z�L�U
�����TNVʑ۬k�j�͡1�8V(B�D�\N�0��#G(N�sI��z�����St�U>f�S�(���k�G�g�#�ӐtH�<� Nl��m}O[w׎wu֑bշ�rz4���w� �׵0��[v!ݩ�8n�
gr��ԥ������4MT 2�<�Zu��3��S�U.�Iy�&���P<!;�  ��ԃ:�]d�2�,s��.;X���U�)+r�HS�wDr��z�R��N�psK�ʫ��C���#���Hm��w�-A`BH��a]�Q?����m�]kE����DMv�嚘� }`��!�ڗfH�-vL�Z{�7��ek[�]Z8�TT�S�GuB0o�i�ࡳb>xKc�v��Q_c�b&Ҏd� �
�	�S�:��v��5��'ή�Y��CS�7rN��B���Q	�F<>�1@	$9Ն)��r���MU{����f2�z]��Q/�3Ο%9\��8�	�%�q�p��Twm"����x�F|VY��F��8;9�ϴn�U�sy��H"� 
6��j�7Cbi��7~��f�񲬳M��y|��y���wؑ<��'sK���<���?�^������+Z��4��Q�-u��b��#!�&%f,�(�#�d\�L�t�������j5�ˋ=a�V�����&�!��f���cBb�p#��|�'�������ϗ��Q�u˛3����hm>�K����� AF]]��j��g+�B��C9B�d/�8}r����ki�Z~^ѡX���K��VO��T�x� �!�f0�L�;�b`���lG
{YX�Wq �
]A#i�����hA�~;��  �:��!�4�. D$X.� Va�d�.-G�`�hk����Ui����׎=]�x����\0����s&���)q*'ر�I��L(kmuDU��*:c�ƕ>$�6]�S�AN3�;��{��]«�+}9��|�c6�mѥ�:��$�%}��D��a�&qa�YB߹�iUUR�fI��9m���M�{u;"���,�S�fz���~� D��I��YV�m��7�f���lW9D��o��e̷���k����ݐ��k���v���֫5+y��P�%��XZ�N�����N�Y�/�xɕ&����nhTT��t��5�|k,Zv�ͦD�g^�2<�P]�������w]��V8���L{B�!��!Y�z���4G�A\p�Nr�2�����JN�U�ۡ�Qw[}��Wf��z�7���Z�[��²��=�I��@G0#�������� F����~��pᆢ�ޙ���!�B�0�Q(����!�{�W'8{�Zy��]*̯W7��6S���ό7C�e�m�h/� �� :R���ռ{�kn�xC���v+𠰠Xa@� ���`#+na� ���x��zWk�6�F�-t!3$�T�.��� m�d̰����麾J��)p�x�]utբ� ��{SI�OrK|	
=�sj�� �3����ʖ��,W2��F3^���ӫk���f�V���՚O�׊�xm�� �ckr�`�1z�0 $�]o�������lZ�~�$�תlih��YN��359����b2xݞ�ɂ�����[:�1p��L��.f�q`�PȲF��C��z���Ҳ,C�]!	���G�s��� �"�L��w�. ��@���]L9��FSLE����u�F��sw\�" �LK_(��QT������b�ɥ]�!�>7u�0 i��H��������I�J8��K��y|4}����R��׍���9�h�0s�f����^+�d��9=tz�TN��/��s߃�6�T� }�3�(q!�w'I˩�׷:�o�^�_���^��5֕/��Ʝ��V��s����;�Y�vAW��P ����D�s @����T�Bq_AX���`i0�#��QP!9_n��҃xs�����y/oχ�U'��xڎ<�V��c�ި��}�D�n ��S$��_䄄�N�Ci1q���IL'Xy�tB�)��$� y�����^�[W��+ꄷhE ��+��X��ovI-�&Є��5rq��g���'yP������3�HN|}Up���'��;��Cl$�5 |�- �!�R�L�2C�|�m i'P��$�t _�kڬ��u��h;�q�D���z�vvK�]ۮҏB�c���F�l�:��iJ�[0�+��1(�b��V?:�6W��6�}S�)�s�M��-�--���)A/�ր��I���/�P� �|�g�Oտ�ڳjRf]]'[3����F���豐 K�G&a!����	?�ЦG��k@G᷉��p����B�ӭCeQf�����+uK�gu_s���5v�����>eP�y��))|I�~�#�L�x��F�C�s�;�6��=���U�q�����#1����9�ل���ff��+�B4l!q��I�Px؆�Q�0b��<!I��1�-Cި���&NJ>r�R�⹹.�b�x��A�C��M`_�;+v�s���� �n��/3f@��t��LӇfA��(�dF��� &w#C��?�Fmf�,o����`�\�E��#����D�>�m> q6���Z煩�P� ���hY�Ƙ��s]qd��DV��_e�)1	���{����7j� ���g���&�q�;�F'ɗBz�?O��c̣C0N�5�ej�7ty��P��y@�yG>��RW<b�TElX ^�&��~�Hv���S�+9L���#�:�0(A�H�\]=S0�sՀ˅G�$}��L��F���!>��e�a�z�gh������0#;Hp=�n[�Q�U"[E��^���5��:�Q?PPn����Ǔ FVC�zP�1���K�5Q���y�:�A���prb �L�+R6²�}d�?��![�:2��'����:Y��{Ac�S+�mR����:���m�~}�<��ޫ���B@)�h���� ���w�>���Y�䐝� @� oZ�_������ѝ�B�8�{��y��պ���\]��r:�U$$}�	�,��z�����Vw����	 [�I-����8��kw�f�����'�i�Wkn=�7���Vi�͝țu�Z�/�C&uK�̢ U�,���2�F��쳵�n)�j�YK�IY�M�N]u�[^Yܚ�k'L�:�\��$��X����Y�*X��&@ƃ�ץR�*љ��weG���]�2�E���ۈ�@�� ��)�����Q=3?)cZ"��@��ǹ���˱7bf���}8���i� B�>�����Y,��ZR3~��1q+�zـ,Q��SYnD�L�$��Pc�����5�g㐗�� P��8b� | �0���s��:��;>bć�w�B�6O�>��M�\���r��.lvwyz���B�pj�DxW�Q1�����H�Q�W�j��S}㘼h37�p�]PWٺʿ�--C.:�Ɋ�l�1Y5��%�����3��/�r�T�9��F%R�����z��sCY�1e4k�ۻ�_atr����Zǣ���;����}C4ﵭQiFv�wNG��q��5��q�c�؏`ۯH�u.J���T���*Fbp���2E�})E���U���	*J�w�b�T!1�K��'#;�xj$J3jZ-�P����R'9/��nfG�n�*!ق �j�U�U�<xq�;''��
�, ���M�V�����"�dQ���Qt5�e�����s��P�:k�<:U~+�u� D��G����9�Ww�.t�����/_�\Y�D@+̹�ˆ�5��¦�KJl��֢�&��m5\�QB�a� }��H��r�8F�W+N�1,�<���\�V�jť D�h$b.R]	G�˷��R`
:�L�?�^l�m<�f��T0C�����7���t�vr=L����3%S�� 3 �vC�g>����6�i�zQ{��`�����4�z�W�J"1��䨒��*���}��p��ȝ�����գ�L}�|�����)���b��ko&"!�K��1�C�?m�?���G՛�N�������wsﻭ��V(י��w��ި�/"�͓�s���^m5�t78 ۬���z�r������i䨛l�S�qu8�VZ���j�)��?�� 
�H��+���7��4�F�X�:��K��4��dZ�����0Y�E�<co�u\Qi= +}��aM �q���0)5F �o��'��{;��(�=||��s۳�%v�� ��l�C꨷�2���@s<��'gv�[u��0n���%��Ln������i-�]��)�t����kuO�t�O�=��3K۵�/�P�ø�78�V0��"+v>;�f�L�w�k�cC�h�ɦ;�ﲐ�ie�;7">p.�-0�5�6/��G����H 1IC�z(��ٜ���8t:��"�um���`�0p�Fs^M|�u��wC�׷���G^Cf��is_M�YV��j885 `���1�.�$(]5T�b��p�T����w|V�>�[��Z��f��>ӳWU��뼊��S��Z����Z��^���(�8�3`q�H��:�#2�L�z����w�<`l:s5#�G�`C�Q��U
��C�:pv�	���l�����t1�ࡂD�U��؅Ԡ	���dd�;�"ar��v���?D����
�L���/��h�@�1�i��[hy/^�һE6'�7���n��� ��֣�c(�������ڂ���	�����N;H>1b�����5^�&�*���J����%h75�棳�f� ��чb=�悅�UT��I������\{�l�L �9��1p���R�1>�o����sk�����b˷t�.�a�X!��t�#(���o3�����Z���|M	ԝ��(�Y�:ڇ<���zv���fz N�G�+��ο<�+�{���	v���ٓ�.��S�j�<D��eJ�WM�����G�����DcFj��J�ӀG����;u:�մ�{��S�3r���|N�����<�@�$��*"��@�͉�<�`J��uڹ�*޳�^�k��hA���H�� q1tP�%d�ML��n5����f�דr�_}B"��7tb����0�W�����NQ��,������G�DD�t�"�&�͆���O�0D[��~=k�a1Yc�V�O�&+�I��;�f&���d��za���f6K��X7�5ObO�3I��$�༣�sҐ1*�̶�n'�̗-z,}�R�D�<�"�01�U�@��\-�3�0P���6�� ����5P�����'Y��ٍ�
b�Fgw��
&�j�����m1�;�qb�7����׵F��=U8�C�(O��[�6l(q�`o8%¢�b��KU��r�o��;�@�۫SO�:���:,B*�\X��| �L"�ۏ�Ա�Y��^�R,����9��F�\n�7�w�݆��!@�b9BU�e)�X�&7-3� *c��(��,  �w)ÁBo���Ę5ɮ���}�b/���q�U
����	�0�$d�.���;q��z!$1<�0�ڊ\L�w4u�{����[��e?�૝88k��/R�վ�(�b�vO�O��-��]��c>���}x�]�90��o(YMz�]O^s�8�?oXa��k
`��F�De5�d���`z$ٓ�5�֚�[����/�y2��>�DM�¥�`XՊ	?B{�D6x��-(<�v���2�'����qM��PD\����9	�S�˧���t�WPъ��^L��b�u�3���4����'VؚN&R�s�V�`��c��ц��O�t����&HXz�����𫾱N�U��$�s%�����,��_i��R�i���ͼ�M�����Ʒ�G�+NW������nU<(�8�.pyEQ�uA���h 9*xM�`͐"�����nkaM�M9Y5��`��+� �p�^���'����9]������}���F��|�8��t����/����}�p���ڬ�LlA M53��8� `��37 +ɈRx�_0؜�ln�Ή�:��`���p���=�]�<��� ���#oO5��v�^R1BJo���C�F��iW��D��HE��vݨT����1Ad�ET���Ns\����|���u���Q�Ũ�e�&`�.24Ĉ�DVk�bs�D!2a�@�n���}0(��v�-�f�l�S2��^���Zșz��>5.>�,eF�J9�9��H�U.��H!���U�Ɲ� A8�m�rd�ENQ���b��r*�8���A����s�MGV�x�<$,�ڨ�@� ���]�  
��v��s�{p�H�^���u��QB����$p$7*&���`�
�\ʽ������#�b��S���n8�����RC΍�5�%��kf��#j�2>���`7\u����b
?�"�A�>G����H��o���b�JI�F�FS�t]��0Dv�����'�jTH6~$�����b6�?�ZhE����h|0���o��OЄ?^�y�*4��sb�:�זD@ķ'-�l;��	(E�ݽ�Uf���G.�eoY�`����bkZ��:f��9I2h�^���!�M[*�^���0�.�'J�����̾�������#�X������J���i�'G���`6�om����m4`n�:3~z��t �A[�C�y��,=�+=��z���)b���\I�A��_<�a��3T�n�̊�ZK�ȇZv��_C�1Y�h"w)���Y��x%mV�:�C��X읉�����3B�U��Oz�r#��~����mD�b�=7�/���l=O,�{\{��z����u�o��lǇ����y�-�m��$�54cy��-ڸ�߀����M�)WZnR�:���7����
��ޓoEi�E*��<Z��@�F��;�5;+�����ͫ8��C5�=vVS���BJ�\Xu�qe�S[j"_G�l�c*���Zu�w���7�7X(YO
S�˕)k�nR�@<U���B�sd5/���Iu�Q�7�J�W^�����ȫFfL�gpy�N3j�&�!�S��42vN��7�cȜi��v���f�Ǖ!�)A�w ���U�zP1�7S�x.5$�ܳ�ko`q��j��٪'� 
+]����}�q'6�6��Š���j=�x�����e7u��v�H�(wWa��ɂ�s*�8⃳"5j�8gdX��x��uh[���n�k/�5�/[�0��	�C�՝6�S:VQ[P �coѼn�q�rI�
IE��8
�jʗG=FgP�5�]C�7���h�����(N(ǌ]��y�� �?��d���(�N�sFQIICgg^�k�������3{GWN��	����]��ҡ,�N�	5��] U���#^�Ճ���b��vNo4�̈́�;�X�q5�^�2tO��4z��(�y�%_=�z?#��ٙ��\�&�ݮ��m3"�}��vE#�+��j�����o�`�R<:.����*h�1��⇇VL�`�u��e�R�;�\'�*�L�@��mY���t��{�\�\��� e�Y�sx�_13��l�AU�7���5X�NV���r��IO�	��)�Y��`A��3*�V�e,=fWv�u��n��v�gg�m\�2뭬꜒���O%w�v��k1�r[��8l���ݧs�.6{�FQֻ!��J��L'�����f-�}����qdRSlC.G����}�.�Z=%��J���`yÉi'Y�,
WƋ�x�6�g��n�Vn<ݱ�9� `����Kq��q�-d�I�z2%)�Wn�ҠxmW7B���[nX�ˏ;U!��N!.ݕ#~��>���}��4�D�U3^�]�'�]?�K|ojgqe���;.��o�KkV���­�uj��@J�O����S+b�_TQ�u�X:���P�� zg��աYu��<�}��]E���S^t��s �Ph���c��4?�F�������8}7=n��}(�B̬��hmn�o�y��׹�8C�P�k�s��NT��b'����0~�4�����J`	v��ʞ�+�Ue��`+���/��5-?5��g4{�wvM0��?�y�5!]����~�>0�*d��<ܺ�wC©�,q�V��Ex����9Q&�Vs"{3ܝ��_w��ڀTQ�rE��^^�"i/���ers�˞!_]�����u|���:4б���jb`|�)f�z�]����ew��P��z��vvjqC�n	�X��f:*A�Th�g�I. Wk޴�=��ۯ�9���xX�Z��˟�?x��B�UR���\��]G��m�G�MO>f}McS1�(ה�>%���j�z�Du�4~=u��h�,��u���g��l�'����c����@��>:���ę�
2>���TK�d?��8!������]�lmM?-�����$��+W
�"�O�[t�/�iA�x%ϡ�e%��>�L�^쫣#Y�F�����ϫ�'��S4f;�ﾅ�@(}�5w����,�@�X\���z�p���6:I�	UM�ڙ;y�0�ɠw�q��B<{�����^$�M
����N�����v.��c���%�w]Nk��lVe������F����*�Of*�׵]�;�tɨ�Q�՜��9�P�)8�*�S?xB
EQ.Tt����]d���Ga�*g���9�)���c-XuK�
��\�j�Q�&9)�P�YƎ��d�T���A?ofk��6��ò�j�,�[�#K*��M��oVAnko��͢�h�,�qn؄3��qU
�YX�'�ǃ�>IF�{�K�vUR�.8>������3�����'�=�KJ}� �� PDX.3���@�鸈��}���*)����|~��D�[r"KPeQ�}&DdF�\��$���Z.ε��v��<��r���]��<�
{����K�v�G1�cƍ����0 �2!2�)m9����uH=���O�vq�[/���DO42L�im�{hf�苉��%�d�`��;	��y>V:�G���͋���in�6&��!�[����w5ה���Ş0�P{L�>�(5�a����r�$A�~^Qd�����,�q�m������.��<ao&��V9A
�~��ld,�*`��0P���Q��P}C�輌>�
P3^��q)yڇ^��R�{�6��A���0/�F�'�| ���?� ��� ���t �,p����]ЀLVܻ��"B D�� iK�_+z�\�T�z�����TfUG�툽�ŏ�+q�\x�a&ڇ���>a��ME\xD�{�j6=���&e]��'/hdv�׾O<�0�5r�#*��^�-{9P≤~��*m��`l(��{��D ���yJ��G"��J������4�Ͱ�>[���p�����5]g���{���D��D�y�H�;�N%/1GS��)D۪����nI�$.Tj���
�;NM0+o�������Ĥ�ׅ�?��|�>#�eM�w��
��#3��0��T��&*���h
D}`�B�l����#Ew�d�5T��W��Ƽ�j_w�f��U��_)[����oy��Ů���sv��]��ٺ�/:h��f���9i��D�X5�L���!������NK׷��U,3�v�����RΣ�Cj֫`'l��7�o��&FFf�Fv����T�֪)��u�C���n�����?�l���#��2˘/�6��Ɍ���Gvg]G�K���6�ͰB&.�Y���/.�Q ��O�uP�y����;��=�6�n�Z4D�#����c�B�~��`�"	�<��ذ�<�̓i
u��!�yȊ��)�g�"尣�9U�~�P��^�B?�8!�/Xs�,����U~̅&*�L�0�CLbQ�ǭC�e�_I@�r�����O��e!P��b#W��%�`+Ɯ#�	'��kt���0D�"����Ş�"�$�V���B%n���Gfv�c
|�B _Z�mɅ�2o��f��E���w邥м�г�H�I�8bAq5�)?S�W$�sO*.(E���LI=O@wrm��Eۺ�D*��7�^��*� �ȥ,Fj�Ó��WI���f���+}=ܾY�$B�n��6r�o|U�L�1?#Prj�b#5�Om'&+(��C�z�S7Yٳ �i�v�_X�(_?_M(�����u�#�bDT�o2Ǯ$^F�s�!3D��>���N?=�/����	�)-ej��il�aPe���1�d��x�l=�lZ�+��^;�ݛ�ƍ.�<Mh��-�SCh�{�����E����'1}�y0.$D��Wx�ˈɬ��U%G��=�t1��
��!�ItJ��Y;�B,������2$F��
��k��y��#a�h%^C$)͗7{,��ύ���F7�t�ClO��f7F�ЃϪ����!	Ǚ���"�D��@��GEȁ��*Xʥ?V�cҟw��r���݀���GX4O�֮���9��0�����P���k�ٵ���#���W�[�ogZ�v�5�q�$mQg(�i\g�m��E8Eˌ�.�c�F����L��R5.θ��˦ys��O�h�Ǘ�o�r�=%R�]�9˼�@]ϔ����2q�-����}�U�l��U�`��(~"߭s4 �7��̮�;�e*���!�Sˎ`ݺ�񈩵���S�@{��փ-{��:�7>3��:��j0!�N|u�1I�a��B�Ì�\���R�7昃�{���A��O��$�է�
��:k�:�s�v�^���
;ِc&[��� ��
��Wp�޾�����"$;R����\[�sڹ��*_�mpU'�S��FϜ6��/*��1�S��E�~J*Ƀ�.(��S}�4.(�9ҹ�lZ3�7������Y�(�]��4~�EcyT.����	>�qQ*�L.w�Ś��͎t�Sf"e��d����	��,�w5:���pĨ�K�*11MB�P����@E�{k�G��e��ӂ{J��dc�p��&8K�]3���5<�ͧ�&b#O�N��L���gь�z\T�����3@4�x92i�3z/��Ҟ�g�<h>/KsQ��{�wQ�mCMG����m���P�H��ʣ�ܳ	��8��^�n�>�w����*��J�'җwݔ0S_�>�C�2�jy�T��6��%�(O�T�DEJ{D�my1�B��*����`��J��o`���iu]�Tu�ݿ��g�̓آ��(«[?yH�l�bO�0Q�|�z�T,�w6`�|�!�}�`ޚ����f�O�xb@C99�F�����xX��"B1��UА��א0"�̞�u�k������*K�pWmq
oI��̿��oe��=8������H��m�%�l��?19P2�JI��
�S(e�ɨ����3���_�U�*F�.�&�f'7D!F�8�>��2�:]�i��Z>ے�I|��"n]��v�M�W���St���< ��}ym�u��N�u9[�v��G����+lN !u��F����p���������&�FuR1E��7V�	d��#|��+����68FOȄ��|�T�r~��bf�����η2����<��7�N�]%3:b&�t�V��(YX��>�*�
�����P, Eʏ|환F�=��EtӥC4d�op�(GT�]$I�~�?*����ZY��"���-��׵2�����q�yo�a?C � ��$�;6�c�Ag=J=Q��ڷ"R�l��Ys��Y�ۇ�+����%z��oO�� �f�?����6[[S&�$�>�h#�Z���q��8O*�Z�J0��W)�0��0e\���]5�tE�Ѱ��*s�v/�gcڡ�0�h��<{��	`��t�j���4N�Б6j���z�`y*"�p��;f=�A�}x#L�W���(����I�ḻ*�ԟ\pϻ:=(ը�}b��|W�Dӎ	�%����3�3����Yv�כ����uI�\�#mq������{)+���IA������"8c3|�LL���i�Q����X�(Q�wE7�){=q�C�1=��tiz|+, '#��(L�C0c��Q{b(�%n3�i�t��|nb�n��_�Z}�(C*g=��G7��1
.m@2XW�-����V�?�X���G.3�3�!��c��y�zn,=�~q�{.�ɥB~c�o�]}8fᯕ+mr�B1ʯ�{p}�$�C�r��6	����>Qm[�b�vD����g�M��L�S&wFL9���>k)ߓm��A�P_\D��^�3��}�g�r|�y댔�^�(76u�����\�Z�#2���f�.��X���� 6fpCA� �5)Hcv�	�-R��ꚗ[]�y�����n��'gp��,�{�����3{�r�����'��90_%����r�nn1��u	P�#�TІ.�&�=}�b��S*�:��p����ס�R旂�3n��! J��V�,|M�TP0fG ���yLvҌ&��]�[�YM�Ib���|�����{����
��e}�����1�~`�>Q#!}��	Dh��sm^`U3�l�0�W�YZ�����!���H��"{%�f�pW��Ay�������(�>s*Ӝ�D>}�3+�]Z���$Q1����챯�b�=="zak�n����[m���Q�1�A���5H8~+�\X[[R�nQ���[E�$z a��e\��ݍ���*h��΀���`R��D]\�4����,���A%}ꊊ:fM���u|
��4�n��|��|���f:gԝm�e��|>�-�?��L׊��y��۔D�O�����0^��	`}�T5v�U|s�R�	�|�*�Ǝ��=�{ڜ<,�2r�9{uP�+���Lx�3�ʉ�^�+�]*��^
5�'��$ϛ��r,	��LP�m�?���0�d%n��cxCQ�^�U�vx�$��}k��4�H1��D�50}�J�8W3VyT���MSƫԤ�P�����1��W�%y��w6^1]�]:�be�p;P(A&��i�S�捻Lt-�j�P�SAYy�s���v�#��d%� ����g�3��� ,���Y��.��1�HfPoJ�]3�6,=Q���l��6.�'x}����NE�9��>�"/eB�y��0.+�󊀭I�j���/gKB��`s�ڜ�\��t�s�VR����&����+�)�cQ��uҧ�N�i�ʨ�i��K�m��7�-�b�P�����hIەKӝBS#{b{��1r�3}ԨmH�YC3�tr7��wc���!}Ƿ��|��v�9���c����T�̇�ӊA�ڦ��ݏ��Vns�T�0۹�B�Q7�g�=ŏ�̿�q��?^f0���[��Lt�J�G�E��J֨~�E����!��`m�P�8����o���m��7Ǭu��v�4�kOo�<��B����Z	���(���rtR��Z�3�:���Oj9]�F(��p��#z>�s�;����8�NIۈ��G7�����u7,��3>҈CZ�.o��,�٧*��}}2��6�}���V*�% �Mu��2I�a��at�g.H�b����dR�צ��e�k�S�����f=�EL&�y�����>�_���l��QF��mg���]X߲���OL�(c>�e	yY�Qi�� �wWPU�:�l\��c�tn,�7ݩ��W։/t���{}�@��P�
�7��K�)Z���+��S�"��j�;�1In���<�b�Pݥ7Q����5�];� |�^ڥ8�)�S��Y���bz�Bw'{����N������`{c��١�p�ML.}������P{̨�w΄����9�q��WL�R���[^��Y7�@�e�@��aT�J��*k���PY�9s>��}�`l�@^5���P��[�1 :�'q��1�9�K�Ny��_}��9~��v�4�:��r�sJȿW��"/��,��}/Փ�Bs�_*�{oN��}<��X�4�;�w�ѣ�{��OV�?om�ޫ�;R�4�,��h����)f�Ҩ���E��"�2�Rն�����9����aTm z���Ʈ�9o����+Z�@� -vt�A��8��8�J�a A	F��B�\�Z�܍�,����
�,�V$�yl�bfl�(-z�'GJ�����hs ��E�nn��ט���f��Ռ�/d��e�"�xm�������A����n�铝�G�;��4z0�r�̃�4>�V$��@WS~��/ф|G��}��`�i��O�S��[ٍvH�!�W��]�x���+!7��BV��_���|����+��X�d5׺˻���p��o�eܓ�q���9���Y(�9H�Qƻ�f��N܏	�uy4�w&y\1ST��HK�.�5���=F�7L��2�KoW���L�\�E1R�~�p��,�o|�!���t�٪�����2r<�E<����9�^�;�N'�|:�uF�j��Ã�G�x}�PZ�Fh�����lD�T;̓��	�ꊛs���{�%v.��r�ʿY����^z
/���I��C�Հl�*4/H��/K����l5MEA���A��P�T>�4����;�5��5Ǣu��~�n��9��1$�/qs �|�Y7ؖ�)��Lo�]�Y�aF"b.���jB\g�� ���r�ӽ�d]^a��Y�G��;���k����qu�n29��&��J�G��ϽyCB�>�&�S�7�F��H�S���}X�I>y��6s6�'�_R���n!�ZL:9'+��=옪@��m\�(t�GQf���cG�E��ɯ�[�z��At�l��/{�D�R�w?���(�2v�0R�;\�uTh���M�}%9ў��MB�|�L���r�Jy/����+��2�]��b�rcZ4���3���wK7���`e�9�})��f�<\j��Xۗ���̮hl�ղ��K�b����w�TU���Cܻ�K��SiI����R����;[K��ռ[�8ñf]�uq��1|�ON�t;&\�7@j�����ws�a�\�k�v4����	�V�#*����l���Q	+�^U �9��Cxl,�,�8�K�Y�ѾC�ВϓNL�V����F�&:��
�9ʙ�_sl�P����&��L�B]J*(��mJlIAgZ�[��ۃ�n�)?;i��9��?`Wk��ӛ~�8L2b�YZ`��������:ƕ)���)�>t�-e'S�*L�}7�B o�Ⱥ
�*2�x��u�&�kn�:�k��Zb��tĀ"��=�����.<&�-����
�zn͛��ɽt	����9ʍ�Q�y��b��B*R���&(���8�d���ި�����N��OIj��o.U�r_�s��k��i;oMJ�9�yDy���W5�r��y�L\@��>�I�L���}�=�G�y`����(m���q����/�#Hq�-��6�{����=�ʘ��O6��b��"�ߜM�RˊOH�}ތn��mN��_D��DMy2jt�F�<ؑ�V��&<��ls=3��f�w`�B�`D6�(Y�ˮEE ��<���
�f�L,8��)�;J�����դ��+���a��3)��Kp{��G����^R�T��O�%Uh���m-l*�^VK���itV��qb�O���NqNE(��n\�<��;\��a��:9Q���ks�
fc��g&�p��\9�����Y��}�\�\A����[���#c/i��`ˬ�F��5�m��}��"4i���3h޺�50%Wxs���5N�2�vX��VѝJ�XJ�%p�B��ف��F���:
�j��U˙�i��0䭫[�m���v��̚�5oeEKJ5��R�[����+��!�(/���i�DP�}W��q�~�����@�����'��F���)a���7����ڸ��k��S�m��(�ef������g��I��w��2GOJvj�N�nٚ��x�m��с1.��QȌ��~���
3�g]�tb�mܺ��l���.qU)��n����GA��9�l�B�/���P��RbX@�Tt؄aͫ�F��ʔ��S)
e�S��c������K���zp3�d��r�Q�&L#��Wx��5Q���T�v/�z�Ku߁��qQ単[��o��3��z�������=�,�r�=�"<7,�;�y;g�˩��=Ea_��8`��p�Bj�*�GmX0����PcG�fz����x2����	L�7B�it�o���Y��~e�/�Ȇ�S�/�j�tU���vM�y]	��o�4.{:B�e������֢�/�O�<ķ F��Hrw�fch���Fa�Kb�ʌ��ZQ�5>i���v��!�W�0�9y����1fr��<��ޙw�ų�{s���576= ��vNFOOJ�
�*:[����ϪB\������D�/3���	W�ۑ?����������ZI|)6b�s���^Q�Ƿ��]Ml�]x;T;����+U�T����}���Y)Ȼ!G���9 *�I@���%7����X{:2��V߇���l3���S���d���Jq`p�;�q�+3we����,*�V�}2���خ�nf�㫥�+}�=��ҽ�49�n#%���|����#De�xt�+�-а$HMeC�%��^-a��R���!�N�e� �]���:�;W�z3���c9��^�ݻ��-��ǂnd)�Z�E.�7w+�c��nr�VM�x��۪;K�R7'V+�P�M��r�6�G�w<���`��>�ް�S��m���jbS�[l^%[ZQ_n�*�d�U�d�B+%�a��F�%'�On���Z�x�����X�:_V�����ܪh�L��Ԩ����\G<ֈY���n��i�=��Ъrӊ�J� �t�ڭx:��r��*��P��p4�X��5�E��"���z�UE�e����]�\��ee���w�������h�7kEv����� ^4�j�	�2@]x	��tR;!�z/�R�	K��a bQ;wt�I�����&�͖>�i�T�ɔ�w�ݲ�nu�U�3%���x��#f��7��)�US���%���Wn;7�{�b�m�5M��"�t�i��(&Z� �Z$�֥А��z��5i��	"�����aN��|(W[���wOw�9B�l#]�u
�f�E^�:$j ���.�����\�M�6�G&3R�ɩ�*���f�F��y�Cd���9c�QQ�4���n�u�à�H��ky�b��Pc�t1p9�
�ggq:됀��C,��
��ޠ�p'+��$n�� iTM]�纛���_�uu2/�ɭ>��ޓ7!�$\���ӑ0w���(���� �����\m�f
wy0�>�_��2��ĨWSݲ������|'N�Қ1ȳN38j�A<�1r����CNj&\u��CD]ݫyHm�y�j�V��v��(�e�{l�}�1�ɲ�=cL����7�ҝ��B�p�"	kJy+CQ���MKEڧ-�)�U�J�D/��5.�1�*#fu����*(���qoC;��5��L�+��V���!�g�u��/��@���߯��B�A�;Q���co ����2�5l�{/�<�[�g���;r+�V���_vo9)oj��������V;Ӕk�j]e�4��RK��ڼ�b/U�wV���G�f���ז�����P��mnd~����);(��q,���3uJ��@���2�����A��:^�ɸ{Vr2]�CX�P.�#��Z;tvU�"������e��I�Z�s	��b���4Gi����ŷnq�i]�}�V��w�z��w���;;���5�ޱW��F��v��r�N�&mP����x�s��
)���n���C���D+sE�o^)�:��1	��N�����Yqd�였DC�0����cU���Q�q�K�mIu��۝m�a`�\NKD��^���Yx�m�DszDv��_�8S�K�
��TfR�ջ�ev�=�g2�4�����S�w� 	35��O7��:�.
ӝ#��^>inQN��o7w���+���Y�����	[mJud��8��
�jǮs76nKs��h5n� &���&�+����B��J��[�Oe���ND(0i�:�v���&Ί���`p��7�_�ysL{t���1�é	�;r�&3��0��"y��X�r"�"�f\1�n���fLv��~����&��t{��4<�0��ia����ҋɊb �%�f�߬��H���XV礷��+�j҆���������̄��U�o���\h�iz�Ԯ�%��a��M�+@��(��*���f?�L�
���[o�pA�>�Ν:�}�o2��k㺪X��<���(�,�L��b�}5�ŀ�(�o���d�lA�?6L&�	"��4����E�s��c�����ݞ;�-�L�c��c�u�Hݽ	�~��껴]Qm�|���K��PЋ����M�X엧k�<���3���C��e�v]&E�H"�P!��ݺ�#�1�vQ��=���Jq�U�MA��\W�TxL����q�Uz碑��<�'�[�g�����eY�Z&���Tv(񉑂�֚e��b���(�4>>����Ś[YXM���������6>�����s���zf��΢���[�����m /�$�׭��	�~��+�Wu��^��8F]ld?-��eؖUa��+^4q��j�	�7Uo���*��R;8�Jv��]���l��a�:LJ�x�9��
�X�Y��y���܋4�:�5�%:�pn^�*�H�ݒ�Ң�S�bL��F�P�=����Jْfѩ#�����94$�Q�����:�ٺ.�,�M;������%�֪T�'~�����U�L�C�/�й��ة"���q�юC�%OA����6eY���GU�p�U�V�y�i��dU �n)���y�C��W4�� ǲ�R�`}�q�O��^�U���@('6�{�qWw`�	��N2�B�I�>�^�\�mw�x)���G:�v��F���1;3�!ޖ�D�5�4��&dgِ�Z��B.��\7{z�ˢ��yuG]�]0�+�o�?;2�c��_P��ٵ
�*[��qN�)�uóy� �O&g�i�[<�w���T�7ҕ�Ǯ��d���"s�(/WKzri�}�1��c.e���Պ��:�z�`2iTH����6o�q�@����{\^`��^�������?~P1=_4l�3�3���1�W�Ef9s���������\rF%���>���Y����N��]h3��N�W�)�/���<��N$�K�<z orV�RϪ2v�z׷v�
���C+��<��Hr;�ڡ�x��\Dv}ڲ��~�>n>��?
�X�ͷ��4�N�~r�wqaC�P�EӃByE���gE�Ӷy+�����t��ַe�fj5$���<�ؾ������~���9�^'�o�wY�˥]V�o�Z|)�S8�P����&n�����W��?�'D���byy�P�([��g��b�Qv��{�s:e���u=��fή2��o�S��+=�;]��W��}lS�^p�)��[���Ce��M� ��;�n��9��c�	��?�X���3��x7(��fI����8�:�KtnC�oL����S;s�q��	8�`�ʁ��L���g^��,N؁�Cm��k%�roTKsV�Ģ�z�+�=���^��'n��s�"��]<>��	�_<섣L��.��A����򆷙��{��՘a����}՗S{���N}��4ps�!�L�r�0=���x��j�q�x�Vgp������|6o.��{s�T`�����O&`v�!lg)VzBa�s������Ԯ��-C0����-��s�2�dx����u"f\y\Z&8�Yu"8T�5Am�O@�1������ �����[�C3�������Ô�ѾT�{�y�� .��Ө�1�s��y�/�����
ݨJc5�\��k�(�Vt߻�+�(C���_��:u������$�Mku?-7�}K�ɜ�+|��|}�����6mHq�u��zf�Z���0n���=yt�xo7ϔ{0�kz�4�a��"�
q���=w}wj*�Y/����*���V������Q(�{�J��xvV��o�F��_���a"��]���!v��̉�gr?<���2�>v-ǩh�f}=���&ȅ�[�ޤ�8@��7[e��h��v���ږ�^��~���OT:�a�9U�R�#:h��:+`���O��n%T�3&��=��r�\9��c'�#���ޫ} 1�͒y�]V9SUKW�xxz���G��9�Y�`5����]�	�FP�ZI�E7�L�G�N�<i�f��"�u�'�,�Z���� $����UA*m�t1%��c���ؠtu� c�
�R�αz�J��9P.U�����B�&�����#�'�����=�����>��^����J��1���QV�����.˘������{X�1ݕ�dz��9�F@��y\�V,DՉw;�������g���)���j��`p=��3r��YPtt���s�<�.��l��Mcج���q��YP�,7��帓�'>��~�U�4On�8��w�.:b��'h_U��=��v ���r��5��y�XQP&�MVϵ���A��}�-��jX�V����gybA����"h��s�u�)��S�����5���Ǫ����.Y�qc�Z��m�s�s�R�X-��6Y�&_��"�F{ҩ�{��Y�y���!���L��DN�]}�u�^���;5��<�zm2iD��D����E^�b_�7@���UA�w���}n����z^)FN<�#�������E�1|�#|�0�#�U�;�ϭ�+�A4G�O�1`n�T��j��жz��]����@��,LixT$F͌��O�\����5�웄u�'p���j{cqݧp�E��I1L�'�*�;��U3���meb�pz��6�O�6�^S�nc��<Ҍ:F�.QT[��+�䩔�xr����o���+)����Bc��j�^Ϊr��/�!�~��ҕ9/��Ԃ٫q�wwK�R߳� G@s�ȥN�7+)��x^w3;�WQ�8�yq'�$���u\�[��U�q��A�6q���d�6-���e�:uXam�'`� n䃴�"��)�	�/2����J`��6���"��P���l̸��4i���p}E�`�)%��̵��s�v7���-U�Ƙ&������镻��ґUQ
t�T�:t~�=�[����&���h��J߬���
OZ�O�7|:�^����j�܏����~���ϕ��1\0j�����*����%]�b��Yz��^9����*q#���{"�����wk�`-�~�;�nlF4ݭ�5���R��.�����,�RZ�k~Tp�O��3r��0g�)�VS�t��q�%%���ϵ��_a����=��~@􌓇�$�*367��맲�H�8+�s=6��p�i9=�;p�<k��N ��wN2~{9T��mO�-�q���23΄�Y'� D.��=��C��^^8@���Sc�)��q61�"��@�^p7+'Y~��[+���k�Uo�\b�z��8�LM`W|��w�}c�B>�q?V���7��"�y��b�3�[�����OOh��}�-�6�\'��^V�VE����BOiW�77�*w�`fSN}LMs�_��۫�>�x}p2�fx�`����T�������d�����L���+J�U#�~��'ϜR��ɇ�>�o��ć�~�/�u|5�w����F�q�഑�� ^�m��\a\�J��_Tq�}���ׇ%n ˫���m�"�o)Y�,k�U(݆�����)G0�㵏o��:Yi�?�1���a4��~9{.eȒ���&� ��jb̫�κœ�M�9��5�/2%�V]���4�e��+�7���L�Jx��kV�T8�S�I���������x��ǠZ���'o�/��W-C�K��.�����m�`��w���^Z>u�;��q��2�|�{�<y��p�-�Ex���^ځ����gz��"]F��ΧK��0��d�6��{��.%^E~�*�[=�fbD{��P��c=��ON���2�T%**H��� ��)�����;f�/��c����'��Q[��ˎ522��h�=�h�;���9O?Q�D�~.�.eC���z
���'&u8��Ѵ�yg}�c=˪�ș���U�Xl�ڵ�x*5#���N��=��cd3�۵ZF���S0�N��,����>��9b�X��,�[Pg��<��uK}��0�w�Ϋ�p6�2j�*�D���c(��������NB�3�*[��ɪ<cOL�ꖲ_�D{@�V.l��B3aOT���~JxӚ�YSmg����+\�o,��݋/��`�����g��̻.���%�2��@6��ٱ{A�M{��
�D�;����4���v*���R�+���?t� ��/�w�z�YR���eׇ}��*"x��r�\'��	���f��\�dϟ��Mޣu��g��Cc����l���,�T�/Lx/�Ұ�ʋߜ_��iR���teY�2�Lك�{���tB�u��<=qj��7w�n۴�Qިw���Hw˲�1�v�����Zf�'k7̭b�B�R�q��p�p�Y�ʫ�)�����*��9�rS
��O�if���*-�}75��O��I.0on�L��u`RVc�׼�3�e8~q(O���$���=�w^���;�F6�f�r)���_kKg�f��l^ѭ1_v���$/�8�� �t�B�Q��bC'��v��uf�|�g0��2R��9j^NI�<���هY6jl^v{0���D�{]TP�o��=�|H�zr�Epm����&��.�_�um�r�m��+��Y��	��
;�x��������ꪋ�G���e�	#�;6#�����-d��3vzo=7<���酲�x��8.��g��w{*;4 g�}�9���ݓ��>טT3�:S5��=�w5pn��>>r�:W�κEM�*��_mN��#���)9wl��{� �Jf�,���R~�Go�U�I�H�l�еɞl��N���vfi{���c�E�t�=��8Q�͘j����
%��/��>-��=�Y�WUk&�g��U�9AW�v���9F�[����F�������ϲ����-��7��]9��2�E��6�~ѷ�_u��+�=-or�	�����G�Bu��Jd5�$��T�$=�1�ۯ8�3x������u�Q$�m�&eH�W�SZ��F��l'f]���+��<;���-�?2�t��"���C'M�t~� ��`��Ѯҳ�)d��I�d��<��*d�a�x{�$�r�Y.�OpL��a�$�E�i����B�}B�!d�Uu�*��v3(�n�27�?D�R��*^:y����.��d����c�X�2B��Y��&�q�*uKb�М�@�8D���]�(�>p7���0��~�T��fA>�A�##��魡>Q�#*��^Ţ�j��vW���6)�mTq�ܫ`�R�=w,�,M3�[�}���-oމ�l������Yi�N�L�[i߶��J�﷮}�������f�o�9v0��)FlL�o#�?2z�c��5�}Ep=��3��P�id21rq?s�m���C~ �F9�*Eglb�O�2�|���E�ٴ}������E|���G�����f�|�O<� uz=�U�"
�v۞(�y�Ҍ�����/ξ�Û�*�F9WN��m:�"�oy)�'�Ȉ
Z�z��������g*>Rzr�
�P�\򽆷2.1(�]�s�_b�ga�s�҆O���ga����i�e��U�"�IȊ?�?��y��z	�f�P�>յ�=uV�����t�A�:
f���i��@T�������{&T2F鸮��#��}�eĻ�������Z��Y�Q6~Vve>�Z{���^�K�^s9W|J��yu���y��;c1���)|��cjZG7o��hU�o�8�<힄��!a"��GZ����0��;�la鸧s�c2AH�V.f<n���͝XS�7�J;ȱ��	�w�hs��L"�EPOv�=lI�oE#�
Y�yˇ�r=>ӑ�{`f(��n^�+9��M6��dPۘvQZu^�zeٗ�U�-;[Q`Jz#����:±��L�=��_z�����J<,��i>}8k�����/ӵ>9ǟ�C�/�UW��K���T��w��T-y,$��:�u-}Ĺ��׮�S���kԮ+���}.�%oq��f����P�� g�/��9�v�㩙�eσ������
��
S <�ɮq�K9m�U�[�:G��2�����Y�����ڗ�-gnUZ.s�����6��̧�_�3u�{�pgg3SZ���CsC��^�s���O%^�5G�ܷ
�Q�_�SB#cY�=ŋx���G�-���Oiar�)v�Q�]p_ܻzHjCh%�dav�f���qus��A.�7"u��c�f׮�_�o�/��^�ۤr�}J�{lw.����q�k׽14��Ǔ�Ff�l)�W�^���� ���s�/��;Y��GJ>�F#(��g
D�q��w��j�,���:����򫫤v����ct��_Y�h���w���U����3����"��y1Y�Pj��S}5&e�[�H��^��gve�c�� ���D��Գ{(w�����@��{�S�w��=������xXo�p0��"�	~��EtyȜ�]B~`)��r_ϻ�j�Lb7�u��{�X&�w�[HXk��hdI�꾼�;s��[���c�Y]�i���i�5�N�%W.�����i��P�S�7�r���5��~3v'�덡5mUq��P}����ދ�i�jne�}+�-�j������u,;�]��2��_��`aYX	��/������ާJ�W%��O�DG��ybYҖ�o��/��jn�=��,�W��ͧ��g,�䐫Q�uE]�ddj�X��rz�처��* ��Ǒf���n�ſXS��qOه;�����$�=�6�{i�+�_V����u�@:i`Ϗ�f?Jr���@�b{*FOe[�c�*n{ف�l��̜W,�����
�������|��HF�з�.Q_\�<���#_���|��;�|v$�獵��[�u�`����j���:�@�Hp�1N��+��s9����rZ�M�rVӧ�����e��C�tcJ �a@��u7&�*�>�:���Џ�:��:���;�fa�3�ƭ��B��Y����j����3v⇬�vN�~"�w���/�������|5�����}t�����N�}�O7H�X�5�\Q�HVP�N�˖~�'�/�����_{�����^�:ڟVO���?�q��"yb�)^��Ƣ�*� �Z���l�%u!����V�<'ϓ�j��o��ѿ;�;��u��y9�!��#��X�;F�]�Y΂m�q6r麳}Rh�UY�@q�4����`h�<y�ue�&��]<���t��2�f�D��\����a�UI�堀��ёi���n�>��-ֺ��i5n��1��t�2s%$b�|;��١��t����[/%���x� vLqN��F�ף\ё�ͲlStB����bV�M�\�HX��T=��9:勋�6���fH�Z)�噖�0�&]ٖ���#r��/!j�@#��E�*J3�(	Z�ՏJ]:���e��Q��J�{��v�,!'A&ܴ�"��e]\��"F�%�40ө���)���Ky,�cj�Զ�'L�v��"�)v�fF��l\Lj��_!f��em{�.��W+��N6�n�fub��j�A�ʔ:�CR��u�.�`J��)!i���k��Vۣ�ʰT�mܝWtBf%�4�kLN$��W�㟜N37��7���[s}[ֵ��D����s�q���w��b��D�O/,�w����uj�b���}�>wA�2)�,5���6����Q-�WG��~��W��Ӄ�ԫ�x���Cr�P�wۣ����^��n�i�X�mX�b�k�ej<q�c��@x8�_V�P�^�5�� aE��z�n�N��$��Ʈ��s����+4&��zX=�����L<{B��"s!%�4bn�e�ᕛ8���٬�OkU���j��t1�컽�IY��5^ҋ�X�뚀w�K���u;�� ek/s2������5�$����Di���^��
.u�*Io(��GQQ�y�#d���1P[@ͬ�u��7A�����@OɄ�E3GQ����R�]�j����û��)�u��}Sw%%�-�]ҟe=sn���֙	yB����g�wid0�҉��`�0� �]�ovd~�@}9K�t�oV���[�
J�&M�'���S:����Cy^�B;K�Ý�HB�8v_gN�2�U!7�bP�� �U�ٹݼ�X��?�yw�N�,�����1�{�yZ�J���M�24k7���K��C�C�l�)~�Ѯ�l(KAA�n�u|�v��
F�6�K���6�k�����&S]�S��[���4iٕ��x�EgR�@�D%>�e�B��,}S0o%Aۭ2�k��U9L~L`�C���mҦ�72wO��O���T��E��wq*�X�"������^��D񌞏o�D|�Q���l����bFn�[4�GX�0@+F�l��j�7@�"��$��1P�%�]�Aqsc�*����'X�y�N��EJ�1����4�<��ju$�݈ Q��Fn�뺳'��LݾzC��ҷ
{����*������p4��5���v8i�+�{qj6h#Xv��o�*QF���_�.�)�q�|d�w7dYC@̸��-pE��s�k�~��J�B;���+���������d������&E^�\�GtV.Fު�v��RLl�hw]�>�,vegeus�6��h�Av�wf<���pkr|�3p ��a��҇k%���}�D}���qyDWM�0�r�A��|I�~�nj�uz]WNމ���kv��,�fT<B�����) SN�ei�{�
;`EY��n�2�@<��Q*
�ı��oc+�z;*^�r����R�+�|���!^c����ڌ�5}���=z�Jբ��T�nւ�������jR��P��TR	ȁ�۳:r<9����yf,�:�� ]a����+26��%-�9�1ΧX�n�Q���}�^���K�Z��e��C��g^s5�J�G#l�xӁ�)��Ò�39=
 �TЪ�fG�٘��Ô���f��d�$V�Z�*��F*~އ�Bىӷ2�k3� �oӎ����F�vO��ٓ�1R>Ҡ�볃����4�U*���Ð߲�_������_�d;�uc�-�]+n
��4\��}�e��{̓+�;J6�������70�[S��B�����gmf���񖵾:����/!��Pnю8�D�T��`l��=��R�Pމȵ���G�ο:�C�*9߲�At;̚[�y�S�q�u�RkT���wz��y�fk�=�PXty��C#�1��IB�5a�&:�^�7hcG(�Xj����Ĥ{=��	�*[G^�~���_y���m�K��}h*�E���o����$��6Nl5p0�������p���qf�틞�(����jƳ�7��{ <`g)�IY��{�B���@�͝V	�|�i��T�@��y�+����&Vfә�N ���Ȇ�	WCC�u�ޛ\f��] �̌�P�Pn�iƫ�f���Q9�!6���u��KseQ���=�>�nm�*z;��H-�&Ș,d��:�Nnz��1Ct��9�_okFu��Ƽ����㕈<�x�W�OQo�*�}r�[�6���6��[ �<U�C���V0!q\���ټl�޹ٵ}*�˶�K���w�Fj6���Y�wF��q@7%��LJ���a��Nw�3��n	^�U؎��P&��0]�ξ	Ј��ؠ;�r�]9<���U?T/lO]�*X��rߪ�$ă������?�����t����5�!o'g�)����@);/�n�8�
t������롈��>���R��g��)�渗�ᐧ�b���mA~gh�n_�O���U̎�t�%�zȍ)gt��C�k6�8���mD��c}c��/Q��C�>�Um��������?�N���<)��{�U6&�幗ȘWޯ�^�����9�j:�\ݸ]�p��*<h^"�{2�,z�[P�VoVGRa�zP9���+��9�c)��r��"6���E緭Q��W|'qb��WZ���7�窫!s�eo�M�հ��8̚�*k]��Z����S�Q9��˶�xrs�kN�b���S��(�jƬ���їJ���ԝ�6��Yť4Z��Dkm�=�5z��p�eH�cCۙ[�+�A��u��kh��{��ݦ�[�I�������^��&xrY�S��,�؏]8�C0�.�*ZM
ލ,U��A]D<Ŋ%C�{�Gr<��Sܭ\�zZ�^�#�XWm�c���|-���*��S�z���4X��O��6ftU ��[5D�*���-��@[U���d�t��� ����WC��/}c��y>(�9ك���YU�K+0�tn����O��
2zyEwjm�g�g��-�F�����5+c2N������x��ߛ��t�W��%��c�˫}���4L�v�&���AGZFiN��^��.�u��vN\$�z�K��mZ��;l�Q���W��kƼ�E%�iC��o��r2��aS�0J��u�zj_�n|~��|���f�����ݞҹ�9G<jN<�����]Ĺ����:\S��~��u./�¦�[0"^k�>�.a
A!+��H{�k��x��=%Y1�!���fx�mï$f�rr(T�Ӹn�9G��a>����jXY�%�Ĵ�+�����a����Cν�Q�L��\���d}ӥ�䟵G8�'R�`LdNC��D��y�RF���S��Ua���2\�WC��l�\�m��M0ʰk��}N��b���܋{zh���R�<J��.[�-lO�����BL�3Mؤ����fߨˢ��ޙ��e8��;���\�8�2l��*�Y�u�g��I�岇~�����M��E�/�q��q�}�e�=O%�ѥR�Ù������r�i�`Qv�j�B��+��ipf���!�:�Zn��8u=�<^q\�Fl;+;;��x�UOPy��$���7�i�gڬ�I���iᅕ]wj	,�$U�3���ܐ�+���Q��xP��=\�*`�_������B���GKU��������v&oj1O�V�j�{o{��j���K�_3���Jt��o�Q�vM��s.J}+Xwﾌ=�9z�75,K�D˾�!ͻ�1�R8���Y�7s�7��O�5r��3�����F�X:G�y�vşT١o�i�tq�^~�Xx���7K ���W�N�o/!Fc���� ut:� U���X��⮽�/��k���^�}\V�G8�|����U�l(^������|��b��(�O�Ս~�w��a�g�K�aþ�1�}�7EN����:��wK�U��$�|p��z�A�:����<�5�/K���9��6xo:<�:)D�g����o#d��p��VO^d�o����b��C�$��3�j[��y-kxP�[��qɌ2����)]q�����Otp�G����%=յ僵�S}6�_�Լ���<�C*ki���>Z�)�MV~��"��o��� 4�s����zXk�2j䈖�+��Yg��eaΠY+rO�ޚ���f=���C�U���8k8N�!-|y;h�7KԸ��{�wQJ�c����:�s3{��;���x�n��\�� Ά�Vm*Y�ts��L��G׺ws��ͪ2\�m����췏ot`�-'}v�,I�B��7u��lG�=����h�~㶎��?8��?I�eʑ��/��ã�y��S�,E���nLyYJ�>��!�|����Q�ڭX悋^U���>Ɔ��Y��PW;G�y��;��VVׄ���U.�����nIV��
z�um��=V8�'M���1��=bit�Y�����
�Le�%ga����g����	�ى3���r��{<(�i՘��5��ewÜ'�H��Z/����&r��tB��{&d>
zxQW~�9$���k�9�^'ڨ�WObp@�uGUq'��V
������@x������A�N�����#R���-v0�cQ�
�T�;Ӗ#���R��/C7��*���t�s�Ra�u<��p�t3���9���a]�q6NE%�����a�1���*�+4z&0/�]��t 2RY�-��J=��B7=qP2	��73��>��x��1�L��l/t�e��}aWm����}x��4����,������ �V�E�=���yc!���
����=�!����_{ɪ�3��F���`V�&9\���<�(����>:�>��G�l��?�a����>�'���W��epg����
��)-鯪'D�sM�Vŀ[�|/��!wwYge"vP鼳	u�ݾ��s[n�$P��e���R�5ݗ��SK.�VU�y��q�Ե�@�J-�yr��d���D��QS�0式#��>f:�Ubm�ڴ��r��m�޼����]����BY��4GU��~���&��ȷ���k�6J��"�qY�/���w�]�Lz�Z��}�S+Q�ܙ��i�N���_0�a�����_)`��zj�W~F�]�k���x�7�	Y��;=�Ҭy�أw���fc���ԢX����+������� {2Y���Ỗ"���er����N��a������өƷ&��l�k�LKb�Gk�ɂ���ź����Wcgp�!�Ln��~��MX#�q�����e\��u7'8¹0��L�Jm�^(�9��K3}�Y�Z��L��`T �fb�
�nz.3�&�ܱW��~b�?f�)�&���ZʱQ�R�Y�(�7&ζ�b����/5�������1|��_�WQ�ط;�7�϶�e�s4�}����.Wt�DD��x�����]�
���*��7T���y@��}�K-ܡ �' ���]��*6����J����<+���'�_��>����/:�n܂S����`"s�˘���c�w���Y}��9�a�R�	0��z�MG��Y�L�3�(|�gM�]���G(�[�Q���ẃB߆0h�BDvC����&(D��0���	6�Tà��]��8���Sק*V�E��ʻ�y���7�T@�;Iݖ�w�u�V�g���:� �gf�y)��6j�z�%�F�AS|���aH_I+`��$p7��fc�x�!��cx��p�f�K�6kK�yP�}aڮa��o1Û?�/ި�_��#&8W�&v������ҽ������	���_.�b��<5�W�\ �=�������0�y%o:��&h^��� �v�(ο/_t�U.�V�ю�ge�Z����P��s�dy��� �ˍ�[�/��5=�#�����=�z�� �Y��_C�'ި�x��*��}�2v�dX?X���Ƞ��F�ta��#�[s�����k���X~�	ty@#Y�-cw�SGx���T:��^]� ��<��~=��K��y��^��+����/ǀ�d���Z��a��>���?G���u�>�:��������4K����e��FI����y�ǜ�D��Z�섰�q|�n�
G���ف1k�LQ~�`s�wRs�s���՝�"�������ՔLk<�Q�ǡ������'����z;��'�մp����o�u5��;Ӟ-��Rژ�n/}Q��A�������*L3_Xuq�t�E)�y'9�����Y�ΐ=��ȋ�n�W����pѾ�^�Ob�I���D��V��V�m���܏t���Ț��/=fI�6�SgFEг��c�:�f�u4Jͩ��F�>��'b�u8m^:pF�A\nee���!��>�fǩҧ�@KP��rP%-MI���F��rEJ���}�p�(�w6B�Q蔓�{y��R���L�ؽ�]�k:M<(�ȋ�b��xV>�ϲ��A��o���/�a�]���ȿFF�����{�v1���q �0�����|�䍪˲�ђS=9B���Q���j�����FL�~�oz�"�zGc/��(��Z�)T8�k�x����a�RCۨc�^�31�*%[���彙K�o"a�%�S�җ�{��%�袐�"�^�NY�<��z��#��*���|_|�Xh�<�jf���^�\�/��&穎�b�UkQ2
�!H��}�o�,V�yUh02���:���^���؎o�|y���k{#z��W>Ok�n��]�r�ͮ����N���.=k{�L(%B
��p�M���峀��6����J�=n�VY�vb��n��
�5'b����9ӌe�oy��z���/�z���k��rrJk�k���%�P77�y@8����ӥ8!��kU<�dܫ��T�n�f�ή�w�g��N���5MWoF6���~O���(ݳ=��⸔O\n���A"�c�y��~��ҕ�
s_���Ԉ���;�a�r}��2/�	
L�O�r�d:�vp�[�t���176 64M��=��*�(蒶����K���:V��n���xq���gҞ�	��2d�My�����Wǰ��师[��h::�:�;���x��@c�Vj�˼�!x�
�r�K�*R�Vc��*Y}�Ӑ��,��:짩��$=RW=�||.�?v����|�����}F�TX���-��W��dVNQ��HP�lN��`�t�s�.D=dF!����~�c��8�o�F{�jVD�CMF�z*^a�޻��Vfqؗs�Kܯnm��ut[:}��������|k�"&�Y��`WQ&�����cb.'"�AX��B���g3.�ԙͿh�4n�����9�=���.U�M�07$�~�-pȣ�̳W���!uS�0zGه~��^��-��k�3�-@Õ������p��zWƷ��������'z��ا�L\���Թ]�D��՚���v{\�Vf O��l1z��>=T�(<��ԌU�*�٢f�R,�w9mt�]�Ym�km��oL�{�4��q�Ɛ��C'��rr��0{��NA�2�ع�8�̏vdN�Q��X*,�7��P[u�OZ�])L�>�����MK-z�z��7/���%O��;�Eϙ| ��錈c����X��a�����N`�h!E��r%�ęi7�!uR��9�{��k�Ui���Ӥ�1�fB�1K�f:�V�<=��J>��O����TXp���٘.v��S��P*'L/���Z��^�Q���"��J�Ę2�]����y��a�r���Fa�SD��7�7x�����{B�����<�Gv~�\:�sv�2�f�������Z�P�ۺ�&q2�DǕ��h#���Ǘ�:s�/�L�D��f�qO���Dk"�y�ԧ�أe�h���ǃ{j5���e�>G>&������q(��2����ǽ�O�M�sb��O��Y?YW/�}���Z���A��A�VTe[^��=�[��7Ad̨�.�/{��c4��K�I�|�TM��`�%׾t�*-}���c�����J�N�_/���haU(P���cu�&�(g�ߴ��|�2�3�1=��6Y�9����̊���p���F��&�b���x���N.�.*�J� ��Y�&,��W9�*�B�S���:Lx�d�R��3}DUT����Ҟr�4����e}����E���]MEh@%u���� ԙjǦ0�L{sf��\-�����#2r~�5WQ[�l���2K=åQ0cC�L�����s�°�.��2��e��	�1>����\Ϥ��֢qrpZu*�5e�c`n�Ӗ(�fm��{�'�GХUz��q:�"��ކ� ��Wp�O��d"���S��`�����J�:��ϖz�m���՛��/�<�Y�p{O�Sxc���f�ܑ&���B
*{u@�ntˁB	Z+8�[�ؼ*�_+SH�UC׮�N�0?�.��*)9��oY��N�N��@:���Cq��qX�&�]����V]����p
'8Y�&2\����N
��2�sӝzȒ��.��	�kB���7�ݬ�v��s1Z�+�*�k�;6����W�Q�5���B��j��a���ފ����ؑ{�.��î�ƨ���{��=B-�fn�D��:�ɗ�*+{0R}���&Xع�xP,ܣZY��+)g\��|��p:�,�םxufɎ�X��=�I�$�K��&&E'7呵2\L�F�hba�,��[ԤطC����'��Əe�"�7z�]΂ѫ��>�bb��=�����I?vSŠ=ɶ%@,ƪ�fQ��!��jr]�X��L��ז*a��la\�g �1!���j���G��s���*f��Db���C�i��n�jdPK��TCL1IQ鵗�l�.t)ݷ��x��sE�3VV�=ӹ�:Y��ִ~�.�%�K��UtWlX�קN�9��b���/��2��e����7u(��a];��Y$�t3l�X4�J�N5��S���������U��6mk{"�d8��uˏh��ҹ���o����if;S�ӓ��fų�A�P�h���Aī����u�z{'j�� �T�5�(�"���v�w�2\V�wui�&��meKy����f�wA��e���إ�z5�J-������3}a����]��cG9��w~T��NV�7yer�M��r�l
�B��u�
Й��۳�v�Ӣ��dA���X"Cy���")�ϥ�3/z�e�H��ӗ��s��uZ�F�QX��s/65�\(�B(�F�畒f���1�:�*]�,K�V�J�×[PX���/²[�Rۼw���ωp�e5���\H�Xgj��_i���Q�Ky�ٹ\4�6�c�,tsM<*�6��l��-:J�X����=MM%R�W�fN��޲j�f;2:Z- ��T
'��[�5@\=-v����[.�t��U�Զ3"њ)��[���t哺�6$��I�3Ua��o�ڲ=���ʹ���$�ǰ�Ӊp�[��Q4=��*=��1���hNXn�=n�xW���/�^&��Ŋ��x�o��9�5���j�w����w���X4a\9*3anY��:�QCA$c��.�9�1@p��m2I���}�N�/����k��P�jTX�^t�a�*���N��K��;��=h}]ډ��J��5kB����Zx�\�o�%���ՙJ[�F�vA�X兠�Y
w�9],4� l'R����Ln��@4����h�����a��d�mx*r�K���&ҵ��=��f��X��+�A@�۞�{܉��(^��i����+�3/�:`�w��;w���k�{!.nM�.\�H�I�R(\��-��U�f��z*8��Ԯ�yjDsY)ЭvE�����z�8�M��S�W�Ās�p���VT�<~����؆�����׍��+f��]J̻Վ�6嘆},��ɽ�-��ȹ.�;�����oP�Yռ9W:�;�/�9������嶨�ޕ���)xr�]�/l��8/�Q����*��m���)���OL�&�������;���&LvKvM	mY�q�T�t�B.�=�;�ǎ��1h��y&��5hY����;��d���m=�ڼ��>;�~�#�V]���/����a�b�K���SYˁo�#;�B7��HIP6+>��'D�XR�׾VyG�ϖdÉ����@c�ҥ2�3�8~�e+|'����*{�y�૏&�|]���%5�P�?LNܬ�%��ǜ��c�ve��	���^05R�{��I"�bm��ɢ���M�����[����R���*A��y�����:)�UM���O�{�x{�Ǣl����ݔ�Jܾ��[�⣂C!�sw�+=�qw�_�cy������WF�aU��o� {�21A��uP=�{�5Ǣd=w{Ӹ������;EP&=yB�_u��ugE�X1z�_�����G�����.�*Q�4wk���5t�#EN&5����{�vd3'4��W8���k�������b�-v#��Loh/��^�������Ê*h��tn-���t�&�X��/���Y7h�� �IJ̃t�E:�5��e��+���xƪ�F'J�F�.�;;���oS�(����B�W�o$,m�u�[(�h�J��{��ӭS��[xnHL"y�W`e��FEa2P«S#%l������98�����U�sm
W/�o���>ȗ���'�㷛��Ce�F;�� 󡸛��c���=�SlB�P�g �S�H���ټ����6���tF�o{�w�}�vhv����D����7����#��((�U�|���1u��U�9G��=��|L�_3q��H�{�Y�4����3/�o4�R�
�Y��B�y֎º^��\� ��{τ��\�ˊ���tf*�y������9/�';���S�"�N�𩻼�q�'�EB�i���6席N�q����L�m���S���ۢ���rug����M�����"�u��?�7��*,S�ĕ�B�u�����E_��_�B}�;� z�[���q��r6MU����Fm�{8��ǩ���E�������"�ʫ��w-�T�t��1�mI��r�'��g�.R�t�*�,�V��PY��UZ�F�f'`G,�mL�����FUL�B�	
l>$�L���1t�hܪ�=1 6��b7��*r��a��ɉ@q���#��	�~�8���n�ܾ�����bX�oX��ٝZʓ3��6�n�;��V~j�3S�[�66c��:���R�V7�ut�n������]2m���I�AWfT�u/�5�P�tL嘶p�ط;�/�a���A�9ip���[�1t���X��*ɷ]����8t/I��5���E��mzf�U1s{�B�������ib��b���Ta�L�����^{�ə�8�����*�j����4���
�x#Ϫ$aM����N��*7i@e��n𘩬Q���Yԇ�r�ͯu�.�<���M�����d^yJ1oTp�����Ok>4>.�̢�K�v^c���IR���d=�QYlGr�\r�~u=�T�uF�gECͺ��RX6*���F����r���3�� �����P=T�Y�z}L��34fH8i��ױ���\�� d[djw�㟘�y��c9������3NݨqA�::7��	��4�f�k���*�+�k9l��>�#��e���y�E;v�8�u��Y�z��tuMlSfy�ܲ"}���3ח�������УXM]qxk�8q6oU�c��^W��g
*4���ؕ���9�Gi_��l�߂���"m�3��eCaj�TE+�� v<��'�]0�z��@=�f������q��Yب���~g�|&�LƬ���)�� d�^��6-�`n��gC�A�A����Cd�4W��G=l��ə��k5^n�0��َ��bkp�S��h�^n-$�h��y�6��aְ/������"���`��F3�A�Uu�E9Y�r�2���4���)���#�79��B���ptK3N����ҚWLCZ���m�J�j=�3w9ˬ���q��#C��|o�������\zTƚ���~�x}�0So`,��"�_$9nT����x9�H��Oz��ҹ��=tD81c�w�}}E�N��5y���L�(��;�	w�7MS.�l-�v����$tV�.$�]Hw����j%��g7�÷���ʤ\�ʅ�gQ�Y��߼����V�����~��W^�ٷ���1Ub���uU�6�ή��ޞ���w�����o ��Փ^Ι*MX���@X��+l��·:D2<3�}]�>�����ϴbŢ�A������|�ٚ,N�&g6�<�0ޛl�9�U�3���S����;���VAY=j$�0�_ͧF�`�?SU�^��ʼ_)>�Z]�:��>����/ONu�9U�t$�&��3�᧶;1:C����2��$6�dz�&���!x��t� gG^��v�fK�����	;�#~�)�"ǖ�P�gޜ�ǾE��I��P`j�2ٙ�-���,d�Xs�h{��^fr��a���~}�!/ET+�*:W�x�'��#��\�kܢ��=@$��L�߈����R�+�Sq�խ�J�V�|=�'�������[(ň�ҍ7�5�o �>�$���?d%ի��d�ޔ�>�[3]Ǳ����{0V�H�����w0R�3j������J`�V5TD۴ĭA�AӤn��J�љ�����i�]�	f�"��ꛠL�Ν����G�&Y�/�uu-�H߅�٩�C��K����6&�
q�����T�	�ð��l"~�&��:$A��]��;��Rx��!��p�ex_h�3�룵�ڀ�UΊ֣��S����ǵ�>&�|��+oD�T�[ U�=�S�����]���i%�"z��53x�����ss3��ق���J��j���9�w�$�u�Y�O2
�*�?XX0��JMx���	r��@�\�(��eǻ�·�}�X��e��4jLi��}=�)X�2sf�Q8UYx����Yp~�״c��w������R�w��>Frz��l�]ԫj�"bz/_wj��D�9g�X�N4uH�Tw<�����j���h��c��!(y�y5�$A�:�Zf�R&�e>]N�(��gf/�O��R��Z���"�
p�}s�\����ʴEM�(���<�)����q�Q�?8��3|�*���:��ȧX����\;�_�s4/2�9J2;8�S9�-T͹���sW�ä×P̯f.�.�д�Fi̾�s\�́f��e�N��z~���D�W�H�s�U7	Z��[�<hlJެ]�p��5�S�X0㠭�L�n��ot8�ve*�<V�CDQ�/�mX)���k��&�nU���dpVh��U�b衭䋍��r��_ �){v������i;�Me����a�����vDf9�RYI��&�xeKwF�	hR/u%5wt���G��辞����V3�)�`���E����2�=����d�?g����XO]$o/�f$����Qp粗����I��tLN���y6���Fc�9�^����u�w$k�w�fj2���y �קlJ�r61!R �=��o��Jc��4��2203�U5L��T��p/[X�L:���=�D��u�+�M*.��wV���� ws���tv{��Vk�yy؎@w�߆��}��V���!_�_zTk�fr�5\žM8�xəs��n�`�����s�QYʮM7ש3�-x��[0vb4Y:�=�;Z��CpV	�Br,>�g&��/��ܦ��]���(������퀣�8�������*h��}.�mV��~��`W�u����{�d�����5]�UF�x��%��e�~}����j�������g�(:_Z��N@�}��32;!^ с�n�C�t��Q1�ᮮ.ȟ9�f9ud�q�&f0����ʾ0o��G�2�[Ʋv|ٷC�~�if��uO��A#�8#��/fxi߸�g��7�%m�P�xj%V��b�\�{�55u��8�`��3��7õ�4Yg�+w���\���N��,p��@RT3Y��S&YQ�,����v8݇���-�V+WԊOYr���.i�&��9#Ϩ<��U�rZx�E><^؜��Ne�r��p.�(�(S��+}����BvO�2�`���rK.r�O91J#��}�۵{+GΡ��82g��X�nyO�*z��QKɮDt���9!��6����H%�O�P�ˋ�ڬ���ʦ9-��̩]p#S�C��⣧�b��^���Q����Q�B��䄝���;-E���/�$$8SQ�O+��9�V{�y��n\�ū8�&|��~�N�w�t)��p�!��u�K�V�h])Ò[����v�s~��1f`��LWf^֥�\�k8��"�����Lg�l2)}Cd�0^GS��]�uB�s����ho\��=v�E�CޏzH~1Q�s3&�rNx��>��Ɛfiهmf��^Wl4\����׿ƺ��7(-�S�db>�{\��ٓ�����>�6k�>���f���E�e$��!	f������ޣ���{�)�NM���2�H��=>v����4�`>�ư�d��s�`&�14��Bl�Uv}O����r�{m.@�v=1>�^��D�Aۥ�m��^��6��yo'�rE�C��x/�tV��&�'��f�	�Ԥ-]0��e�F� ���rVr}.M���Y
¯xxP�>���{vw��QdX�0���\9WwF�	;�C�]���)����T���0���zw6-do�3�V��rV��7L�y�-�	m
�C���BN�Y��
Y.�Kq��"5̭t��0D� ����Kf�bU��Fi4�NQ5��wo�@j��iQ�,�r������e��o�Vm�P�ߎ�=��;S�6t� V9�:e���:~��J%U8�I|5D����{��|8f��f�=���H��V�#�zvG�D<}f�4K�*vP��V�Z��h�;�@���]����@���E�Y���i�TqJ�w��3��=6&*s��ܛ�Qb旼Q�+��Q`�8�|E"�7tـ;mn\I6��yT�i���oSϥ].pU�7g�.�];����g��?9E7#ތ}6:.�Ê�
s��Z�!m���i3���lɼ����!����Q���k�V��t���\fV�]%N��0�q�d��/a/���w����'�wl���h�x���3w��_�3�ì�`�:��/t�o�Y�j��!��q�nź�c�9�2p�[�`3mEz�)YJ7��r���Q�\C�R�4���C�#���Mns�:U�t2�цNB�LJu��~]@T�/�Qm}o4��8�t�9s.�ژڏQ�mwV��1�Y@�v�z�*/���	i�U�/cP���NeS����b�&�R;j���9�*����y�Xo3d�sucf�"�z��w{��WM6ȭ�������_!�r8V��zvr΅�tG��S���Cۨa:$���Y[�/\k��]M�J��kᎋ�֋it�+
�E�2ui�q ������F��1V���sf��^�3�v��n���]��P��eB�.������35�u*Q9{F���6z-0)�O7½�7B@��-�!��K�|�ۗ{�|���G��B���Z�n��⭒���|[��H����lq����E�z�ສ��+�S�d��٧���`=C����/Ӽz� {;�8���ʺ��y4���w��g.��ωL��ר������=���/)�"oo&��u��>���I��uϊ�=��BP���j^{�n��g@��\o򪥔�0��S��ZO�́,.XN�y�k��+� ��ߔǼ��Ag�1veހ^M<��8� e̻�U��̠l�뎸��N�����������X�LN��~�ŎU+���u]��L&'Λ�,�>���8��^u݂8��}^��u3��&I��yF�R�~�o}��؞�inK�Ecu�{��V�@��Q� ����:����|��n��^f��kP���N�l�J�b=�`2�9m�������2K���y]q�2�d��j���Tu�N�� �zD����n�����s�A�@�§��d�9����c�Kk����Z���N�R��>�����dP�jz'N���N�$�q��d�µ�u��r��B���N�ծr
��St�1�`]�x �`j����/uq,n��t�\;��"��+�J�A�8*�dq��+���?m�V.�JvCc6e�֫��Ra�(vb�����J0t��<������K�CV���B����l�*��`ߣ�
���)X��7�ih���7_��]�N)�]z���o�-^�z)�	n�nc!�}f�~2[�T
鎝u���G�� �zDX7.�B�&�^��zf�,dk�|�!},ɮ�9��q�Nh$���9��ߍs]�G��c1B��O)���<�/�KI�W51�:����蠾Z�y���(h��,m�Fv���aL/x�¬]�k=�תd�X�r�Od�]�`zn燨ɇj�u�+B=Q;�:��+/�ᛴ�s۷\�O=.�F����%
Q���M��k�,e߹�Q�v���C�N�E>\��}�=��W�l��P��$�&\n�;�ʘF��WF�OE{3������}{e���D˂ߖ\�3W��5=��KI�1�$�~�}Eւ�m��_ .{;2
2#7)�E�Q��գ��)ݹ�"��K9�C����j8]�˜�sE�^&&4�Q�u{&��R�T��D�ݫ���~�8��f�9Ef泷l}��:��5�x�4'�ojVl��R��d�=��9��{�i�-�z�r�b� �G�Ө��Ǌq�й@Q�g��3dƗsXī����pu��`�g�]�}҅)������
����5Q��[��e�g^�V;"6n���_��Vk7(��������QH)�����1W�z"UsZ0�U]��b6I ����O̑� '���sT2�����{=�\^���z�L`¯�}�gu��9��{ns/Ơ���h�"�۝nWd"��p�~�W���wz) �i;�}鬬�w~�*�	8��a=�}�3{;�{;� ��6���j�t6�mݕ'<�PK��Ѝ�n4J0l���#;��0�0XB0}�]5`�VF(*d9p���i�'P&��o�}�ǈ?�`m$7���~ѳ���D*w][�-)9́/�.����[14��w����7Q%��VF�b�nJP �C,G��8�[T�ɶo��3GwGGo�$}D���ò]��Tq�ƴU�	��qD'p�6�,�M��t�y�s315�����\^R�WwSh��Pc6q�JJ���9�Ah�QgT��ݾѻ��@Y!��g/0� i������=����o�l���c	� ��:�N�I���v������BS#f>��.��o	aB��	���5�JP��1*�n��E�F5��+�7��l܆L�7���)�����kol��źc�Jea��0����p�5ZW\���r�%��_}���(�4��>��cf3Ta���`b�2*MH�!$"i��6�:f��1>�k�CN�ff�L���[�]�����'sv��5Q�x��ֺ�[��ޭ��qd��L����[�d� BFň�j4�`�.��Q$�����[ ���K2���/���w��k�n��YL��OO5�R��V\'��Y�@
$}	��G7�gD`�i&cD�B$h
h�����f��`�b1�n�#�~�"�����i��	S�w*V�}�P���^���w$3����k
��p�Y9�UUY�/{a��ő��Xpu܌���ԭ��l��t���b^����F�w3R�Q�UNm��x�ɸ��|0�[�5^\-u��:�5�F���}�ڂ�*Qs��KBQv�%��8�1���h��Y���z�A}!؝$$\V=�Bэ���t��X����ڌvq_���'�;ALΔ���l�V���~㴹՘;s����:��^,3w/L�1ܰ��h��������{z���{��v��R���e��w���]6AU�;l��X
�A#B5�[���q ��A�ch��o�.���u �l�f���WU�M���%����&��ժnSK���_7���ݹ�#�S��B���lsѲ���,�n��,/hv_� �j̫���79��W"(p�mH����)f�9w�&��m�X�T���""���Q��uu�����A�p��,�u��f�>o��fd����=�gj�a�l�Pv,wu.���;R�ݕ��7��iV�̀q0���A9,j���*f�k<qnw\[@��7�n�޼�Q��x����bKśp!%-�ҊJKkrn�u%(��u��9aW�uɵ�ᩅ��늤�{��ۖn���	7�2�;Yى��YC�u����L�[�m�!��@�8�����m;)�o�h�Ӱ��zi=u����5D��w����1�Y6�T�}�dg��n�A��Xɹ`��~���US���zU"^A�Au��Twz>ʳ��2���e櫜��3
��j��	��������ӧz��\�����=Y���C��8I+c�W����UieZ��`%ŋ7��;�5����� ��cr��=Y��}NH��ULvV�,���T��p�
���)?~s��':}g�V���"<y�E���[T��z�fO�@'��i�=
Ɏ��O�.dN��fuA}W��r�t���� {��z(>`���q���U]^ȕM��U��q~�E���2���;�U;�T)�^�D>���8�єvr�oěD���z����թAհ�{YX��G��P��qw�+W��5P�IÍ����J�ی��TS|(�5#�4o��+q8���q�o�t����s�.��f*kl��P�f�Ú�������C>�Ws.x hC��:�2�^0"�G�����t%��A��toK�����Q��H�8�30�ݬ�O��ў6�q�f����vde�L�3�|�o��b��������ͫ`߱����©OϦ�����S
-�D*>>���b��*w産������`�D������,q����C�R{�c}Qf��Y�]>Ms�ezNf1�����kB�I�8a��n|�U���݂�Cy��&Ëh��ßQz�s�R1;�@5����E��@������5*�X\x�1\��h���N~��rf�=��_Nl��V�=���,�J���ժo��ۍ��'n�{�K��9��9s�9����R�|s�p��B�z�fE������;W^q˳კW���p}��WM�3�,>E����=�]~�Ur0Ǽ�P�bwx����iR���DG�_f��T��~�؂$fŬ��tTKf�D���&���l^�**���=J\����^{��*[���@�m��]Ѱ(�N�G�1P7&W���x\��E�x�,&3�e��%�i3D��^� �yQ�C3�����d���=k�{����\r){��x�T�T��F�I'^/S��\=���
�ѳo�F.�,��5����1��Xyv���'c�4�
��]�u�YP�@��,i�/��tn:�Gn�~�R��y�7I���r�:#$E�</�OA��쯾`�ҏ���F�!�,��Ō=rsu}ck���\q�B.��d��G�0�6�.�wOz]�p}P:sO9Y��}����ڍ��(�Z�p�~����~�/oG�Ȇ}wE�{�%��w�GT	�����R'�8�T�)Go��l�{�X�!%[���r���6����w����d�<�˲�։�$ι��`݆�+�qU7w&^��Ǝ���Lѽ�իS�����+(@�Y
�P��&V/��H϶�r�^�ڹϯ51��D���a�D\]����J�]h�Y�\%_<�C/�{$��u��Y��Z6���k�p��ɣ��3 P�t�2k*��wK%P|ߧ��5n�-iJ~���B�ǖ�C�q��b��0=|j*����l퐪N��+���
��ht����^�8*�Ke�Γ:&��w��Ϲ?p��Wɇ/�e�s�s!o2���b��B���	w�D/&����@xN��
�-̧6�A@]Iȑ�F�;}�2�j/a�լ�ᅠ.�7����{=��~�9�����"��F�ķ$@Q*0��Dy�5�>�j�mm�>Q��gL'i	�a���u+Վ���5
�s/�iǕ�>��jO���O�`���b���`�]�l�؛��}S_5�G���/21%Ҵ��F�p�3��176Ǻ=�q��Au4ZAg�����m�D��y'O�=RV����-5_�S��\m��.���ͫ�$��NA�8���ނ�B<7n�����*7i�w��y�]��U=j�k8J�Z�J�9=��o4W>8t����5ˠj0�*��tRVX���#f�*ly�>�2��s���)?�Lhb���a��)ܯd���]�Fľ3.n|����3����x<��qwm5FyA�`�^��ܰ&�p�]�n����� ��ԙ�{7.@I�J5-�w5��sE�uv�=�+��9v�ol�|^��W`.�cXKz����g:�3�D��k�L��ݶw�X޶�Xq���l	���M�[aX&�><hi&.c%�1���ڤ���/:��ƠA8�Fj�p*m��ޯK@Ÿ��@�sљ���uKpO���Z8���W�����&��q������]�CeH�T`EU;4xU���k�l��m�O'H�S;�t�E{�{��������@�2Z�;��4�
̫yN&랎L����$�H����ҟY�s9N �kv��S���R5�=+��4\Z�y}�8ՙ��u��)oӪ\��^��o���B�Ή=�Z1�`�����P���p~��S�u	�/�"�V� ��xv�iI����������Y?q5~vWUÇ��t+�Vm����rK����W]]�AQ=���S4ڬ3����o�4�-��%>���is��싼�^�E�]7�<��T��k:v�1�:tG{4;�?%P���(=P��t\P�7��sf�u�G6j8S��M��oذV[s�ҹ�}_���>��k�6;ob��wq���K�2�x��Zn�1�8[V��(��+�|ש�S">��z*���.���},�푥�ˣ��%Td)V�^eHNQ���by���s�V�ܠ��P�-!�wNӖԬ��c7�%���uK*��Ф7�h<�4ުko����[Z�:��JB�WZY�J���s�Z��*�we]���fB����sp���-� ���N��C����5�����1x*��՗zڇ;X�m�U;W>��mO�;�&1����2�>ߏ�^o���p�Z���ۏ����1�#|4[���̙�˨���`#��{^��o(��k�댟�~k��&�c��-F��>k9BQp
��{���d2.��k9�����kOlˑ��KtR�z���b�Ly4�{|�š���̧]^�^@��vX�ko2f/��1✆��дd�ܼ��ذF���G�5���	��:��8�6��H;�ϫM+����T�{�	s<|�I:3[q^=*�J�����8ܝ-�@���cl�}O��<wc���j����තxS q��kn%�'v�U+Vہ7+�:+�]�Q��
��Q`��A{rc����spQZ�ζc�xL �&�g�%w-�\�@>��|U���	쳉����n���!Q�{T�1(L�C�+��r ���M{:� f=TK�׮�g�K����6b�@�u��$��9f�"9�jQ0c�r�Ga����}���0��h��|
�퉺�Ӕ규+Z�\�O���K��f��������н��G�E�,]J���&,�r�]b,���u���oGu*@�a�2�Vk��yՆ��L�D���!�@,s-jhA�a�I�_^ B�9AG�����jN�����44��=ݩᔭ���4f�\[��A��͂_�6��r���j�{=�%�UJ��h_\c�"Q�}H���K�FKXǧ}Lg\Lx07N�|��S,^��:���E�/Gzd(�ǣ537��;�N�ʗɟ�v���,�`͊f���8m�!F���h][�ͭ��S�s�k��\��*{���	�� ���w;��O�-��9ަ�	R��vT�ڿT���9=3�7�w�ij;�G}�c�o��4Q�t-�49����۪x�5]NLס�r����8��`UGY�Sf�ճ����z4v���pv�>�d��~��ꚪ��Jr,�ۋEA�ނk�W׽ݞ�x�R>�Lq,R�{��-�y8âe�r+�����oR��p�ęHU^>#�3��Љ�ܣ��e5S�f(�Hɮ ��U��W?U�}��X�3f$�/���C�w7�{�y�:�\V� m�"j�ѥ�nk.O?�]�m�r�xfx�1�UzWh�wޚ���ާv���� Q���\e+$@+4U`���x�v�L;�&h�ѧƴy5��]8�/UZ�Ƕ���4���8*�M���Q8�+�@t*�����K���њ*���.������S[Ai���	2�g^�������|��zz^� ��R�XηNm��j�Y�����䅇��4��N�Ù��H8qX(����,�+�ò���1�u���>`S�vAW}8V%e,�*�|������s��N��`wX�EQ��e�z5:7���b�j�8���*�{=�k�
]�V׊4ˬTne�*��Rv�k�yn;ǧ��ؒy{��?O	��p��Gs�Y�.&����Xcճ��a��S�'P��UV�Șy�&�o5���Q���q�\��zuf*��v �垺9{N��~ꇶ0��\ʈ�0�Ud���nS��u�dt�K�V�A0y��5j"��@ț9������)����4e��x��}oy��%N������R�r�J�$��@N||�K�_r�n��z��U��هJ���:�����Q��S�;,{�<n;��y��J<-Y����I���G��9j�YXe=�qC�u�{,<ut��W?r��11��OBn8v9��ͯ@�C`��Z�8��/w��bK�@��4�ۗV�M�w������c+U'L�1}�|����+7��Jlx\�Q�i*����2Ѵn�[���B�x�iRO�т�ي�)C��湄Fß�=�<�{�F�.F�������yA�^�6*B0�$fl��{&�@��%��T������Ҩ��X�G��#��+L�{���4e[E2zMʜ�"��m��ę�P�1�M�@�K-����4��m�f��L�;�mPQs��". Gb�N��,\��{ᵖ����sq��Y������C�x`�iBq�mc���"��Q�^V�U��o��踩���$�wӑX�����B���w5p"�۸���]�:	n��j;~��f�0$ݬ.5�ve���
�Z��1���х�̬멝���z��OT�������\(�2�8"B�p�Mݠ��_���}F���;� �f��}~��G���]]��c�|f"ť皎t�Q	�~�5�\�tꯌLd�:�;�~�����qv�g���y=���x)G���Df��ʷ�q��h�V�Ɋ͋���ܠ�d��~�Π4bn������	Y��Ǟ���`�鵫�|+�p��Of���K����ڝ�7[��Z Z��!��H���X6�sG	Y[bCS�ܺ`��:���DƇ����E
�m{�j��pBZm���}�����Tf��Z�"xHu��*F?g���-��vky���"E�\�cِ�\$�J)\���?NE��مa+���5�m�����3������{D�W}3Yor:�2�yM���n:d^3�"M	A�T���ե>�<t*��0ai�����D�7�C��J���@�����}a�����|.�
�@�+*ʫ�\��)˴,�{v���4�h�f���Ձ����e�R;��j"��L�xu�X]�&vy��I�1��s��RR����wj��R]��×ڛ�fx87g.:�<�u�.r��:��N-Z��s�d�`��ș��A�ͨ�,B
��)�uv�]�~��xT��^��Q�Pv�~���W1vb��*��>��H[�[�%�r�ܪӰ��J��*��Dc�טr/�X��z$��-���W�<ԇݦ�_�%�϶
��VI�7N�D�bqW>T�2{�Y�L��8��<�'���n*�eh�pu*�p<�/��B�t��ee�\,GUL��<�9�����e�yv�^����9����Q4(e�µ�5�tx��V	��gXBk'���,-gF<��_������2�dsb�_B��9��	P���m4t�S*[ױ��A5p�B�7���\yog�٧��)�Ǧ���8���}��N	!�3��23�ç<gh�����]UYu��JU2X��"��9�*�:c��tT�^c���*X�E�&�a�~�2<c�U�=^|+ ����U&j9{���C!g�u���.~<�n�'¶�Z=I]E���X�&�i��bYf6dc6.�o���e��ט�/x����1GG���'�jp��v��S1��sA�>��`� ��tO�XV^���o/uUF\���%շ�Z�U��������h��Īp��D-��w,��ymK�;	�4 QJҖ�iX�@��X�^�],�Y���8H������6��☳��������t�u��+�Ep�����v�ex14>a�rt��Qg�<�*,<���d�Qp:��*Me��b��3�{��\��8���I���0 �縃�T{(��΍E�{�/��.�(7p��u��xtL���&�N�h��}}�q��i��D*�Sy�cm�b"�)����]#�J�q�Rƾe3NƏ��\<��a��}�Zm�8/®���0�/�o�P�ݝ��m_�'$x�U��T�ﳧ��&iT:�ET,���Y3ΐ�^9,;:~x�i=��9p��s˨��o�>	�k�X����(�b�Ț�n��A���e�p{2�v:}�pf�� ��=�l�/�1�{���53m8�6��|�ۗU��t/�������I���7��f�\�I��r��{�&��_�h�ߎ~�j�UPS'ʽ:�
�p��������j���BL��aG�u����S�T+)�^`� �1�X�|#�CT�x�н2 ��U�L�T<�qGi��P�x�t�M.�T��j
�_�bk�}nܳPL��x��]�&�\�R��$�SX��^Z���Q�K�`*�>�����w�sԕ��GS�0V#qӾ���WW+/��M�r��;�b�$%������q��h�f����Ი� �\�ym��iVf�����Ti؛�h��Rvv�p���ѦW
��tZ؏)��K����fyD�%���؜_l=��oyXon�����Hv��y�$� ��n���}��z��]}�����܆��!���#+wc&Ω8����}��lJr��C:�UF��,�V�3�b��߹UY� M0���l�o\�����o4��_RS��E�X!Td���Hu;���mAX��J�b�a�Hp��q�1n5Jji6�}X���S��������	I$��=@ad���h���k�I�W֮ r>���˱o�rV��,�2����uFD��oH9۝ߞ��I;E��\��*�Vj�9���Lj��$ �v5�xz��;�UG�n�n�(�_Vz����eoo>�Lê:�JY�Y(�}G^��[}��a*�����V:�0^��-�.u���i���t)�Qx�u��n3r�0�Ǭ����b""&LDE8iBOw�i��K9�m@�3�YpZ3�Bu��Q�{��k=~�7P1��몯h���p��FG��%�_�GS�okpu���/g9Gw��m�v-��[���ZyAA��/f
�C�҂U1X�	YU9��Y�{�ﲯ7��d�	 u�g�z���Xm���u�o(�S��JLJ���.���!�׎a���ԭr�0{Fk�箽B�stu�Ů]ִߴ�kwB���5�����
���ذݩ�?)U��bMԪuT3Z��#\Iov�k� W�R�^T����vq}ӲA�����(�كD�|��*�\��ˀn������N��X��r('GՇ��Ư�%�e�i �.��lK�"��)t���U��/.��j�M��%�Ț��j�I��i���|wwFs��Րa-���}xm�+9}��.��%s2Ct�yM,9W��ʧ~�bl��%JܵF"HZ{�Ie���jv�*;.�ot��k�e;��X��ܶv��������K�N�buϐ���]`��c�%�<��g3�$��Sb	�˾��F���ZE���V��x#cYr"˽�qF�y�J�������,�T��5�6�u]�*�;��Z��أ��7{�Z�W��]"�4������9����b�BL6� ��h٨�T�+sP����o����Lfn�䖢j� �Lv�Z=C�u��7��V,��������(��Gy�!fY��\9�����ֶ�n�N}R�,�C�]��I��i��L�7k7rJ%�D�m�m�7��x�a��at�Ф�Κ����������R���tfn�4C3��j�bZ_fp`�;-ե�eZծ�e����y{����=%�][v]�|9ӾI���:9����:��t�!��:>y�<��m��%^V�M'�0	��vY��Rv�d�RB��(>ˤbꋬ���nꖮ��s�d�t�\4T�ôճ��EBd.��%+y��l�;���45bU9�I��n�E�-t��k)*mK�yg:���7+����x�(�s��*�P��돆eL���ri�V�]ֳRJ/�:YyՄ^�.=ѽ[��^�V��'5�}�+.��Y�I#vf��V�`�E��tV�߱�������9i�0U���j���f�;�HO^��uen�i
�e�UͮR�3֫dn�R��N�a�b4����n��sL�Z'����MB�YƬwe<=Ή�����Y[�L-C+/�) �af��2	�mm`�����*H�$(}��R���NVq�f�A�S�=����~Q�7Ce|/�@sG4�S��ط�[���*Gz㑙=�b�w7��Jp��`����c'��[ami�^�̋b	;��O#`�_UFg<݇'�؜!`�hb�y&�\ߧ����|_�/s��:k}��}�ky�X�}�/:qћ��.��v(Ɠ1�u�t	��N=x�l%V���9��RL.����|�e��xd>���5�Y{����H��G����~i�[1w|C�us�1�a��^��B�K���l���`ҊQ4{e �볲�f88���4C�O��츰n,�bÉ*YԀ�<<�=�v�Mxle/f�L0(�q\m.�Q���#����
r� ��n*)
;1�jG�<~�	u�]==-9�3':4O^gT"�A���o�c�Y�*y%�0��z��g+e���Oq�}�w.2�x�˃�c��9:���?=Mq��*�uqQ}O��|�>Z��6��s\,vΊ�u]�:������5�4�{��t|���\����r�_��si�U�T�˾��A*�.�	�^�b4�{y,Z�$�����T��k[�Ew�i�݋�]{s5˿�ғQc�n:���{g�N��$o<Զ����N�)�`��;rw#� �Ɨ��Q���7��ꉃ���"D;��60��ħXѭ��w�d��ڴ<��&�������	����V�'��[�bž
��Y�[���h�P�͇�&ꢌ�#�#%��n1h�6W�1kFz�=m����ѓs�R*���I������M���3��U�	��`�׵���n^|�]X����2���rL�K����,�#�>큓eh5���ߠF�>��w����2��o>��R��w��v��aN�&�=�Vj�����Q;~���裵����p<�w�c,�]��}�}v���̉��B�*�����L,lڵ�&jq4#��b=��]n�֒ņ�n�����`��I|v���ޞ@��>u��\<`�Yr ᤹���N��^�]¾�@b��g��f�f���d���}��Ц�ı����`X�N�cܬ��z0�a�����Y�����S�8�:8D�8�re��ω~P�'�3Ӈ��{�<㇏�t�m�Ͻٜ�)V:;�h��[��΅�{H������Hc�Tα����C�M���f���b��SA�af�	n��ۚU�c���m���l��Y��!�oX��L��߄Zn��Y��U��^�헺�pm,į�+���U���vѼ44��}�r��Z�
�̼�u�^��M��	FiTU�z��E���K}���ڎ��>w�̗�.�p����iF�{s#�z�往m�
�� U	L=p�ؾ���[��	f������y^<��*W'��oE"}@PEo�`�f%Fک�^)��	�#�;g}�{�����_A�up���8��YD@��}�� �n�
(<�OAB4_P�C�I5���g^��F1���q���Ys����C��Yܻ k�5d�����|�B�]�N���Ѓ�h��;����^����_Vz�9������\c"�JZ�R��i=��4��k�ȸ��WGM(��f���=��7R앀o0z)M�vTuvYY��{]3�q.�]����<B�������(֧���Ԃ.���vE��A�=�B��4��J��2�-Qc'����ݾӓ��WW���DL�E�f^F�W�P#�����#��F��7}Jj�t�*��}����H����Y��u���v�]�%\��|�yQa��B��;��>����x�|��Q`�B;:�.�	˘n�}
�5.:�v��6��K����y�.�}j�\ͅ1K���)K�8�-Ւ��.bĪE-�s�2nc U����R��w_�)��c��y�u�V�_C�C�8Ŵ�z)E�b��ӋE�&���	eFCT�31�!�բ�=�-�(��c�{�����.�-���luiY��¥��O�������OIk�aL�r�����x���Is@���EEe)!��	�S�aPw���X�8�-W<�����;��j��C`,�O7�b���ǲ��p�VU��*���J���~��S�k�L_�i��e�SMS.��b���5zY^��彷�&}!MJ:�}��;ݮ{�0��q2�N��6GA�Ω�Dߢ�_��CՋ3���!���)a:}���i5.����s���:~�}��5�����]]��l�۝�/���X�g=gs6�r�k=0bk({�1�p&��kߑ@j4� �i�Ós�b��y�sq�ug�zQ��S��p_Ռ֓�6��V���L{,��"Ч��;��^}��D��Vr}Ӣ�B�*��"�bI����P������3~O���K�{��;����+R���ȰuK��OgnYK���L�de;�QcBYϦ��8z�4�ϻ��xz�1�Zb���tL��d�uj7I��v�(�c�:�:'#X��/Kt�U�dd�/A'�f0�U+zl'��Yk2;���QɋJ�}�����_0�m��W�qi-�������c���m&�58��)�s��шf;K�0�����Tk�=�=�t�J��7x�tVP��L���L��fufm��~���������K+&+�'�,L�tk�V�T�q�7�I���rѮ���	QfS<�5P�.gn��yp/��JWa�s�'�F]�}�
��]�0hl#��v纭x,6O�����Y����JK��죎	�g��c�>=�	��U?]�l|E�#�����-=�w=���;�g��s#��p��}g1f��őj3F���ؒ��Qos6�kxS��2�9Uu�;:}�XA��F�}"1�Ӂ��%n��Ui5;��S	U���B������+Sl�|�S]`�׶k���w(q�.|)�z;����=E�I�"��� uz��Ց^��e@����&�{���n��E��۰n(`��4�@�о}${� ڋ��=8tT� ����ta��+'ǝїtI��^C_!�*�u�riz�燎�Q=�L�+�9t�x��3&n�
���.l�\�@�Vp�3�d��x=Ŷ�f8�|�P�a
��Lʚ㽓�b��]�ԴD��;����͓it�^��-F`jsΦ�tCa��}֢nh�Д\��\f�bdK�zhѓ���2"�'ެ�l�(A!���X~�P�v?(�|vX}F������p��(�D���M¾ov���5zQ��5�3�C����/7eKYʯ&s�^7i3l�El͸	x��nR^���zd�*�#^X��2���pCyP�����%�U����2��w��=�m܊��y���4:B]$�u�z�YqT��XA��9$���������;�ߩ���+C{r�&�fº�HE�c���U3Yn7pT,��]���ǡ��lҺ�&�E�'�_��k2b^�7Gf�O�bѠ^2�^��5f�b�N:G�{[5u��iخ_+�vs���@��i�<������(�y�
ӣ>�o|�ʼ��&�X3<�u�oޭw`GJ��X`N��P���S�kУ��5szme�̐8Q��^;�iJ�{�o2��ݱ�ټ�Txd
:�,�6/n�Z��H�0�w�k����R�>}��ʲ�̝'/̅��ե����C�8��2]#����s�6�30�1˺�}s��J>���`S�S�.�{�d��s��v9�~����s���O*����!�h*�igl��h���u汼S~��z﬩�r����<���U͊� �y'��X�O� ���V�����n~~._�s/Cs���(#J�t��C�{��r���4���|=Wu>S1G���k�D8f��T�.}+0գ���~�nc��rD���f����3�-�V���輺���	n�w�brU����k~W�!+�(�����3�-�@L��,fem:�1�#@��țI=+Ty�l��6�T�K��o���\ɫxU��
�m:�R��vU��x.��`�+��jqLE�D͠�NdN��,�i̧BF[*���32��\t�9�b8�\/�l�>���@ܽԾ.����%�n�g��1��<�S����"�g�-d���s����t�}�!�	��<�G�F�A�Ug�s���Jp�#��L�rs9��%b}G�׸cͣ�`�n��ED���Yy4�wi�A�i��csn%�r\;5�X��u�Q�r�ӥ�[���8V��e�ѐ1rًʇJc�;�;'�1�=2�!^�T`�� ��.��7N���Q��#<C���
���R'�RFOI�<�(1.-��6@Y��\P��@n.�'G�lW���/�4��(B�Y���3��4���>�s�����CAY���*<�3�pyrl�7���?7���ȇA�+��`:1Y+�a���j�l��tm8��M�/ec�UP�5����~�#.OW:j���գˣ%KG�0z4�5�*��\���"\^�U��?�}��zCsl|,�;.�L�e�Ǝ�ud\F^�
�y�
�0+�LuH�&uTc�B���k�*(�����X{(b��w�g�{#����d��Z��d]G�#��(']����NJ�R餴��"��>3��Pʚ~�]�U�թ��m��]��wв�v����.��|��a�����ϫ�!G�����:�$^��fVc��n���\�@�w' @�4��7����8�]Q�LS��i�x�.��z'+�.��������I��<�h��])���K�o5c��8]�vb�&$��jh{
s�A�!-�OP�����w]I+5�+^���A��5v�n��ζ������ʫ[�aF����L�:TaZUO�y�Uo`u�D�칫����o&'�.������R�W�5G�T�'�����'��unt�"�y8��������G;�Y���3$ްz��_swG�N��[�±�}��l(0r����T��p�L�1�n��$[�6z�
�ՓɳP�B���6{�;�Z/�l��TNv���ʄ����VFEI�r�Y{ˠ��d+{�H�H�@ �Q��"�6ﯲ,�$��0�r�bl��@�k���ԴVd�=�M����uMqy�m�MF؁+ Z�Vz}�3���aeR�ͭ��U�+H��Sw9J;���;����}�wcQ���z_!EB���}�6"�B�hc���qf�+ [G�Q[��0��;��s�J�X6�J�Wǁ�c�t�h�qYj�Ǡ\��	x@V����fTvr�����jݺ+%O�����f9H��Xr��s!FA��et��p=/�j&:QU5輘�B�y���m�!��T�i�*0M�l��FL�zoՠ"�	��ػ�uH��[v�X6���b�eh���u#Cw5���k�ʏ:��Ĭ�>�l@2�:����JWʳ�a�ԅ`ۚ�Q)���Ѻ2��!�N�Ĳn���t¸k���<�Eluڬx�PK.���ފL�1��3؊�����Tt^�#���y�����u��?h�>FW)�@��#��}�<�p�G�휊:�e��(���1;V3���]�(N�fȣ�����{�� Wݰ�K���8���L�mNO���6r�6`
�_�����>}�����DV�_K.O]>�f��z��W&{����bo,���t}��q�y�Ek�T��gn	�b��^��KPހ80)�#o\�봷��>CĨ�Nl
�V}v,��n��H�&�RVOzfp�����	G�_e��~��U��Ec���G�cωN�)m��!�tsͥK-�pO�d��n~=��L��i��WH`�������g5�]���v`+$�\]�q�>�W:s�,��vf=��P�M�e�X{�lM��QnS����ax&l.��Q��/g�:2���:-�F���-��U2XY�dDZ�(��Ugh����O��������m�}gǯ��{OtL�yQ�m�	�f]�\�[��	�K[f�ܫ��@�0�F�`Q�T�I|��soL���תkGF�yY��,�ю3��n�u�8�IZ��lZ�1;�sA��w;K�*󲚝8����D�Nf�ݠ�n�����D�]��5m7�Z�N����Q�8Z��6�x3)#|P(�#v�u|��m��Ҳv��x�.����Հ�y^G9�O�_9�o�/-<���V��,���;+�]���g��y	�*j/H��b�0-�2>8 �8�
P�W!du��f�g+Y��&1����Q*�w�jqPS[Ȭ�2�v��i���ƟM^�x;�|���4'�lbtl�$���o1v�D��dj�ϯi�Ԏ�'�,�%��ߌ*��s�q�4Ic�^鍗.9?�ⴺ����`WO	��N�td�*����	d ,p{K|�&F����D��a�Ω��N��T��Uu9��9���G��F�F���ȹP22��@L������w��v|~��k{[�:�+L�%��r�3�oA����}u��ȅ|��Y�����t���N��>�={Z��%1V��Ja��/"�Dx�~�<�Z��v�'��}��l]��ur�T���1)�T,r�40@�7./-�����Q�R4��rwB:W'2�RP��\Q�j'��[d�.b~|��2��@S5��	[���7�'
�nBtaDĕ�-Ajނ6��,�9v�\�9��2G1fU��+E��r����#�^��:kw'
t�����6�eCM
���L7C�æ��yπ]9[���T����]<�]�"�0�ZgIN���LtVoxu�깺zF-ތ��d儦�(��S׮�V�>Y���%����njm�q�uz��^��w�Z���z푮�l}�1��J/F�Љ�`'*����6�Sڝ�\؞ʝ����1��Xx֪оjJg7���5�Ʀ�yp�(!|����8��S}_�T)�r���dV3�7f7\7�[G�(�Wҹun���f��sG��Z��L%eD8�p[6�a�����w?`�t���BDv|�\B
_O�G]��eUM�A�n�`�2�X�؇('�z��Rv�u��%i[���G0T��� ��j�Ǚ۸c�̻ڬ�F.#�*������zd�dw7��O�w>ͬ���ꝣK�~͢���Bv��v�P�����J:�X�U�"���pn��iAE�	:h��YX�ŉw�PV���Q"m��4���N }���sz�q�N�;I�C2�?G��y�(DU����Ҷ��$� �� ��� Y��NS��+M#Q3H)E�OP��[O��Z��Fv���̇	�+�"�E��7R�R�[��f���{�
wt���n�g3]F�֫�l[tz�?���l�9f��+A3.+)&����W6�#(���n��	��6�Ӣ8�s\�ksB:�a�)�|oy+㋇g��>�JI����uڰ�\ˠa�`F]�9#��v�F�1W�1J��S�^�ΩWʀ�G��8p�x�t����z��7g���j[Y�Q��k�ZN7�Y3�ðh���\[2wV��k�I�c��Lf1���Ig@e���A����H��Q����
�  �ci)$`�aR������ N�wƮ��K�J ���n��V�άń�ٕ�����&1І��;�^�8������d�S�P�pdT%�9�ف���7��sH���ø�#6^{]eQᱸ7]or;w�i�2�i����o%�}Z���[-.����1��`nSq7�hW&wQ$Y�P�d�	�7�f���_vvݫm�w��2s�Lm�q�gI0.Ѩ�\T�z��
eĈ�X�ɪ��ֹJ�cz�O;)�x����ܭzy��Mى�H�zc呡El���4a N��J5
,��=�����ۡnv�6�]��su3�����K�IҾ齽X#l\�]���ƊӸ@�3R��t�7�'k.��+*C܆�X�ɼ���]@э�XN��G!٣���\�8�-0��ںڋ��_0�f��ū���o�Asu���(U���#Yw�[7`&��͔FR�.��ƍ��r+�xQ���j��j.�lq�O�4b0̰�_^\O��nV��)bf��ۅ-p�pâ�Q�t�/rq�צ���L��,��b� ����l���t���8m%��l���\
���m4r���r�+���ќ�6�C�6\\���d���'2I��[K,��\{r�*��Dar��:�ձ�l�����S2�ĩ���ۂz�F����ܝmNvr}:�Ve�v�A���ʓz����8��E���@Va����#����+�祧�hex:N:V�;#z]�ĭL�d{�7�Nz�����{]v]���o��=�ӊ��9����t���qV6cF�.�T�ǒڌ�{�L��D��ϑ�nrbӄ�Һ�ͯ`��%K_���W�,fN��Tӵjk&s�s7���V�دvL�@�h���}�6*y�����d�1���wV���3g�v�0�j���_\�<}�zs[�{�h�^�J��D�J���ĵ� �Ġ�yv��ĻS�w��=������`�z��ùB��*M38߯]Q�gy��=��7��aE:�6������K���ە�|�s�r����;q����bN��QR�����3R���*RB����=vg_W��5���[fa��M��Q�ޘ�b9��߾x�;ج�ͫ�@VX�;�=�� �tL���OFҍ��K��zc��t�>Xʆ.�V��R.�COg\���ѯ����OKf�<��#����d�#�`�_������ł�arw�Ө^I���+ί�`53�NBP���7]8�A��d��~\糚��\]$�Y��MN��sN}&<�o��rw7��hum"n�՜߯э��|*>f�̓�1�|���@M�xz�OZ/�:�;-�q��� � �#�����	^�%4��,H��C,-�_9(�77Z`�g����ܙހ;�s܂a?�M�i�����_�ec{}���u���9���7E&ub�;}|��j畸Ť��q�팃$=ۨd��aW������?��4��ٖ��G$mfu�,L#a�u��
a,5+��Q��?.�Ç��8�6Ȏ5����V��)�ٌk[_n.��Y,h�c*]n�"��zzv-:Ŝ�{U����|���%ed@A*�7�X,�5�oz�W�!x��ب�Y���ƉZ�_O��\]<����gpx�ۈ�Ue]&C�ճ���e�g�
�*0s�G"�[E;jxVH�y���t�̘WW����k��m|{!����0���ln��l���i�(GU���
P�;S�]w�ݹ�-5�ٛj}Gf��٘�Ǎ�JR.ޅ���E���t4Ӟt�+|�o�����u6����4˾Tա*����tcѭ������c���WF/{%��u8U�l�n���&�4�Ӱ5��|�N��5g	|e�#"�}��f�)��І���8>w���ǸlW�x73c��S[y�%p��� p�$���b<?ˠ&0W;9�2��@loLtq��ͳ�u[� �ٝ8<C:d�t߸ִ�Y@�t٫��rDdW��Q���ʊ<J��;g��-��R쪅k`c�(��cb΀��4�-d��b��]�t�1�th���V'Q�kj�N�N�뼠������d��W���G�k���N6m1�M�̦��}�rfI��ۛ]j�җ��\p}�?b�pIzb�-������m�����E�Ft�Ovם��l��1�nr:&����^���g7o�۴g1��!�gҲϽ��k��]ő~�/E{d�\D�[�w���6�ӂG���8:��'-ʻU3U���˺��ϧ� ���f������;����ތ����u_D�辉���{l�a�@;.�.�ٺut�H��^��L�B��m��@8f�#�D��6��z��h�v	;o�w�k��͙���<�<�Bשl�M
�
�|�իF���>^�Ӯ����m�J����<+��u��a�D���U>����p�n����]���5c*0���vuF���P���X�	=������ҫ�tc"�ƌ��.����r����\4!D��w<'��{B�WK�'�֎�,��V�\fa|1w�9�SooMu��g���Ү���q1�Σ�cmN=N��l{[.�D�*BZ�E[o��,L��c2=��Qi��������޼��P�m���l�����J��>{\i�*]Իշ�K��Q���a�NLow3��(�w�r��[I�T!0P���G��vy>�x�^���;޿~}��3�c;�#���[`T��%d��e[��� �`�����1�2ip�d��k��۸V�u��l���zڭCY|��u���F����o"��=V[i����r�A�n��K�9\�ɳ����O�F}sd�T��Q���|��R�ejV$(p��,z(�2⛝=�Qy�ٹ�"�S ��QWf�FdR�1��(*�������@���J��NV��=)Yѥ!���sQ��{ѓ2�/�1>4o�-Q��2��J/�h�n]^�n�m�
U��ݩ
��\#3�=�m`s���SR��4� E5���X{�41��x�;(��Y	��6��5!w����Evo�v�1��Uv��t=�O"��Ovq�0#î��oz�(�����|luȝ�WڥE��]L&!uR�%�1�e�@�����΀����l�[��	�鹊�=j]>j9!�ۊ�z[��
���#]�Y��F8Rܺ���ga�'�:�FǗ��ǔ4��7�g3q�U
On��oY�0�iɯR���j9cy�vL cX��Q[8�Q�+ƶ��a�|w.�5��:(b0=z��y�W�m����u;���B����+���z��x��s�"����x{T�=\�N:�Nz��p��:���-�,�'���T��o�na���:�*/Oۻ�C��2�<E��qJ��o,�ch|v��ީ� Q�+x��uw��]��]0fpĸé���4r��V��^������6�ѷZ/+ s�ųbާ��e�(0��S��(	�t�X����	'>��Hga����Zt����7R���*�V�C4���c�]K�'.p���v	ۡ3�u���D���Q���>s�[��^E;���%�#j�!/Gs�#�	��3cG ◇{o���[��)�����S�p�5��N�Ln{�ۄX�P֮�=����ֺ��m��o*2%��7eEϜ���`g
I�h�}��PV�3��K����ۧ�j�y@�+e�ث%	N�)bG@��e��q`�:���]�w�-T�����,�o4�,�rk-�)�fd@����J��JX��wɻR.yǗ��t�?5A�rg�ӎ|�Z�@��i�\�+n�%	ɞs�MA���^�I�[Q|"���]1�ri���S��	�s(f�i���8����}�v�q2@��n��C\Ź����y湳�=sq�.Ds3������oP:�e�d�SNT�����T3-LnL(�s�ߗ�F��L�	�l�l!�~0�\�@��fjϟ����v/V�9�2}�):)1KD��>���Y��W¤An8s����ǲ2��]v�DUonDQݒ%9hp7޵���蕎�Y���ILL=��E��kpe��!V��z�w��z:�cGU���t�A��̑m��Fmɡ�y���6������(Mtпr�Xo��2�u�,��WKL��N]��K���Z�X�%C�V��OQ��ÞF�:������ʺ�|�Qt-ʸ=r�OaBpͳ2�_e)ˍA�=S*�g1�����.{�����]�C<���QؓW��W��og���n�9�=~�NYJ�]��s�u�d�I�\�0�9�њ�j��r"��ID핢;�pw<m��t>�f��&N���æ�s�:p��i�̜"��F`�q"T���?N��T2�5
�5{�~la�]n�(:�~��Zr��i�!D�"�X�"t�_��hF�C�&�u,���t�i�<�F�O�X*{�����Wؓ}o���-�}4��,Q�uݥ�&�p��J[�^��Lt�
�J�H��B��k�#��B�k�8sX{I�O�U(	o/�Ϯ:N�����'=�/*���dr�̡�eO��Ai��Z5��R+O��V���ݵ�9�"b��L��W�d��M�>0���X����|���N�� �ͬ{�j��=�	�	]��-alhP|�D�㹣Y��������.�������}��,X�S�K�Z=�s���Y��D\��i͠��c;��>F��8ڎj3<3\w�_��};���	��[X�x�G��ڦ[\&N��-Q�X�輫���6˸%��%]jfZ�B���ul*PH�{�㼮���Gi����1%Y���u����ni���v�f�p��y7��t�X��!Y��N$��Tn�� �r�)5t�_��߮oŨ�wac�Jl�	��+�eI�^��n�^e�AF�Ԟ�3:��ϢRO��~���_מ�5�J+Ah7�&&'�Z�����L[��k����Pvɭ���gX#�_��ifǉ�;�L����*s�~�>�fF�3�x�`�؁T�:��x���+`�b*ר�Q��B��y�t���<��+aK��zP6�
Vڬ���uI���/���٬���y�����d�P{��D�"tvI��_�A�M�\�.�(�C��f?!�S�2�m��n�M
���T����K���e�*�\e.����8�>���{uܪ���R��o�1z��tV�k�ZY�����8a�K�U�(�J-��po����O@���1���z�����2��,ֆ\�g�A��Η��A�I��9ƛS���{ϗj��eg�v,�OcP�m�g� �)TU�^T]!�<,)��<T���2��vA��Zg=:��'ջ<�^��Ϥs�lnסQ=J^8g�|�=	u�!�������=�A���;��\^�| �˅Y������;m���]��tl��.�x[:�R\�8-_;�;Vv��Ӿ�eK׸hf��$�\� A�3i����knH{�p#��y�-{����S�4�=�zv>ӑ��&�Vo�Q�ػo���)G��8�ֶ:VýC�*�&�	6�3��k�*]�}]]Ov����,g�9�����.���zy�)���8���]�&�%B� �*l�n�xf!���0�X�&'��%�-a
��-\Q�[L���� Yo�ǔ�֯j������	�t=�S����	��CojX�d���&�9�50��G�(��=u������\�z��]�*"ǅvx�h�|�Q���~���VO����T�+�혧��r�"2�R�֭�	�p�;���FF��N�\�b�qm�מ��f�g����xy��꫑ʢ���*�R��@i#>y�ܚ�^�|�z������*�Oeĥ�^G��nq���@��g���j��;�ou�� ���A�;\�b�BA+f���ϞԔΪsy
V=�z��P�����%�N�D^����gJJ��cTP�f����uqh|{/��U�bF�c���3��4�����J�@�x;�zu�N�挧��^ڼ����1}�v`�v�
�����S �����	�%����}���^��s�bq,cm�����7�o��&�����3��'�XlVi-����e��)i�E�=*L@��K�0�R�a�B�fw=�{�elZ�Kᩭ:%��:����ߵs���wtw���.�h9�]�ϳ�k����~����Eͫ�`½�uU�d	��.ݾ�����Wz��s�أ=��J
a�kx��w���;���Q����כ��������|�B��T�����w5�]1��r)+=�#a��B�nFc����r��nC��^Q�@�o_<n ����;�U��ȷ�$Έ3W�Ρ�ӤY������v��E�q<".�%��1f��S�`��y��4��U����E���Tld>�|d�t�=�uׯ4d��x�_�=��iR>���M`"
�ҁ��C����B��n���H7m�(���~W�G�� �Bϼ��ZN�q���NIƞ���� ����He�l{��#f+��$5z}��3~W1�E>$�$3a�s�p#s,���ȭ�B�����~��3D���̉��w���`ٳZm��������@lCsog5�	ay�H��j���M��'����J;[�d�!�L�C�_5(��۸�<��B�LlSU�u����쩟B���$S}ۘb̍�-nفq�K�no9s��˘Q��͍9GZw)!̸�r�.��ws�]����fVǯ�+��ѻ;��)BT�ɉx�ݴ���;v��]4fP�<D��\���bi��K0γ���,�v`'W���4P�h_E��r��:G7��&f��;Ze��PT�)�5�%�mclW�~�a�-����Y��篰��
�	�T��ʞ�H���}�{CU9F^�
��(�`E�Aj�%���.P`@�v̙ݷ��G&�R2�ջ��W
�>aVwB��h�����BO�vY�ȉ�٩�5�z�я^ �Au����¹����F���ґklzxJ�&�v���tqԺ�..:�l]E�'t^�8~�>���	�SNų宍�΂�a�K���*���ݳ=t���&��K�q��c:��ȏ�I�Ѯw��sj[���Wa|�¥ʽ�}6tT�mW�|�b�O�����,�ԕ]νUQ"n���ܿkd@�R����hDwK�~b�O[�� �BrD���j�t�����ݤUxtʾ�,�9���?m��k��Z�9��rg��b'�3�󸛧��s^l��pa}�}��<��Yh��7�D["�+�ܕsrU=��b�}p{ޫT�GW`u�B���U�S`�5o��2-��6aЁJ�C�n�u��}Sr��QA8���Ք:��ik�(Ɗ��������ﶼ[YT�{2A�uf���	TN��Bgj U�`K!��ż���*^���M;�1Κ/�20o�fZ}�,Up��-��_E����d�Z����b��6�--F^G�:��[((����[h�`����٣w��o�	�'0����u���@�8�friY���i��j����T(R�g^Va�NFnd��[�sn�7�s�'2�;9�)��{���>'r6�TpBK�µ��`EN����ݴ�kPƨ���k�F7d� -F��.�:3��O3I8eB۶�a��]Y�'�}X�������&d��%*%���ڲ~�m���$D����Z =�(Jt�w���K[U�A���ł��6a��W��@����hu�w�J�vn�������o�� s��C����´��@�����a	��;N�ô�
�P��M�n���|iuF�)wn�WZ��XF7O>I-�BȊ!NU�hL�a:˥{$�x��¬�;�+iV(�J�r:���^q�v�nC\���[G9w4���ǵe^��X�9�H�;;h���`0�Zf]���/�ܽ=C���xv���r���ۊ�mMÕf!Y']�<�e�([N�'��W�u.V�N(��,zE�5�*P�׹�z�"Ƚt�,�:�j��t�J���6AU�f�A��g��rNO{���0]�\��f�67pC��7���F3�mK���S���י���F3NСswp��yH޸��0��� �i�q�����z��3��w�m<�9d6��(@�)�S���D�X��;,�Z��W)Dzomb۾�2�K����&�͗��R���z>��ӥ�bj�sr�������k�T(ސtF˸Z?6^G#K����Ul�z3uK�[*�ܜ��/�on]J�6�ڕÞ�wo]#�N��+^�b�=�ک��/�IX��D��� mK����egN���(�V���M�D�9X.q�כ���}�m+��bH�_L�Zn�J�iy;���f/����q�ه�j��[�rф����'���J�j�n*����k��;N��Ł.4^f��;��g �ۢ�8�h��1��km��\�I������m���C�p�f%����V�jÒ59��l��K���t�4k9T�k���&�D��I��cMm�k;i	��H	��K��b.k�+p��env�t�K�]�
=v��5j�%
<�D�"�pGQw���b�ҳ�:��H��v�̔Ug\�p��OY۱�1���Q�P�*�.��k^��Uz"�n��!��C2⎼ZԸ�U��#�:;���3f����k����kk�&(pP�B�3Ew�*��7���Bj;w�R�[nElE�)o�9�{�B���H�gu�*窭���O�ҥ��&
Yp+�6;f��W!�,�s��Zve�ٱ2�x2su�]��1�ݠ'F����.%��3��y���E��ݙHa�kf�W�嫥n�v�&��Zc��,nV멚(�fvu�'�ytc����3u~=�q)w�5���[_��	}����-�����Hp/h,jr���s�
7��rqD�ymb�f�ڛ�z�������&�2�E�J�h�e�vMեygp�Id���q�u��1u�1��鉔���E��'$��h��f4��f�wFe񊬭��t��G�B�(�h�O|�}��+�݊L�]��G���;y�7w�&���[g/�jZ����<��Wڧ��{��z��t��ۇ^B5�^�撑o|9yWb�jd �y�ac��]�V��i�����a���S��L'�agZ����@���(�q�%�{�[�1KW���ػ�wAk�(x����Y=+���z|�Y�%�[�"_@{О<m�vX��*���D;�޸��:0��H�+�{��Y��jQ��8�0`]��= �UG�35���ǽ^�=�0�⢁x�;7�o;AI��=M8v���7P�%T+���ވ�1��
�c-e��E�Y�C[6�a��g�M���Z�^]����v�X~�����S·8n��S��p1�h���w!QUj[7��^�$glrux�"O:j3X����{}G��?\���n�V�{B;��͋t2�y[G����� S�����E��m�'�0 ��5^Q9���iA�(�ˡٵ����&+qjTVF�lHH�n��5� �����9�-��Ynп��k�b�pV#�߸���';��D4��a���*�A�:'xjyA*���Ŧ�~UI���(j�0�(��-H!��Uv��P���c���77���J'�b[.���|;��1��.���c=�Ӱ(�b0j�J�t��9Tm\�p�Շ ��so[[B&H��BOQf۩�p$nh��k�Rz>��sn5A�
�wq�-:N����סt�ۀ�v�/:���x��`#Ն=8`fI���5���ƞ刨�T���za�2#)�@1A����U��Ճm�뼕;�̖�J�Y�~��|3��"����]}�kyY2E��(*}C���T���!|�(@U��~l��gם]�9�ʹ���FO�9\T�F� �f��C�@�1��
��e��wf��Ec[h�+�<�/��Ӯ}���!�	"s-�d�snUXv���{��M�W��:�ŧ�>��읮��3�<�1�8��9���i��Czu�y���o&�Z���0��xѭ�Y�Z�i���<4!�f+�&�r�)�?�E�ŲK޵I�nT����P|w�F�� wU_2�����@=A,̀�{+��4Q��'{iX�2�Z����9���jud7��>X��^+�/l�:��nb'⾡uwnV}�Oŵ�D�|�|4��}�]Se����x7,e���p�1L�����oL����C��B����a��9�Y6��m�)�͸5v��M��V/G�͈�x3��Lͺ��Y��c4hy��z(C��{@�1Y{��jw�o��?�f~G0��|�]6��q�V�3!�w�8}����l�j����#�c^�o�9���y���v�Jg{�����䘸@u�QKz�����Z���v"���z���/K����PL0S�U
��O�F�tV��Fty��>����.^b)ԋ�o<�T����~�����:T.�s��A�8D��zg�3{�I[��Do�|�2�~��/EQ��<��N3��1�2R�h�>�;;>�xeZ;]�r��<�2 MlQE�[se���Yo3z�:>r<�����"~��맘��2���ٽ��|���bX�{m���A��K6ZI�ԹV�}�����3i	�V8�ͱƐ.���'Cohwe�a"���(�	N&݊齖o�O	u�u�@B����a��OtȪ�
���F�K*�]��]9o���%vX�)��-�t�%L�#��r�I3�M�8Tᔚɵ���5���U�|}�}*��]�(��C��wæ�������1[�z�I�rWx�蠺�ڡ�9�����R�9�����'�UJ�aXQ1�M�⊹���{���c��}|K[T?d�o^�I��� 8��m�=�	��SF�e��]]߽� ȃ��-�v{���U�7�%��U��lK���:�l�n��	�C��.]+�O=窾���V:�ON���v�)���*���_c?/���(~���`�_.c�_N-W�QR��^�ry{�m�иn�յ��ϸ6��r���Jh�W��{ހ�^ǺTv5c���P�K����͚]f��u9�{==]O��c��x	���E���N)��u��sr�S�~;t��hoZH��}����f&���@�������U@��?X�V��?�����W�;�67n��'�_T&<"���x־A������n��ۅJ!�S:R��1�պ�9| ��w�B��78�nc̵�&�׳���-p�ډv�\hn�j��o&1n팇��b��EΛ�����ڤ.�K�5ڭ�[�y�����ٸ��o`�����R��Ӊ'uf>��{�s�f�]u5��雟k��z6�/k*�zʁ�����fy��Hu��c6<���z]��]X{�q��Ԟ ��X�k�vn�k�3�{�MB��������1.�H	o�h���o��^,�ZV�/Ԗ=������2�.��̑�cm�5�~��>�����g���Ti��f=��W]�ۖ���3!�y;-�Ҥe6
��i��y������gp���;��6��#�~��m�o�F�{�Z��[����f綑s0� ��ή�pV��R*�r���Js�{����Lc�e:�(�ڏͪ��U'�z�0f�3�P�y�w��A�=�����~F����(���N�ڌ��@_we���P�{���@�k�T��󯾱�/����a�Gzr�}!����w)��f��9�s�����9� {�3�｀���`��ꚿ)��A뢦����8��PU�˺�ܘ�﫞�3�g�ڌ�����\ľk������+Բqn�r-�������l[A���8�.Jԥ��+y���|͗dXCNcg��ׁ�/�T�QFD;��l��U3�R�n��WZ%+m�N���s_e�]HZд�����{3��X�Ov��rD��e��g��C9֡�˨@�Br��g�/��9��FgX����L�n��z|T3:����ۄ~Zb�Ω�/J�^v%��vT?yў��r}��>��߲^~�Υ�0�I�-���3ز=>��1s���IR��1�E?y�"w�b̞��8�vVD¨&�ȑ&NVC�P��Ո7�י�Ѓkû\MP�`�/��:A̪�7]A� W�u�,n>Y���������	f��M8�!�F�j�XP=4���<xǱ��Vr�>�>�v��~�.|6�Yv�(��Q������
77��[N�/DY���7�����9�q����:��X�`�m�6��_%8�d���o��=`����hsA3�����-������0�wn�R�q/�|{�SH��+�f���W$�ӌeܰW�
���F���n���>��7��{���揭�Z�ߚ�����	<�7V���x�.�L�m�����z-�ۇ)��T�o�8t���n��s	�Yl(8��������Y����V�3QK�(�VDƪB�]�GBqcD�5���In^A)�.3��y��Vsbsɺ��<jҸCСY~i��t���~��N)��8�K��q��}�ʰ�����x�=[��۴���HY!.0�SEwNn�mfWw�����F$�\uY�"��y����+9���E��F[��O���1��C3974hR4xs��3�7����o��M�i��2��u�J�Y��={��v����u��[��{�S���bG��e�WU�3�779e9�S�p���G�ت��J�05m��RM��ǣ���-my%0[śI�;Sup��=�V����(����ruC��tP�'�_�A���`o���h���99;��h������Z��fOc����5y���
,B��߫/h���S��6���\��Z��������?�ف��}Jynl�l��>du�gn�x_=U�6b�?7}
2C��nj�l�6�ƉnJ'���n��f���e�����\Vm]��Y\VW>Z߫����.heЀ�.b��e7"��w��"j��J���t%L�n��g��]KB�ul��?
�_ZI.*w#��hw쬲���Q�}1.���$l<H�󊷧k�'�Y4MT��Uy�wY.g2��H�EԘ�q�r}�����V27]^T�P9���L�����X���ޑ�GC������d�
�hD�n�^
����t�g���5�K�Y�/�>F:*|v�;�/~��DU5s�瓹��ǣ��������}R��ެ��G�}î`ؑ�vg�*�c�,�Fޣ�*���;a!�ݩ��\�ѺK���65�zo�3<��u�t�SY9B�&Hx�{0F;�gݝS����dW�| <�~�7�Ez�I�4��Fa����c)Y�
C�r=����}q�}ц�e��`*�/ۖi��$��Zzg¶�z�w�3�b�����i��έ�Sp�r�<ѝ�k�]�z�V��Q�q����;f<fz�\�\
�v4uw�؝�㹗1�ft�U���^p��dW[�#N�98�����nOO��׈��f���'�]=�۷�U�S#�n����?����K�SP�~p��
�_���X�E+і3��Hλ<�w�U���5�+o[��M�7/��{��Ŋe��|'Sc T�"��b�׸1�=�w����Y�B5$�k�j�0�"*,�CPE^���z��gs���ļL��,�D��p7[΁s��x��VA���^^+lW֢���&2�rx��Z:�n�l[u�^]'���"q��ᷫ3^�f�1��H�&wʢGÏ�߄ ��0��}u�������1��.���Ь�E�X4�=�y��LU��oʊ�H����.���[���1�wg������������18�BL粸L�U��ӷ;�8\-�y��8������BG`xi-q�2}<ܿ{��#��uF�e=���*���Dsb�_;�VC��Pk'`}�Q�T��ڦ�1�OLle���>s�7y�6'�}�3�'.6է��fwш Տ\r����}��߹�(���a��Ǻ;xP��ʻu�ډ��j^����J�����0�K��߫��A�SU�g#���չuF�5VO4'SAhx�������퇦^�>�m[q1�Z��Q�z�TfR8��ΩNZTn�&0@;8�q@�v�}��(9,Ou'x����Mz�/bY��v媐'[�hIk/1��n�0G�~O3�Ν1��i�#4�.Fm��V�fEV'SB aj�2��BӋ��lN[o�[�?t���Wm�P�A��JͰ��O�K
��2�W�?�����î��`q�Ю?歭�眷0.�:ѻNA4f�Ӽ� ̏i�jwk�ܿû���u�W2 ������{ݑs됋\��
����[��K���˩bG��2��uc�`�K��zt��x�9xz��e��<���c�J�L�3��싯<�Շa�
R]f�f��z�/��
u='�v�+a�0m�v$� ��8��r�Tע�ًcC��G����a��㍋�Ib�=�0��d��mD�Խ�M2z�� �*����4������q���W3y�V�d�#Z��8@��`��;��*�qC��:Y�oS^y��1�*�wE��^��k��Rٰw׈�Ȣ�q�4kB�TD���g�!p}ϔ�͋��X�H���]\�L<7褠�m{ �U~}���G,��i��#u�üz�h�iԨĹ�r���]����hf�:���ej�W!:�Ew��Wr�x+qS�㰪�nd}w-:��Еo&�X[�[kW��f��p�c�:IѲ�y,�j�/9�;����:^JƙǤ�VP*���Y��od+r���7���']��PA��z�e<�r�Z��C(%Nh=���7�ڮv@��Å�n@ci�JJ�^R��h����ܜf�п�R�zlw�{��S�tyf�G�"w�N�
�F͕��ցuX�,{�����K�ݻ��7�H�g`ր�hy���bSTxCN7����Pvh�n�)s���YJ
�'y�7*�'ح,N#�����y�Q.�B�e�fm�b���S����u�B����F�O�Hr��r���Í�7�b���J��2�����x�p&��4(lV�؛}�JL��J}Mu��f�ʻ%h�s�n�Ta��܋U��G!R�3G��
���hd0���es���n��|�����ub٬�b���+�<�����<UҌ^�.d�\1��˱�>n�A�&B^r&�Nк�H�Yc +Y�4�wi�����ٓ���n;�Q���]θ���V*�/�j�ܾ'E:�t(]�!]��rn�c���wv3���Q�;o�D�K)b�Ҕ�w�>��Y���rl*�ٰ�	n,ށǃoxF
Oe:;[㛟9��23��[w-1+N��=ղ�2a�����������k�	̓��;-��h�����3E_�]�n���\&>*��]d��F�VL4�������JiC�I7{����1M��2Ӭ��.�ٛ�u�Jc�܇n��*�_=������q'愠�K��d���o�{7���n��
F�����4B5{o�f��ދ�(���U�ㄔo]�Yv�!y��^*�L�=vr�i�c0��6��bu1�v��(�����+�|ͅΝ��\�BJQG�X�����c�5�of��JA���u��oE����M�FZ����3,��ɘf[�'0��!�`}F�,�4ų<˲�0tȨ{a_��2�4��4r l�m�Ui��H�$;�!��3���'E��rI�aJ�Kt]֎�'��������f*�;P,t���Lơ*�����]+7D�SRY�:�2�¶sz�o]ҫĉ��.�j�)}��:}��ޅ�X�i�솗ta�<��+�.v�P`�$���"�����d���ZWG6w놹I2�󱕳v�	f�`ŉ�pF]���V@݇e!%�OM����wFEc+���n�y��H��o{1<�S��e���g&YB!���{ʆ�:���IN1�1����u�=������0���R�79��L�0��+��=U\��3!y�Z�v���k`W�5'Ӌ|6X�:$z��a�Gn�M5$��W<:ۭ�ՙp�����Nu�}OYwaks��v�i�%YE�C;��Z�����l��s8�*�^�(�]���q-��^7�۫��}qڨl��8����;3N�<,��c�����df#Y��j�w|˩��0�����f$�M
&�d��M���興���� 7�0�l�O!R�ն�Ю����N?�
�i��f�ʼ�mFY�����׽���Qp�nI�]k5�;5ۜ� l�0l��T�T��B�@��[��+Ux4[Ɵ�����Ϩ{�����~��%������{vx�bcg���dG��IK��e�/{�5�����綴��Ԫ/��r;3Gtd�[�#/=;O�Yן>������b�xF���|C͒����V�ܨ7�4�����{a�'f��MvuȾ�+f�.�����ö3+�eb�;Q�ko�j��G;<Ϝ����~����~�s^Y�hdĲ�+�|WhsEDϏ�/(���!��pcMfFrtb�q����[{��kk�_�˥GqV��Z�w��.ǵ�/nagEo��	c�v���=W��h����w^���vj��L:�����~/�Y����s'��E��7E��d'����z�^Oh�E�x8{�d��6�Ҳ��ͫ����堘�"��5��Q����S��5������{	�3(��1]��h^f�d�rL7����2�4�ͭ��{�\/f�FH~�wsf%�dU-��-Ֆ����������:sJ�]ήoM��}�t��cw�V�D���F ��ORNl���Ȯ{�\yVPf˝]�ç�u
9����T<H�&��`�����NGU���륟��I�΢S��/su���g�t|��F2n���*�0zv�v{��&%�t��Ex�+=�B>��N����u��9o�:L�|h.}�l�^�NֿQ]A�����
��&ì�7r=ⷽ�V�q��2~>��{sz!CR澰8���ݽݜܺL^�KƳ�p��}�z4�B1�H���C������rd-{��~4�h�oT�ۊә����&��P�� ���T+�\���8�Qk-�X #me������>г��oװ�I_�`���G`oBY����c�ۄ��8��✜�*�Gp�}ku���~!�Y&����V�Π>F�t�����p��;ޮ��m�eK̷�nR̶�#ތ����Ok�9���ۚ��^]Q�>��9}2G��U#�O���ҭ�/Y�i����1�|��=[4YޤQ�w���\+����'R�{ŽL�r�C�����.N*�[�-���/0�4�;�҃�����w0TwY:�����u��O@��H@�c�N�力���.�h���Poc��o��l������wv�����V�y��7����#Y<`�Ǧ�8�^g�&s������R��3�`lӳ��s�OW�YS�D��I��@,n~'��E6�0fT���(����/d�Џ�lVU#3��d�.y��c��0�X�/'�,E���w_zn^L�F��	pPeZS�uh��,c���S�eE�w�Uj��Ug�a�z�r/�
;0�8qL5�T��%���0�4�-���=�9�0��7�����~p5U��7P�2]��Ϻ(���L�tl��7�ڇ`%Po�諺cM}��疟��_~&ն�w�N�K�o�WXC~ܗ�>�����Xz�}���:%⺍ؘ�7�
f��zA�����~(ߢ}�}ZY���l������P��Y��wp�*M�����'�(T{"�z$��5���Y�p�s�<�Z� ~1����z�f#ۂ����z=��Nə�����e�Z��O������W�8�:���և '��B����Qŧj覚�.��~����Y�N>�4&K`���;IV$�7m�����.�������A��KueΛ�Pŵ��a=sZuh��j��Q3m�ɰ��y�)iİ�I�38.E��v��o����%nV����zY���	��/E��<1��n��^o�x�s]�{��&Y�K�/Y��g�z��Gձ�^X���GD\X������~�G�t���W��Ǿج92*������W��tu�
L�{݋SG5���c#��y���/�>����z(衕�/:9�=�s��V��ؙ�Uu��p�?
u|�H>3}d}�{�~��&+��0gC��^{��x�h��p��\��hKy7�N3���Z>�^�u����|r��"ɳ���h:t˨y�dy��i�g���{kU�I����>��L��jW��oSko��N��z���t�{~>�,>� d�c�~�R����;��s⫔�<��Q�j�@-7��n��zc2j
|��B�i~�����<u��ي*�3g!F�����.*ݱS%�k�B��~IF�q�G��K�.������,*�+:��9��K��@mE,=��:��XsM�q��d;[]����LkWBKS�e��8L��j~u��z���Lꥅ���kt�:/cYL����y����޼��f��g[P�Ь��K�ր��[��jwl�Yr��c�US�/��;B�8�U������ތ�rr�ۨ�U-�)m������Z��� 6!>�Ov���a�)���e)���]�ŋ@z��X9���r�!��H��]j���lq5��}��g�Ж�0iaJ�סӆgz�����A��U5u���,}y��KV�<��Y�.t�O<��C��>�Hy#<����_���V� �,o7[Oj�)���yC�m�{a�B
��}����]F�p�I�=�� ��:o2s��Z�d�\?r��cyc�񙵥؇�z�T{z��XW�?VK�cFFa���p�Ձ	���nf�N��,,��R�~��V�ى�9���c/W� VZ�v���o��إ}�ϗ��\��}H:�sގx�-I�!Xgٹ9s��{!��v�;z�vϡ����u/�;�RW2h���S����w���
����'�m���s��� ���/6&4Z3�#R��
xފp��]C��ywݔì%�e<6X�,E�}ָP�}v6�R<��j�㖺NyqC0-=�h6�pG�7n�����Kq�-l�ƶ�"q�$�V���5CVq^v�}�Íb7ͺ�2�>�s��{s-f���}w�ٜ��B�IG�c����ލ��ϯ<��7ۿj����߭���T��5�1v2�UB�D�e��x�kg�n�LvŹ���t�Un��0E�A"����XJZ�n���x�wRL�b�Qκ������{Kz�fY�B�省Dхuh��J��6�����;�8�/n���R�1���n�'�c�4�՟�~>从��^���b��]+m��գ�Q���퟽&�,��l��,��i�lTN?ߋ��
p��z9[�Rm�j���zu����m<�ݐ�&,Nd��e⍌���n���׭?{|;�q�*_3}.�X!d�9����R�O���]}��=@����B�o���>��?+��D�yl�Ѵ�Oe����|!xs�kcU�j�ULz Q��-�8HUV��kd���7��y]���r�3�We�z���^��Q]B�}YBR�Þ��c��	����n�J���j�bb���.�9G]K�\��4���,��5�u���\O���o)�Y9G\)S+#��{-�̮����-!^����Ƃ���39����=�������6��h�&>�i�}���^���=;�o��cr�c���M]��S*��������^��k�"�S�����s��W�i�Z�&5Øb�{J���q)���ʞ����*��u��l֭Y,F
ֈ�=�f��q��8y��m]o��P�k��g^į~��2�f6��/1��ϝ��8�W�)�j.�#�lQ��)vn"�˟n,5���Z\�h�{7�k}���6���5L�Rb��w=*�p�F��}���Wla��:�Qs�b��Fo����Lm��q����|{C���q\������:�]���� #�l��[3�b�4}IC͜��EO�q�#���w�������k�Š���⮴���P:}JhIY;$����]P������1>(�հ���j�==������<�Ԥ��Xw4����c��Ñ�>LT��u��Jcu�oM��#wD[�yQ��`ˮ?��t�S�*T(�n���.�J�U�-ɱ�֜.�3�7��V�ǝש�=���Z��)��c�7��:��Ĵ���VM.T徑]Y�NPs���Ⱥ�Y�� ���Iˎg4`�ݿ����q�	��s6��'�[N����]*����X6�maa�S*Ǿ�l��_��~��2��~��;��}�mq��IyQ����h�Iï2+׮��!%�sn�AQ�Lh�UQ�s�jD��Ҷ'
��0}o%�H�cj��1����G��a����pKr<��7���v�Mb�Q�m!f�Ҝ���xns����"N�C\u]�:�W�\1�^���ʷR���F�sp�^{�x� B:z;��ҢǦ�{�霊+��׭��r+�z�5��x�~3��9VK��uǜ�� �S�W�p6}3�}����gp�/~NZ-J�D���i��^�Tw:�Y�W�*��e1����o��/��,J�JY?ZN�]�Ύ���߯����m�FM���.���W�]K��f:�ef[�ͺ����O~� ��N�H��F��C#2�f��2���oHN�P����;b'k�6�U�¦qե�`H�CH}ڸ����+�Y�X{;�V���}8��k��e��2���.��7�B<"H��i{��f�]��3ҟg31"��M���`�В�q���γ�\N[��s�=�WC����qS�q�q�,���:��lI��^�Ǐv�=��+�=6L9�����ں�oY�{��^�A�y� ����gx�x�[Ր+���D:��j�`g�GgH���.��As����K�>̫.�x}�ѹ�~̌��|;�4�j�
`��+Ȧ������4{���˓��>�_
*��</�qQ}�>�o�FE�Ψ�&׉�\U�����G�6N�s�>g��i�u</l�3����Te`"�@�{c����= f#-׷�Ӱ4
�gbH�sT�%J�Tmc��Q{��֖�{k7����Da�h�bɿ]Nx׋"���1��v�i�J�q|���*,���G|���J���=tVn�<讳�D�|���f�4	���#$�[��킏b��1xz��¼�O�z]��tP	�N{rj+�O�Xu
W��n�mU_��lk�9��S�b}��r���>I�N�`��+���хt�A��$A�r��������oy�4i�CCS���K˱t��r���(�c�+piޙP�S�M^�p�(�ݻ�G2a��*|#�j\k.p�ê�:��Ԏ���Kp�ҽ�cU��]�� �b�K!]��s/�m<;��wx��9��%�FV�㛰�I�kG��M}Ұ��7|1xL�`;>~��M�t��˿��Gj�)�F-�Z���ͮ��8�]D0���c	�WxPݦf�����h����ς��c��'�%9���˥sF����L��t(5�?T$�+�#��q1����e	�>~��V>�|�� �[fL-���3נ_T���*,uw�Ժ;�%_*������ڊͥp�U|� ��g@��O��z=�݇�9"�}:� �z�HW��ܕ�6�1^J���z绎-F���������÷�wv���d��PXY�cKs�^�'p�9���p�z�����	�
�Md�g�3<.��o�ݤr��&)GI��X��7��c�:+����Ψ��3�R�
�5���<W�34��>�$d���)���GQ)n{��3<���}��ٯ����.Ck*_�HS�����˪�9G7qj����y�}���^+�9�����{�@iZ�2n��P�-�r��@��᪥эp�`-2��V�!�/	�/E㶖��ͨ�o���_�v�.d��79lyv�,�������ߛڒ�{^e���V�dچ��]��ٗ7���|3��I!�yI!��{>>ݏ�"��f�)[����b�*��(��iD�TJk ����r�RBUߒE'�/��������?����[��_����/�ï�3�������������$�w}$���[�מu\2����ǳ�RHr���ձ���?.j՜����~~>?��2ݻ�X��ȟ�YIJ������C%�f� ��"��f�X���AA��oJF��{@MA��*P���]	*��$
��Nцm��@mK�O��̷3S���� �x�n,7+���t�(���d4[Q\p�3s����x
R�G,$]�Ʈ���;Mm��3F�i����u��ܚ�1�%��k&���eŖujV6�0�)G`J��
�KD�f�6X+PTko9z]�o.���%Zo%]lBVJ�)�C�I�CʽT��ǖH�&MJ�b�wk���i�fj�x���^U�]1~Ut.R�
A��κ��Za�y^�CIi�6t�D�nn=�1�!���p5���v�̸Ց�ESiB���ݬ�ѻ3g0�.f��7���ք�6���֖Ѳ]�����46����n��(��\�E�ʳ{Zl��q��b�{�uRc�����y1�H�h�"�ݥ��=r���$�U������B�6*�$��a�
m(�2�5j`d�$,+�(~�*a���2m�"��6p<,k�h�m�l=��n�B�i(&G�u��[�1K��/[˗�쬈Ѵ)Uۿ�_9UP�EL��SSO%iZ��	���"���l���Y�X��V���t�~�R�Y����L5��`��m��k/6P�F��Zʻ���b7,�s1 �m*�.C1P(;[aS�ї2���h�F�e��(Y~��E�i�fU�9 ���U6�ZdM��-ݷx��5+l�mGVl5F-$�۳HJ	����KЯJ�X���gUl�Z��w�0������&��J���o��K�խ�N`9�dh+�yf��f]�ǎ�sp��Zzn���L����U�i�J�
�֛Ӕ��*4�� i���V.Z��������#sk(�q�^G3o2�"�0 js&Jbg���a�A��Ԓ[�:�6��$�eӐ�r�4�Jw����i�oie��)5�V�%e��e]�ttۇhc͹�%d/sd&��wT!Q[%��������{��f���d��fB-���ꗂә�&q��^���/tǔ���9�VÄM�i\�d^^�D��Y��-Q.]�{��aC�0^�u���Q2�X3i��݇6���v୳k*�]�i��3%�f,����.'y[a�A�B\�P&V�]�9M����S�ہ�nX�d;�U��x$&CjJwt��Xح�g("�>�*�1�t�+�A˛TT���X?����V�"Si��VB�[v�n���r��ڼ�Î�.5�%ؚ�`:0�$��zf�2��m�u��2��z���	! �HI V1AU�T�
�*�H'}��*�
���
������T�R�U0����^�U�)$2�s�����m|<6۾w�	$�G���f�'wߏ�6�u��$�Gmp��u��7>$�C��e��YHk���m�$$���>1��
!ˆ���d�Na�$�]w.����y��IE��f�WOW��o��Hq��I[{5���^f���i�d����!BJ)���O^�m�5����p�I$3;n��{f޻�u$��y��[�^������)���/���U��0(�� H ��1�|>�6�Tl�l�ʒ�P ���
�Q
UR�5��@D�((��fR�D*���)*�@ *T�OlMi(�PI�PPEJH�R!ER�U"�4��TU )@Q($���*�HU*`0�4(�Ap          �V�p��J�#��   �@�=)։=2�J�5�RRP�ciV���A���@��-���ѡ�@�x���zx�p �
����4�[$v:�z4;����A^�o{xO-�H	֔�"�'��t( A��@g` � ���B�3�f��>��u���{�w_:o{^��O�ۣ�������mb��=���w��گ����nk8�y�{ǻӻo������������7>a˻�=yS��n��Ȫ)N�v����*�{�_v�W�}͆����ն>'��-O��z��gί��vl��;o��ϵ�m�.��`�vju����yg��o����V���]�>��Ww�}��^���3�����}��b����}ꪥ��#J�RP�I�����6���3�=}���_{t�{=��w�;��9���Ǉ����f�uV��s۷-]r��z��e��=��u��w[=ۤw���׭�=����>��mm��=����'HS�L�
*���l���1}�W��lm��oGS�_wT���=⒛w�����v5w�;��[�w]��Ǿ�Mzܭ�we��'�i{o6�n����X���z��m�
jPQ UQU��T�3.�r�:v��Ϡ�-��u}����z75�{\�kaw}���vW%o����ڻ���/e���5�y7gT�U��s:��}�F�a+� PO��E�m���ľ�����y#Kc�󽻫��MW�T]ʹ۶�|���ky��>���,n�o=����������2�:��n��4Wt�����U'�iJ��)�uvһk�:�����<���]e;^�^�}y���n��}�W���r�V�׸g-�X�s��kk--�f:�����yX�i�F��L�Hz�TU#%y�^��g�s{(5��5�>��mf�o���S����o;�ݧ>����<�l��w�w�__}�;���vOUt��ݭ�;l
�A��w���^����Q��1@"�$�f_]ӈ�;�{ܾ����n����vm����^}�ͦr����!�}��z���=+ޝ���w���|�X���xc�v����}��&͛V���7��{j��[�B
+�R` �? �EJ� @ "��I)U   S4��@ h �~%)TLd14OzD�UT�O�  &���%6Q䙨�F2~;�?�~?/�/��WfB�|3�-Wy��4\h��<���j��?S�|���!$���	BI�$��I�@���!BIb�$$��i!BI���!$��$$��/���G�������{:w��ګ�-	�֙1��"�����E�{-�&�hU����J� �;�"ۖ��Y�l��2�b�]hݫ�j��.KZo`M޺�����Ȳ�	:"���ƚv��Y״�f9S�"�%�W��*�efjdJ�7ndj�&�%��ܰ�B��3I��̿�P�&�Ҳd`ȠА�U��Xtn��!8���ޚ�L��{�Ǎ�Ő�C����5��J��Y�4�#�PV�a�4��v,MkU���:Zȡ$4�/�f�`�(�\�Ҿ\�������T�i�!$]Ja��Ma������4[�ݨ�7��G�t�.�F�]��*"���2��mQm�v*�n���(2�U��Tr��p�4^�B��-�y&9(k�3B+U�D;�Gq(��E����(,gE��R!V-�P�)�b=�Z�Փ쵖i<���pU��*�!��9)T)�0�j�SX�̦Wu���PN�zko��Z�P�k!$5�騲�2��R�+EZR�`Z�~�1��AP�(�яNt�MX]��Y��ԝ�<J��`,�k;z^g\/��켺�{r<���6'�)��c	�DR�ۢq1Xh9��f���r��f̛Y��4��Ѣ��� �&̕�n���l2�y��F��Aٔ���wB�c�tc��eƨ�I�kdv�m~��F��6\ǎޫ�ˤS��e2nn�s�)�O�j�l]Y�:�mXgekLJW���oHl=P��$Xԡ���ӂ�&ƽ�zY�^֫f�b�d����1�y�X��(LL����6x��nʫ�֊zʭtv"u!ޖ 5sq\KsPʫ{>�<���ݤ��F���p�̖�xw��V�l�c��4���T1�VC̘=��e��ϙI�ŷ�.e��hR75�J����˹l�UWF�X�udJ.Xt.�ׂ�M`V7)j��s2�K��yy�a�2�j���K)�n����Ƭ,ܢ�n�\��R�\G�m�(0]��-a���;��\yV����t%Y5Ǟ���m�����f�v��ԇ_1���!ěW�X�����AQ<`9VM�:������b3�b�ƈ����F"�`q�������L���֎g�n	�"5�VV@��`uiU�" 1b�h�*�4;pԆ,ʹ�f� Sn#F��@">~A1Y����û�#{�3c���wu�_|��!�hSn�駯���������X����P�H,!�W5�6�;���;�<6�����F�E,r�ݤ
�e�rÆ6Hڤ޺̶��I���?�ܱ��٬��v-�"�S�$�υ�g�uq��JLD���HX[N��޼8ͽ�bK�<�y���QE�)\�������|w��s���iN沼La֪�Hm�D���w���T�j��E���Zw,�)�o�V���� kM��l�+%gYbB�}�_24��a�e=�ɩ5k	4罿o��f�L�5˞�Cݪ��y�;��h��(��(�����`T���&"�!�Xb���N$6�Hpd�ć�'���� �1!�P��(������*M�a�i�䇜`m!�a�)9`s+��ɫ(`.�Hy!��B��ZX�I�I�I6��C�!��Y�"�@��������c<�� ��`��$�Hm�u2V���*B���!�
���1 �
C��������2HbC��8���d��7}~�{9n���yNk�w)�ǜ��,d��Rͳ�n;��Y��m�5�D/&���&=�4$ݖSWGi:�5�ɔ�hr��,�0�o3�̢.(�R����VdG^@I����J�+j,	٣�T�5�K5xm�E�ʅP�-�XX��E�1ݢ����2�9x�����j)&�FjAi���[�E���Y�E9f5wP<���P̬ءY��Kt�-$��MZS�+n��ʒl�W��<�j���/r�ܼ�PLVH�bƩ�*�%D�;�ER;�v�� ���� *ø�Uf��P_�C{DS}T��O,f���b;��u	�Z�+���K�^D&\��
��82^��^�`�ь���PK�&�G=�ɶ�L�;�C�Y�HfQ��d_BdM�KT��f�����&�a��S@�#w!t�,=�w����,��ظ�f�6�K-�d7I�+te4��Gܕ� Eq�1�yZ��{TA7��&T��jAlFA[�#8�BI�dܕ�T*3YZ���8t�[�H������W�M@<�T���������������ʅ�_i��X��,�]���*�JJ�e(�F�T8��"�4p��mȦ$�7u�#%�[Z`�_9vr6�OH�����{S+��鉨�JVh!u�����0��hHF�V�V���&��H�9��Ż�LZ�a�	� x��k��fäQЌW��()�	X��!���WF�
JB�&�U%�)��z�w;���wx-�x
X#X`cE�u]ݚ��'ZO�����#][��GP�e�Q�ٹ�'�0*����C����&�T���4�L��=;�[UD�F�e|�W.c�w u�e�4֣��Z#�pehJK6�K��u��)S��n�U�ͬ���m��5��[�F���DA�D ���tbB�r�YZ���)�0`��:b��)v�ɚF�Y����~��m��N)^�nK�W�6����^iY=��q?�K0l�	��0��CF����l����`��*�M�J�L�utS0[8������]�p3�����y�����N��/�gRñ�C��U���wt�ã��"付��sDv»yĂ-iESK
ӻ��P&�:n��a�ޛ$�E��1A���ʻ�p���6q��)h��]��y����2Ze�/,�6T�;�����o�Y��b�1B�j�[Q�wX�d(�ͫ�bk w4����n���M=	�q	�+�����-)YY��i�&��m�]�h�D�
S��7K2�5���4��Kn��ʎ˕�&uޝ�͗R�W�iS.�J�؞leSׁ�����4��'B�l�ܚ-XwJl�u���Y[	hX�\k�GMf0�QC�9j��m��Sifݍx�I�p{�`�ĔswO��ڸ�4�d���3��Jhg9������s=Oo�n��������Wc&�5#mm,�����U��jҋ)���C�]�x*�?=7.ɕ@�n� �Y�Beкo2�97vP �I/5���2[l�v	T�uU5
�'J��
̩{��P�V�wv+C��T�n�f|q^Zr��C��Rf4"��t�������Y�^�Ո�u�gM��ѧh��!"Ì7�3^����W�`bc�^EdY�����t�]`TZ�/V��|
9YR���%&�B�ՌCW?Rd���ʒ�J�ǤEO�h`�mY���-)�H�4P ������{[.k5=J"��Eݯ�̪�;��[��uB&�m}n���s41�cT%��� �V�8N%y��y��1�'M2�<2�(<�r�!*.�Dt��[��A�"�5Y�Iń���3���P�a�N)#$`j��6F�2QiU՘v5rC��]]����S1	�YTڳ7)U�r���X�D1�	���?F"�+�І��)0F�I;�.������Z����cM��J��5-��ېƍ&�aҀۣ6����Wr����,�A
AS,$�n��1y����"���2����%h.�U��A;A���mV���1�C�"y��L��O��7��]J9,�QDv�Y��� �lf� ֮7��g��l]�˳�yr��ڎ]'fM&a��/d�3,�o���ե�.ޚ
�c�G�&h��S7^��ڌ��7,#*�VZI�V����chV̂m#H�	6��.T���g0�˽%YŚ�����fn�9pIjô�]eĝ�C%FjSlXF�4HT5"46֤�3T΄�L��V �X�ڥyxQ�Z�/j\^���#�����-T������S����X[��j�c)\��!h�o�4�A�% Nё����9W)��Vs���f��)k,�e��˺�bM֧r��tQ7�H����wf%�U�����3"V%6a�L��T�RL @���&ԊQ"D������I�U�?eS�#�i:��S)��(�{��ѫ�%�*��.�	�%`�(�d˩T�,Yk�\��6yb�Bbj��#��Xً2T�Å&�i��S疚F�+cܱ��-#H�� 0�V�A�5~�{*9��l��h9��m["�v%�N��-f�܏mŋ����pԷ0��&��lZ���ެ��动S������7D0�fc'`���
ے��,�]�%��ҫgiKa�t��.��1����ؚ��)d9v�ݕ�i�;�c��V�J�8	"ɶ2Z�9Jl��̢v��~;��Q�m�F�Ĝ�5_Z�{�P�B*�(k�R�f��/okX �KGlޣ��ʽ��ұl��)]\6�E��f����n=�$�e���F�J{�"T���(Ԧ��&
�b�swNkw6:[��x��� ke1��,`:��t��H��2M��@6�suJt͉��Z�[_�%��0d9���nEQ��JZfAaX�w]X�GTǌ�&��T�v��9��,Hu'��b�e-(�<�8��w�4�$���a�����{����۝��\�m����bAd��.�M!�b��H�!�鹮�ӷ�X4��QKU�!k͔B%�#Ѷ�D�km��S@��n�h�%ǣURdƩ�Tm���a��:�I�H�]{9Ǘ��b�|2�䢊�ތ�Y2kNT����Xެ��h�2�!T��0
K��[gpM���@�@��{*fݥ�ƅ�'��ܳ���L�-��3	wV��%��ɶV�:��ڑ&���*�іAӆ��m�*�
�3Tv�T��5��Ȑ8�i���+�Xt���Œ��g�n��Z/Qj��f����ը�`^��T�F�C#Y��GD���f"�����iX1d��re�wU��Q��A�=��P�cP���N��v2r�7K�KXȡSgq=tкr���v��n��#ՃMn]�p;�A�vB���Ć/��n�,�aT��!�wsJ���VR�������A�4�e�/":���fԙe����6�p�.�L=��Je�O��rFq����Ï����
�9N�YC@��wM��N��ш�J�n��yXBRTvh�O�B��	O?D�5r��Ld2�ұ�&Ԓ�X���QPTY��P���@�O	tC���[��Qfn�xࡩ�f0UR)����Z��T�e��P�%�ճKת��+e-g+p\9j�nM�b�{-� 
�V�鲖���C*ر��IO�ͥ5f�Ӗ�e�����,��k�3U@%�+��_�X�T�2l��� 5��B��r�S��R��3�XZ��@���p��t�Sv�SyS)^����t���0@df_��to�*"u��dqm�ȁ����Kt�3���lE�� kV�� �ե���V���.n�N�E
�
�#
��0˼̔���BM���6�e�r����71�����Z��	t��-�V�zBZ{ytYB8�nL����`f^ٔ*1nbǎ�n����ba�����Y#5e�L���^iE�(K{���]*X�P�(O��--]��Y���n��#q��0��W���nf�1E�i�Ք�D�-p2�GG	��n�zR*L�B݉aBQ�*�N�]�l��f��|�I�fC���F��Y�IҘv�1F&b���J�\	�G"�&R�ؔjTv����[���qɲhq���8p��!�F��2eMa���BU�%��	����!r�	Z�R�r��ǵY�S�)VP��S�R���r�B[h��V]���#U��E��<z�2�;��dhkoSD��Mi����twn��a2�E��Vdw�M���eFXM�y�ㄼ�-`z�#�ͼ�ݬ�n�c�-ju=�(�Wm�M�0Z��`�L�v�YJ���Z�����Bʽ/ZD�y����&+����L���O�� ����5+ao#D(8�&�Y�R�B��f�²��LU�&#�O��2Q��X4ե��piF� �O �[��ƽ�T�V@ԉ�QI�d*[�)i5�d2���)���]�8A�kq=4������6pV�͡R�a�Eh�d��QU��wLm�5�F�:��l�]�-n�n�֪,8��V��x��ux�栲�D���`�>�{Ѿ�G�H�I�#}$o����7�F�H�I�$}$�����7�H�I�#}$o����>�F�H�I�#}$�����7�F�H�I#�$o������G�H�I�H�I��$��J�Q��[���Y���&Ÿ��b��
���4��)������DZ�7pϳ�2�a��횷�����$D��݄��;	���X��mBpۀ>�ξ���@e1f�*��(��f�b�TVyI�sOgE}�����h�U���:v	�\xћ��eA�"�厝���.��*u��;ӲZ��sZC7�h���6�Z{��v�5��FK�cq��;U)��.��η2�PL�ۇ��k%��d�w",Е}�{rT�'D�x�Oٱ���vqi�盛���̸�L�ܻv�;�>�f%p���
���:`�ޣ� ;M��e�, 0�,ݡ!Ȇ�����7]FF0V���B�~�]�L�����B���g�
䨣ζ-]ۊ#�%|�P��5N��d��v�U���9R,���.��_m[*��o�����M��N� �#��a����|��}�'�_]ei24	��ޜ��Ovn�WQaG�)1�!�='��<QT�r��'��$�s��um�)[aN�N0�"���-�3�-��-��ee�^k,f��J��u��;�1܎��:#7^�Ŭ��jJ0r��'����r��8��v]�j�á��,�(�(j���N�9�d,�I��r�����z�F�6�h�����Wͬ��C��ʬ��(�E�[Qm�����`��j��n�����y���[��ti���v�O�A&XV�W�[�ꑾt����������׳2�����:S�\CL���W��|�$��	���Y�����#R����ʹ͋�����c����C]|����ڇ�`���(]���	�!�l��9{ֻ��
��n�7�QZ9�!�d�kkF�O.��a��glk�ßo@r�͙����w�8���~����d��P�4V囲��8Ff����nNv�.��O	ë����]{;�ׄᱶ�դo=��G}]�>*��R�ם�v��V��Y���I����y�+���Q9:����q�s�R��v`Y�������}����d�uv{o�u�!��2�4�n��RORX'&u���k5�NN��S���*��-,�0h2[�܇$�:�/����?]�:v����2q�D�F�ŝ��;βv���!�Q��:#|��rc�X��6�Ð�le^<Ĕɡ���24y[�y�=���{�R�73��"�_H]�r]�>׌�T{�����1K�&a��v����}҇C\1�����0wdt+���k/��[y�Ǎ��L:�N��/�vd��Gq��-��3�8V'Y�zd&7,�b��Y��K����c�ڬV4��;F��s�N������+G���Q���s�C&���*�?!�C:�Qk���� �HĬD�s޻�t�d4�gs��.U�np�"+��fܽ��x�u#�PM�/5�%��^Z79RO�d�Y�i�X{wl̬"�Y�<n1N���3�����h����,��{�+%Y���^���)&���Z��Ã`�#�v��b"����$[�+ag����Ʀj*�)awۘ�4�ݲ�l3����`/2�i{����i��,�0^�z�X�2��4��'w7��k5�յ��L�����8��������e#n��0,�X��cw[�q��s}�:ޙ�V�4i�SC����O�N��y�>���p�QÃ�tv�R�D���Y��:3$�s��ڎ]N9K��+�2�Z����]K��|�1h}��#(�f����\��JM�6�.��B{���}wE��0Ey����e�@�;�9���(ǫuu��蝽ٕ��F}Jí7q��:�:6�_���s��mn��*��W�����Y_C��k�xҨ���Iysuv�]�3aۼ�I]�b�n�� Vu,tJ��K6qȞ��ŷR���<̕zbF���\�E�]��fV�WH�ǉM!��u=����ő�!Q�b��:���YV�����8ˎ��E:��e�˶�����:c1���V����owg+��6�I�"*�����K�<�ڡp��su���U�Zm�f�C03e*븱h T�SH�S[�����_�{S�[b�jJ�S��4:|]�}�7�$)ve�D�0Iy���1b��ֺ	u_X
��8�q�Sq�vr�v��gq��]r�q�[+��n�!��3�cC��Q�)q���1E�����ǻ���#hg\�I�ކ��E�U�y��x�{O:����=��	]�W�t�Y�o�Y�ݦ�����]���%�O�����BqSȷ��v��DP�#����=.˦��nv!�˹`���SUu[}�������+�r�d��}{�b�[�Q2ru6��hZ���Ef<��ٳEfT���L8�u��-�x{Y���QW30^�٦����'K1W,�joj��_x��t�b�%q<n�2�&_۸4�z�p��qU����&}�v4�Ecv�r:�$t�;�a;�l7���+f�� �R�Ł��jQ���]�X�i|l�s4<��rܷ 짘�XY��PUd�B����Ւ�掻swu���׵s%�T�gYAީҁ�e��
�\�3{�4*ܖ�SI���V.��e'֢1ZwW[�(쓉�Pòl�E��g����]��+	� W�v�#{�/��w���ui�yn�n{��l�T�MC!*e��d�h���Ex	�����K�8��y�A�f�H1�r�⫔�*�x��C�'&�QҰ��f�ڰ�\�9A����L��$��3u�N����Z�SJ��e�RUlf�II�,�f&�<���t�����ʦ9��f��c͗�p+��Y��7p�7V�\U�唫�����m#�έ��f�NE{*����:���9֝Z��p�wv�X5��Z�f7�����A�� ��Q�V�'�i�2hKl�t��I;�2�!���N�m�왷�a1���Ҭ���Ѭ��u����'h��Sy�Mt���K��)tWS��'Lss���'u�D��UgE[=DY��ݲư�;`�Q��bi�ts���b�)� yd�dyX>��w��y�E�_*�M���V5r*�Z��uy���r���[�U�J���0�t�#Sy���/B:A�ne����"t�ɪ��\�V�µ�A�Y���
�0v�z*�<Yv��{�ȡH����<��w��f'YgrE�z8K�S6o\�64T�W@\�]΂��xE���[�z��s�\����#mR3=�W��l�vdٲ�d$+2t3&��A��(9���z����t���6��I���c����S��6.,];:-tˇrB���ɚ��p��,9͛{u�[;i��7SE���&ʃ�\4�u�l��#��ib��s[�n�F0��HG]����`�Fʻ��_�ui�h[����!���WF�M�Ûb&r�s�=��~G��2��eΩ�%�ݲ��<8;?�#ky�eȡ�6ȼ�-�1�Mu�˼s�
�tנw:�d�����=.�pa���d0�;4X$�@���郏+��[�Y5��%�4��e��M]�ޡՙ�1q�h1m"�>�$5���W5,9��vz�w�|���:eJ(������x�Y�2�}S3)�Z{��F��}��MΧ�@@b��s��{Kw���x_%���t��������mh콮d�D�4z��������^�K��X+�H*�cN����t��c��IV�l�7%-��p�|=fY�Ge�2~DSs	�����B]���k~�������C���<.�;W��X�0�B_nͩ���͡���⫭�VPe
�O%!�ݐj���Ә��Ί0j�v/r����:�P��[%��ɺK��1�q2ٚ��[���;��v�G9wQ��bV���%:ܝ�3fYb���9p;��;��w���;�<��N���@��w�iE�Y��mЃ�FTZL��f���=�U�N���^kvɈ��ю�z)�Se�F�^q�͵�xl�0;&���x(C:r"�q�#�I�����B�=Y�z.�<���͉5���}T��T���t�Te�բ�ъ!��"�%�U>�ھ�A6�{����u:mИ�v�����{��ʲ�b��DM�v�Ƚ�u������bb6�s�����FZ'wV�ո�L��l�.���u�����좥ˍd��{���v@D���U�g��P��rz�Q]�b<�<�����P�%�x�����C�������x&���b����L�qs�\7j˺u��cm_g�ܕ��;{cG�ƞ��j�;()�.��-W5R�I�I��X��G���n�B�����.S�����I6��vo��1���3i�dc.+;��T:H�t�u���lv&(�8��2�{�歛]���Q�)�E,����/��ST�������5+�639�2f�����v;6�c�M�k'��o^�ٝ��IM�u�mr�8��+�����
�AF�wү�9 (��b����05�ld�}6f��A8�M�1J�/��u����Ȇ��9w]��Sm�A��ͣ��V��$cs�Of��uz��zI���۱�oZQG.��pc��2�wC��T)f���g�Q�*܂�z��ڱ�YSc뻂�]��vX�8�Z�_Վ�L�V���o]���뒥8s\���n=Q�r��^%ғ�Y��^�N��g�kCnX{q����͚���۳y�+0�k���P�	i�'����@;� ИK">=�+�[v�b�Ff�2�P�O��:R۠Z�oa��6[qH���U��h0�]ɗ{hl��\�!3e53vZ����v������ݎ�z:dx�"�¬n�B�}�>ɽn��,uV3 �0"��ȫ�ۛ�/����0B�����2���;��3���ҖI�Z����	�x��+][]����԰��qL�3P/�F'K�e܂�4��5M���c�g���.*��W<���U�|��{/5�F��MD0V[�i��}G-įvfJ��9�aM����A��G�:+�;�0�hk5n�s
=)M����x���),·Wj닯E���\�v�29B��*c��Ydg#���.�`7q ��y�ԛ����з���/wVr�;��'J�vA�Oʍ*�(K#u�tH������V�s�t@�滷�-p=- �ѓ"Y�a����W�f��@�MgqG��>�Sf]�`[AG�Ök`̓�qb]d^w�|2ȫ���\ȭa�������<%�U=�U�dńM�zȹ�����u�B]��6��Vo,Ʉ�@]ѹ{��'`��S�ѣ���1�=��ܡ��l⪉�"ޚi�%-}�$�U��U_�v3���@o'M�mh(�Wk�np�pL�`m�k���j�ίgwsW�R�{�#1�K��o2`���:�f[];2$������-��)m�U��HJ÷RMȆIq*@�N�O�N�I�q$���Ur�=(��z9[�7feڝ�b2�g��ͣ�l�2�CL�ü����3�o�goͧ�(�Oi�i�A�����5Y�y��s�Xެ���sw��;vM�M.M�>�H|�4�o;�˱�R]F=7�Y ڼ��Ԍ���);yR�Κp��p��.�:N�`�34ZS�ѧ����_����e�{-��5Ò�w}(n��<�Y8��|�����4��jo2-���qj�_��3�`"*�L�r��f`�+�7���r���5���E�О��5:L��=t�BC(g�|�ջl]�:ﹹF�g`��
T��!F�S�9G_gm#�m�{r�|��[0N7}�{4�S���39(�o*3���H��7��)�V��f��]���<Rt_>�v_��c���J8��0;#~�����塱q�#��u!�&�u2���Vmm�rk�����&�h4�y��Z�ζ��u]�-�ɪ�a^���w.*�ٙ���!�r��tj�I����s5�1�xn;8�f�����_r���s�w����&̍p�o`�<�C1fҖ_#]xQ]��iy�,��Q�C52i٣aA9����9E�r�M_���?�AQ�D%��M�ahW��J�F�Qv�5�Q���W��*�eZc�\�Nu�5˰1��pe�%��Ộ�]���ꈕ*q��o��[��_\�<:����tܻ��q�6��Z�^s���B�wTnVlK�-��o��緈�4�F��%S*��L�ŀ�� F����CMFm�i�<w�A�����κ�;��%�RƯ���u�\1݄v�-�N�oJ�j��&6�RA^�[��`m�0j*�4�%jf��v�ҧ�]9�s����i�{���B�� �]'��7�����X�R*f{̈́�>姀���/4����+�dr�=��fzz��it���WZ��Ұ� <kZ:x������f�Jԣ�����]��y�7#JP�t'�֟)
����A�����o�i*G�:n{���/.s�Sx1�`"����J�
�I�-�)b�)TX2H��6@k[��sH>�a=4���3 �0�0��[��˽�qw)�[yy/u�[m���8`��u���,�}�Wm����ȯQ	m�;�uE���1�*��LDe��ۏ1�����cXy�PHM�U�c\BU�V�fL����ց4��'J��
WӪ:�Uכ���V5���O>t*���{��x�g;M���wY��$�����x����!m�{���j�B��酦i�
2[�i!>�31��G!��:�L�(�h�Ou,k�ǻwdc��g,+�.��ـ��1t^��d�x���Kp@w
�ϣ�{@��^i��F��Da��J��z��m��lY�C/��=t��Ougf:�/�r%Y�K��n�V�o%����[�\ݺ�b��B�,�L-Π-����)Ʒ��}fҽI*b�F���9}�����<8s�7�{�����		'�I!B�@�?ܐ� � O�C�H!$��0����$1���$��d��H�	$��$6�HM��I� LI'I�B`Hi�Ԅ
�:�� ��, V@��)?�$� N!yd��`IP���:�q�P�v�� VM&!gM0�@�L'Hb�
�7�́� (M�6�Hm
���&�Hy��~�OCI�	���q'u y1/�VBVH1 E1�$�b�%`C���$�Ԁu!�Rz�
�0	� �c<�tͰ'P�,�L�	4�|�0ש1�I2 q<�"�0HVB� aX�XV8��,8ͱ@#�b&3�m�~aԊ.R��CV`i�C��$�o2I�7d�|�I� d�u���|��BiR<��m� ��Y$�Hu���R:��(���$������0XIj�;qXB�졾󺄁Xv�8����2 X����I�BC�0'=a y'+�R��!��ֳRI'+d$'��&��7mI y�� y1����9BIǬ:ϙ /i��IԄ$%m�&+�XB%`@��fw�i$��|�N3N1BC}�� ��l �a ̄�t�	��v�J���قI&Z>��ϻ���<�u�H:��8�I�	3V�5+7�'��lTd�q�M��9a&�̄zϒ	�C�D��&3��}{hk��Ӥ�q��D���ݼg�2����{x`�x���� c8�w� yz�>@�t&o� ��)	�ā�� ����C�Oz��\�k�b@G���Gz�>ےL��
�� fZ�4�&a����wz$�d4� hݽMa&e�Ԙ��C=����Ir�e�_}���R�|��La7���RO�� ^�{�	;��0e����$ګ q�^!7�������[��8��3;a*�,��(K��@�{��C��=�rH�\!�2�M{{~�/ל�}j�`:�h���܅~=`]�ۨP��%M}��?7v0h){l c��׸C��:�$�9�0��j���\����@oֺ`f{��l�ak�͑�t����K#ə�5�7Ǻ��.P>Tr��>2��o�l�9��t�8�]w4N^>�=�>K7�6��[�4XT�%�۲s��Pj�r�Zր�ֲ�P̐D8{��v�D򇟐=�������7��s��7�3Pz�s��{ZɃ�fo25_Y�ZS �.�:�ѣ}�!����2�����5�\�{48:��'/3Z'4o&�&�����3�I��ɡ��7v�̓Ow�����I�;2C^u�����d���:\�Rhﰇ�C���̓���I����w!�4�2� ���70�/٦L7����o��>���:!��m�k0�=������h}d���c�}��P��$>�5���#�ӭ[�8��ڇNo	.%��%!P�-��}}��_R]�Έ:��Rx�m��)�Ly�C;@�\�p;�wP=����_t�Xkﰞ�!���܆�q�;��k=�f6]�S�̐�X;��|���Ӿn��y�s���d}�������&n�[C{рk�w�h�S$1��쓻׹����fY=���9��M4He�<�g\[!���z�z �;�G��~���'3\����ֹI���sv���P;���@.����=�@{`]��L�=�}�d7۞�'ud���v�����@�t;�3)ֹu ��l��O�f�P5�d4�~�q���a�ɛ����w���k�d3�=�<��5���5߭i���s��E�m�)��X���7c��)|�v�n�Es�R�3Ka��Y�YI;&W]��W��p��[�Xí��6���xm���4k ���k�S6��H�>׬��;K�	j���h�4봵]������E��^Ѐ�H+)��^}�D���R�D΋���i��9��+�3�����J�X�#��Hi�Ȗ��uw���������3:��� HI?����>�  -��������ꪲ�B��6����)���}o&��f�o+��5�l�f�L�:`�uoh�,q�,s��8V�j���M��|����5[��O\��*�� ��CF��' Z�"4�AG���G[���ޕ��]�bFzmNV�s�3��Iv��U�V�އi�-�I��2��7#��/�E��	D;���#o�m�v(��ޭu�)�z�["֚��H<�[3���o:��=���N��=D��ÅOٹ���ge�V��́�2M�t���usG���� �u"�6�WY,?Ӌy���51Iv��7VEܩ�;77f^_l��m�;��te��I�32���L��Q�U�'��)�x��`-�ʝd��_V����lP;��sF)Z���̵��ix�K˨3��H�͠�'F����V>X��u��t��5zKf
y�7�ooK|�Yx�R}>]�by�H��1��ٮ�V9~5,6�Ic\�����ݨXف�0{��;q�؉b��)�g��e'�R���0���6hW&�邲���[��.��ڰr�u��VoE���҄ɶ�@�\ Ļ��;zw>"]D5m�v��.��)d\]%R8
f�;c]�4�@U�YԞ{p9��Z�����;�\����ii|�7�>uՌ�ѽ\MQ�a�(�nt}:"�'�ߡ�ƌ�U6�#�,z��g������=�q��)��鿯o��xz��L��ˤ�lٸc.0CK=�b�ݷ�kDvCϩ�;�������,�T"}ߏbJ�-f�Z���Rܾ��hwf���3�xJ��C��]�dW?�B�!"���	�	�����1�H�:�I mi�d��:��1�}d�XLd �$�� m�2B��v�4�(H��Cu	��=gXHB ����~߽���^���QDAwj;B�Db+ �WEdTb"�����"e���AT`�1EB�|�*�&5O�֍,DP�"J�`�"�AC�1U��ق0Q��DQVE��E��¬��9�Q��*�ф1�b��j�7���p⊏m"��bqq���P-� ����,DUM4D`�DQO0Ğ`{�1I�EUPb',��b"Ȉ�X��?~��P�D�8��`�0�b�����F�" hIQA"��V#ր�R�ߪk}�����=/���~8��R(u��*~�1�U���g���.Z����HcQ��CV���VEA��k%V,��2cQe�Yb��݇�`�AG,eQTE�§����QR����i��*���LE6�ʢ�1{lY�UU�s��f�bȪ�[�"��M����4 �����L���1ݗT?8�`��H	 ��go���=Ì7�X��j1���0Q�̆g�]TQ`�}J�IX,�DEUt�����5lQQB�FEY��&�\j�EQQU[aD��g�/�V)2�L�*"����B��Y0թ�����&��Ȫ1\g�����c�DF�Xm5��L�`Q�1S)���лj�j|�A:B	��׉�"-��A?AF���Tee��G��t�A��w�E��ԕ�_�V��1]Z��g�N:�DE�|ԕ�h��TE����m��h����b���#m�l�UQ���(�,b"�����z���:J�"H(�A������c��͚��J��m�f�[,���*�o��]w	��®Y)�s���0D�qEEr�n|�Ty~ͦ!��TTY�Tg���C)]��
G��#�h�]Z(�qȂ����j,UU�rfnY�ER���jj�玵YԦ0�Xor�YQ��ʫ������2D�?�Ҝ\�r�3IQ�UX��[�G)U����KUY�N\�XQQm�#�0¹�}ef��CQ�����m�V4*����R����w��Sv��X���׃����AK�
#
��\��u�4�+�K�wn�طV��=�2hA��*�ݦ��*�j�)~u�������@�A%���d�� �I�o�h�Ɣ��o���ʹ�*���[Ps^���[QR�cA�pӤ�A$�� �>^�or��a�����PDq���U�
��fJ�}��$�I!����ci<u$�(�ʟe��luV�0(<���Sb�Z��z�Ҩƥ��:�,�V*��U���{v(����0A%��5�=ˠ�=���]� Ě@J��lx�#@�E6} �2N�e�9��j�B�s��u��f*b��n����^~��I�����o��B�Q�M5w�b����t�~���d2�$�j�xNI;4˽*��:�2�
���!%��9� �`�Z�m��|I��Ǻ��/�^Q*���Y��d���W^��v{�����S�Q�k��Q��007gY����ΣU��5���қaF*n���^�ef^g#�7z��	�"���G�ͻ�z���3�kB#�0���ːPƥ�Z֭�\��3���T}lb���\7���A�7D3k� �P�#�D���(y�d�{�٧f��� ���}��}y�j��O�I � "���;�&�2i�]���aj��f<a0�`�����筞6�!/HB&<�${��"���,[�B��HH��Ԙ�LG���uJ)�r8{P�W����������p��Em�"���X����y� S_&a���� ���p�o�t���PX��Y!?���y� M|H�D#�*���x,(��]\~9�N?k���8s�����/�)i!�&�4SŦM%^���m+K�h5�b!{jP��Y������C����w�}���B�S�5�9n?������B�`fJ羡����=��'U/�ؿ��(���^����w��A��7��ځ��La_Qn��u(�m-�.Mek|n�n_�ɗ��"�ڨ���i�r|�����E��ݎ����o��&X�%�!���вJ�A)\J F���P=A�I ��(���y�h���(�P�A?0qǮ�t�)��8�sZ�OK�拶9��|>�9 ���U�̔�v=�H�!��L�}y�EGP�7 �	i﹭ɲ�}���6�9n�Lc���S;O��6��ˍ��a��Q��5#��k��+���o��sk<5��}�a������1����ݡ�k)����Ͷ���Zח���n�į�~�)��(��Xtmyߐ���sW͡v�% R�RƘ?�O?M�Yy,����y��oJ�p�9J=��=��ģ��[XX(��IHE�����5���7�"��C� ���ڰn�!A�}���d�H$#�.�Q�=���1�ݩ �<J\~~��_2�;Y��-���q����.Ĵˊ1c��wX��J���ڵ9i�U�6�:�k/S0��平a����k��S���=���fťCo�**�u��ϝ��7��յދ5�Hj�3&���	4�#����������i��޷���u-�ڐǛ�K�H���gY��x�k5��:�8��h�f
څ�z&oX�wi{#�	&�J�uuq����.�[~�1�O�eL=R���,��T^�QJ�2өGMK�}w��<�^^DG�e�%��B���\� ���*}I�Dev�����~O��=�rش/��3������A�%a4���6�}��#
���i2�Q*�Mg�I��qGٮ��<(��㊷�=��X�xW%Kp]��>@C���%����E���T��R��.M���5�rf�ֽײ���Ƶe	�BrNU�ㅈ��˧<n�{�}Ï�7�ͼ��"6K��%�|��a���q#�TZ���z�$`H�-L�ba�`��,� ͟�w���Y�xR>]����@�p�4y7D$f(	����o�|�x����ƤAEx����{�qb�l�`4o ����y�� ��.��~������9G/6@�$�Dz;�����+*9l&�f�l��5����>_Y˜~��]�����e���l��Uh?
��Q_�Yеu[��PY�Cnp��řEq��(Sd?/���M"�;�QÈ��!aP�o�j�/����	)(
��)��E>�P}�7Z9�����c������ˮe�����l;��oP�)�a?#
?a2�t�Ć�VL�"˧t��	�M��0� +iJf��������:�jW�hy����C�Li##P"�H3:���a���l�0��^籱ީO.s���Y �2}!
v9��wx]�`����D�93�
�a>�e���s�b��1h���L��A��2nXC�t���`�vKr����=}�n|�' �־�;����{Gu~��򦮭��#=}�Q��ڞ>��b��6���qk�ZkAΗ�
(�$�N�n��V�����ԳG'g
�S*E�ʨ�V�Cr{��NL}~i&��Z�@�����y�n�ff����ny�l�h^�]V?2� DJH�_4~��T����N���J�X!((ȥ��&K({��H�D>��*��(���w��Kz�j��DD庵>�ZoSt��o���@{ ��}AA�Q�[��e��1�����$�E�Eou�����0FCeo��u뗎��(�PL�O����!�d��>qPk��y۽�\kg5�m��ڻ�ǭ�D�"�?��DQ&���S��t�6���s�2������a���ɜ�n/��C�ھ�ޱ��=9��4�j��E�v�_|qPby�5GqlB�]��B�7� ��b�!uWu�-�I��"�����[w�c��c
+��U�`��'5W@�<��>_@\H��zt�$W �k��?3�6mԌ]��d.5P�ɳ�|�)���}���moP~��J�8e��:��?"�!��䁥�he![w�D��r$O��I���m���e��a
|�fA8�.�����|���,��iH�Q7�EӨU|���$�l�Y�;@ݕ��x�����n1�6.C&�Ĥ|�7
����F�D<x�B(�u��h��Nz�$��I��s˽C�6}�W:o����9�n�
��7�{�ﵼ{�m��~iK��j��̴w��L����=�����M���i�ox����:�7�87<s��:R��_�]
���;���鿷~m���7���}ɼui�^
��yM�v�`��N����Z�s�vq��pwR�=]��N��K���).�d̳�r����Ue�o!�_�z���S��ݼ�PD�zn�@�yT�#ȴAvѣ	,��r����� -'���#\���B�c^�g��V���̖�%�w�B�H�K97�����!�������V|rUc�Фp�����m��>p��D�A���Էӯq�� _� _��a�	]#.�Ĺ�ɒ�y������8B~������@�	���,�{:O���Z��Q�'Z�o�$L��/E[j�߇��1��]�p�7B��@ ���P�#����H��D
N��h�H�"!D��~�l��1�/aw��Zɫca�]5:�h�� �=���ﵘg�k�R!O��H�e�y��ovx,����L O�yd|z� �Q�i�ԼBLɥ�_3I���%�CZC�'D����*�7sLw1S[t�I;�m�'�ٰo�T�e�Nb���QYU\�L&Qx�|��S��|oo)CǱ�*��7�d��Osk����S�+�D]4ƈ�<��`7>�k���?1�	a�Ti</�xDH��P4G��(?}��f9�m{3h���a��IIЃ�5C,�
C��ӻ�R���.!�%�}Ɉx�$&b1z�_Y�AP,)����F���>0�k#�+�i}��2��'��hw�f	6@�>m�s˭��������_L����}
�a��&qF��:P�!o{��:?�����@�'�d:}BN�x�G~�L��0�-���E�)� H�\̑J�����m��AQ!{��� C.��p���=0^s6V��C� #��Gi5��=DwgUݪ�;j�����T���C�Z7g.Hr�8Lb����TJS�N���Y��.��f�9l���� ��vM��cq�0���jeO����-���&c��R����v�1|���M{��'�1m޶�)��{���e�4�/y|`tڳl0֬w��D�:.$AC�c�U�=�T��������B�@�AMDC�Ta����u��=�n��*����7͍H�f�RO��ĵQ�`���S��Ҝr3�&j���6����T9!Q��G�<sB�6.׊� C;�@t�?|:�JG�]G�\����uL��/�+,"�D�c{��A��qt����3�e��g� �!U/t�P�D�7����!�����~�uW�^su[*�M)b�#b�Ʃ�$��]�6�n�l
�g�RZ��*�<A���C$�6����Ք��Y"N�Rs��n���Ua�"R��T�d2�4�_�}҇5�qm}�Y�ѻLx0�SrPȥV��z�|����M�YK�6�Lq��:������粪��Hz=7���Q�al�6҅��MJn�g��t
��:j�8z<?#D�cb���T�C5 	e+2�N�ws:�)^��c̖���:>}�=5������|���z�~���Iɘ�i�3nUr}(.�b�/1w��ˬ�g;�κ�u�NC�F��S4�l��
�#���;"��'�I��;L춭1�t��Ne�߲�/p��t3�{�9�u�w��$��k��C�<2�	 ��6�;�߬�=h {�jƈ�g����I	�@�$�Oa~����z�=�^59�+�����s}�y�(���}xb4�Me]���5� ��ӽ���������'��Ԛ�@_�;���Gx^��m���Iv��]������f����A�|N���PH� �r���$���xxf��Hsm{B��_i��*��p���
�׸�[��]�u���A�)��`Q֝�����v�쨂X�%Ȅ;������
"�D� ��C�ܾ TAuY��ō�V7����H6��Q�@�z�3>�!�ni�,�o/% %kv��ژ�l��D7z�����=�x�Y'U�E2����-Y:%@~���!T|�:}^�Ƙ^n��0x�-�1_k�c�>a���ߥ>���p^ٝkr`+ͻۮÊ/��(X�>a����1�t�]�"(�p�d�L�jޑQ)�Xv<_���\�l�{�Wf������H�)�m�a�
�Lױ���; 1F�*n^DH�7§���cL�ǒ��7�f����{4��=�&�H�'1���n��H�^cL��Däd��uk��N��`H}dF�ر�����YZ�]����#��&� �\B����w��v��6����2��֥��]fb�(�'�u+������h�q�{��e?����mY�G�c
RL!e����~t���!t5,5i���$!m�ZY�a<dp�y7�~YS����������W$���^	���9�^�d�o� ��!z�BNT�DF{g��L��؏f9R�QQe�/�|��{�}���Bo�]ԁ��3���C䄦}w���?ō5#���g�=��C:쮻��U��Op[^$�f���+�*�m�^�=�H̓�@��S�'F���_�,�ݫ5Oq��)���G��9,�q��E�=�ݣ7�`{ۡ_u滮/��qᛲ�="o�ԉ��h!�t�^}0���UUz�`���OʙZ�$�W�������U(]E8���S�qo0�/�}Mn���	:Q|$��d��b��@��l�QO����'kpQ� �(�ɛ�����Z^��
"E.�1�~�~���J|�}�{䷝���}�n�=q.g�1�=K�,�6�I$���Tɮ���C	�gG��y�n���F�w�1�y`�M���|�aF�A/μ吝����\S]0K�k=c�xlޡ����"+���B���HP�O��c��Ӷ�?x�G�s;��e�:���燭Y�i��k4ޛ`��^xW����6��>D���yBwUN��n�>�rȇid��UN�s��R�5�G�1�:�*�V�Z/ʢr��x0]�]���ϫ`��cJ����\������´K�A��>?#I%��?H6���O �ˇh=�s�"
i_Wa-F�+�*������ll�(�a����~���dw73ۧԳ]�V�<_��oH]��k3S�͚����P�䈬�S�:{AW�I��:��{��EMȰ�@������b��P��>.Ȕ���HjcZ�BV�)3�����KE�m!؄�g��v���c�� Q)}ݱ<�7�cU�1�}��U
�uk~?�!�p�ɖ̌�)���{>߹NN�UۃWd�x�+@٩d�|�g���;�[e(Mj�e낚޾���J�`ٶWge�k���}'YYzy�	�Ce7lK���΍�9�,=���L�g|J��|���xR�TƉ̰�������栊�!g(s�R��}��}�<�l�۳��Su7�e<0+�5ISd�|�(>�^�^g��q�Q=^�%_� �����mS�Z��m���<#�����A#�=%SN7&u2��_�h(��d���f.D�-=��M{�O�"7r�Y�x(9p�7�D6rH4�$pﷴԴ��օO�RG��x�Ր1ЖYhx��g���O=�ㆵE>pE=Ɔ�eTf�<.��Y-�h{���]Y�y��?�y��P���?�f\<��{V����T�Re>�`�����Z�HЙ�5 ��)��nee4��C�����r�.���j�bm�|l��nFPC1�b���,5���	J_���@�)�6�r�ҰcZ4D}�X��~���!�l���Wm�븱��=�F���5�W!��)c�����}Rӕ6���6�W�:�zZ>D!��ޙ k9�b�]���M1u{��*n@��u�َ�:��g?3W[��M:ru]����!��2گk�#�ϋ3? Wǽ�R���E��p�H2y,6�������UE�e�SЩ�Q)^�1=b�O�b�jZ�1#&�`����r�-� ӱ�b�Cy�O�u�_5��D�·��)�uN��̃�����,����9fmC֘�7m��R�P��h�Jl��[�rr�8%|���ű^N���C9�m�|�Z�W֩����[�|r�[���d�I!�|:�$�=�M�f/�l� ��s֮�]△��9��N|��"hh=@y����;��$�hf�H����7��lG䚹��u8yH�"�[�{�'�4�\��ʱ�8��|>��{Jd��[��� ��L�����;<���E���j/(�=y~�B���u@�EM�D���Mk�U�}碉�!��<q�I5�2m��Z�?�|�]��b}lw!���(&���J�S��jL3]I�����.��ə4�<�"r~�X�HS��(x��j^N��1����u�xW^_�a>o�.Z��8ҙ_S�ԍ �>�>n�W����}� B��|>���"���@�uW0������*ݴ2fOR�T��@���џ!���1��6�ȉ<��6��vK˘|u-^���L"�w�y>;Y���hw��|��N��ٸ
V	N����ӟ��4���������k�e�'<;��~�뻪��q�n��D��> ����|�(�4�m�HG�v��]�G���0�E�6�-��X}�
�|��/�_�eS�i�}�ݜ��ѿ^�G�VM��SA�Q�DSF/�|+t��w=�7��}>����T�}A�JRYN�eI��3#"��lȘ�:Υ�'���gv�YF��3,(�퉋&8yn�T��j.&���ʚ_:�]�0����<��1�R�c�WǷ��3�L� ��K,�o1n��*T/w���C�Z�v��9LM�S/NY��Lut@$ ]6F��ު9{DY�WR;�;+��C�$�+v�?�/����9g�L����4G��B��.j߼�Ǵ�.�"������x���]����u�4)�.�;�ܥ4���q�7ػ��nT���T��p��W��{K۾d�{��cE�����A
a�ZՃ�eE�Q_��P)�ᘖ���y�(t�t�>m�l����m�Ey�}���n�b&8��7����B�)�yM��.F0yMﻺd�7bz��sR��J1B�}_d'f�,�&Rb�w�o(e���h�}�E��-��b��)���$�ژ�fC����V�#1��IWj����8: �T}s�9/[�B�n�\�r������ˬ�"�~͘618���T���b���.�^˃e<���M=L�Y8�V�f(�j��r�%�.�13/b��r�����&�&�+��Rw�iP3�j;��Ƨ8��������2�'-�q���u�_`�n�5�g8jXs�M�2uѹ��'C�
P[�N��L�5���0u��aM]Qk�{KNw��$���s��N��)�`[s�٫��;�C��kѿM��{]���H��c���w� BL�:�`�XOճ���l�2��"x:PʝUnWuL�(���⌣���a��z��"�����;(w"��o��M�[�]���*;(n�X�Нf�uս�ob��zEw_�9�d��h�.�����e�{!�{�^>F�e�\�K�f���$-�5y7�W�r!>��:���N�x��QV�'ryTL헡��v���=�J�C���ۀ��1����N�֙F�v�&9�6l�jI�9`w�GJ�2�$��;M��˻5�cjQ.�����d�d�]�hl��gX�1�L�M���|6��`�ã$$�έ�h�]�f��)DS��n��{�^=��1������ʋ*���Y��mf֋ys��K��gc�A���˛s�G2��qu�G��W�EgΜGK���{o9[Ϋ�8�U;/<;\IKiN\;^�!��,sΣ��%�G�V�& �:���6�V�;�6ʏ���j^��cj�����5ܷ${F��H�a����H��C�X��w`��m
�gz�<�v	��7������vn�����ݲ���p�|�uvl��{�k��35Sk��ڕ�zkX�U2�FWiuM"�6�-lR�D��d^SAg��B��Vp� DקW����tk/�E�P�,J�i��<��N�}����O��i�*�e&XMdr�v�yuБ���s���(���5K�w�����%J���5���=gZ�ʤ�V/������L@�bJ��AL0�~�s����kT6g�Ęʇ�Xi�o�G��o��(̈e,%`��m��ri1��C��L��8�SS{������aG���'�$�X��'�h3=��kT<� �t�Gg��{m�1�Mz�i���6�$���VsŊ.�ef}CL�J�O���g(q<�*i�����c4�	1*O�Q�f����3����k�����x�yP1ٽ�a�� Q�0�?z�SHi���{��O3篻`g�{g�h��M�I\�%b�Sh~2ɶT+
�}�&�X�j���p�I�9i�>�}��I�9pCW��h����AJ���g��1ћO�㾬���=�:��H	+�L��?!���֘~|�t�dZ���,�n�f�b��!��&���3��'��<�Sv�������a������G����GL�����%bͲS�}s/?}��x���Y��J�3���W��;����q��I���LO�՟ݦ&�&�0
��l�?�߮���T�_!�8�I�Z9c�i�CI�Wa�����"H�H�R,����k>g�S�����2M�8�?����y�7���y�������M1�l
0�P��1'\NwY6�l����y=�����c۶}�z�N��YR){����I�S�:&Ш8�����ɉ^���_��H)ǚ�������2��2>�Y�fF��%���w���8��~�˪K��paR�M�ʞ�]nͳ+u�p_�S?^�r������g���6�����l<Of���ئ���@�:�N3i�?3�Xe�B�ѓ�8��{0~��r�lB����5&��|NJ�������#�S�1�ڳ�{�1�>��st���󣻳�R�����I���CN�d�.��Xi�z�'Tq
��`s���)8�U�z�=�ejV�eL������>�]�wP�T��;�b��?"�)|gެ6�+<�v����
�y?I7��x~M��1ө$�]�i�U? o)14/�a�q+��yt�LLd�q'2�I���~���`�����{4��I�%(��su���6�����@�C�=���Ǭ8��ȵ�����?�s��@q
�����:��6�����x��G�h������`����̆��Q�ϳ��C��C��9���n��Xbu��	;���U��?�[����}�����Te�!1�9ݦ~�����=�����r�#72C����1E�d4��=�֣u��f�9'v�(9���'���-tǗ3�9����s�9�Ӯn��r���~����������������)3ԙ���������58É+��r,����{g����F�'~}��W�!��۳I�~M&�6��C��?3�k��6��*k)7�	���?���>���������N��*(���y�<IƤuh���i��T�����`�d��a��`�S���O�Q��1���?{%t�����X~w�_�+��z�־���_��4�M��a��;Ɍ60��O�q�L�`b(q
��8�Gzւ��
��k+��hef;����m�����o�MX����v��p���87��f�|�T��ˮ����/�}���&i?��;���$�֩��L���y��|�XlCYN}쇙�u��i����,4�/p��*M�Ty$?~9�$�c�D�5�C�����:���65�4��/��nW�"�'��?��60�HO��80��j�O��b��Rq�8���P�aԾoY�fĕ?'��`zӆX6�9f�Y4�6��?f�ݐ��6��Ͻ�Mr�5�����?~ϡ�-�������3�m�.��r��>��m����51�Lq����2}���b�0�&� ��LN�jq�+<�=B�H#0I^%���� ��x���`����f��0�}���}��������?+?��fس��$�͌��y�x�Y��q߮:M�YPr�(q�?\I���!�bi��3��·�#��Hc5���k��(u6��
�)�C���k��~��������{������$�16����I�������[�I�?04����ӌXb����f&0�Ҧ?0*�{E7�fߒ���M0��l7Ǜ��B�D4��I�ۉCY�_|mQ�&��?h^�GFS��ǐ�'�~0��N?'��Xu�ۼ����/}f�'�I�]��~�m�����?��1��;a�����:j��~ea���y�	���d��?�0���[g�S��<���f���}��� 0�|�^�����v���=��q����0I̳L���������I���߿~�9�SC�,Y��CHmS������͌������i�'?��e�n�X��~�+~��d�Ԣ�	0�_O�T]ܿ\�]�7��x�\������`�E!
�Q$�w��}��o3���w�M����4h����J���
՜%���8��p�a�R!&�CZm��Փ��df�S��,b�+�l��Q'框.�O'.�*���a�!�u%��}��������oْu��+��3i1���`�� V�/�m�b�����۔k��<ͣ�hw��0	P��wA���H���=�3�Q1�x�c"�Ndw9��3uR�T�����~��i��;�O2i���*As�Q���N3|���̜��`m4�1���0+�8����5�����]2��	.�q�c��/{�M�Ub#�C�J�;'n���>Ɨ�}��!����`������u�T��i��/��5���T���1�A`z\3p�h�,Y�Hm%~N06�͇���&�8ܠ�@�L�/;)�?s�yH\��χ�fE�m^:��;gJ4���`���ҁ3��q�36��j}~a!�#6"�l�G�#��:��S;�]�J�w��q�o�d	Pl��[��x4	����#ѵQ�ǘ�rn��]�2�d�#y(��K�q�����赈O��%Z�v��z���?��?;�� �?�����STy�Z$�skB�c�9��tK��$(\�e��X�[4���a� ��V�����<+�Q�% �`"9�����$�ٷ��z޺�a�?���U�^��ͯc�O^i���U9��2�i�%�#f�!�E�Dy��vgM5��j'��Sz<=�D�f��EY��d���]V���{b.']�N��Y��,h4��ݶ�̃,+gr��x��G�pȋ��γ��
�0���=�/���n�&��̢�V��ZlR�2e4�N�4�2-�`�>��b�����-�Ґ����U�"͐�o���G�&�8O�'�]*�fP�>�+�bD�@6Ȁ�4���{mEAu���"�V� �\�U��B���a�k�m����{ч}����m�|���JB��8-�UܟN�w+4��]Ky�����\�a�W�vP���^����o���7,!��J�_����R=�ޣ1��T:Q`�#�힖�k�G��69Q�6Ǡ����?x|=��j����"R���Y�H���e﷩["�I�7j9KS��DL��C�[Mk�Q~~�0�%AbՖ�kb�����uT�'���~P}JZ�Jcر�a�l����l��� ��{朱��⬙��>�F��׍{<8H��
��Ֆk�sAK!9r\���j�Z�,�*e�ܬٙ'Z+��&�s+g��f�ԇ�I�F̫��z�/=s"h墵�pѸ����%�N�1�vL�v�]�_{3$�*��88�~o��ju��;�d{����<���z�£���HC|ffڎU�kSf�:,���Ql��OKK�#�Mx\&(n(t����;��u�u���,l"=I��eW��kԨQEQl)�[��=��?���~�ar�{!&� ��k�3����{�B�ś��|.*.�V�y���u�#
�@b�s�j���t³��	��*ͮ܊������X^�����3+��^��y�'f��vx��}{n#q%��TG�� �<ئ{"`*�L��&�lV���4��P� ��U�Ӆ�3REN������tݞq<F.}i�N�*�jE俷E�@a��6�ID^J�!�[�TY�"F�3�����q�YR_#��I�r��v�
�v�[ޅ��]]=��������l\���A|P_�f�Ro7Wq�<���r`�螙�K��AxW2�Rfk�cx�pv���!�`%��٥>��IO/l+`oS��QU5���s�]�CR��N�g>�S{�;Nvx|>��k��5��p�;޺���U;�^�N��6����c��w�N	p����{ZI$���<WTQh�C��7�e�w�7G�����)Ȍ%=^��K6j�J�\$Q%4��Ɩ:!�˘�j%�[�������p���Y���%��ywJH�4�~}=�ӷ�|�TMϊY�u��T�^���mVm�b4]����]�i	5�m��qTkp1sQ�]�S�JM|V�v���DI��L����p������]�f�� N��ě���Q%��<�C=�}7EQM�A�Q���-:��F�ecs�ʵ���o��Sλ4��[	�6�5�v�>6:2�,�̟UN�kf�t��	�r��b�B>���-��'�߾�Wx��W~DK��3�4AH6�<������u>��������$��7a=+�;���S��t�[�{�����
��z2uH>jce\���+0��5�-?��ě�+���O�Y[�*"��)C�A��V@>
b��q�S�E5��Ȃ�;��j`A��'=�0�D��ۻ�y�}(/O̻f�m�����;�j��M�"�[���[�~�f��$�^nX�M��9|�uAsc�}%�vz���{�Z��ռ�t�������`��R"�i~w���׹��\���o���LuW��y�{6a��<l�nź��;h=�،Jy[
��y����]�cT���4�i��~�5}�Ŷ�9��]T�X4�ُy�8�Ɩ=>z�ѷ9�Φ�.=ܗq;ӀS-ҷ[LcTz�>�6�o�mYޢ���б���1��Z/lծ�Vn]f�G�c�$k���{�N����ns��5�e~9?$�p��:\�ǈ]���P�iw�i��;�q����>����)d�ފ�9�]P�S���n���a?�}�9�m�hM�.B�T��L�]uM��"���D�]lt�F=�lU�����k�t6��F�`r(�ww:���.\P��2%
��䂜�#e���w�CE�b���'D'��;q��2��%
�$�|ujP�uUr�}}+r6���g9G/hP�=��,�I�_y��)k���Nz&gD�ڊ��O�ӱ��*g�`p��]Ƞ��C[<���h�
L�?� $����Ȕ�$|�`//K�vt=m��˝�uV��*�L�s2�
{���g���
�V�/�莉Gg�������������#n|T���W!s.-�[��e)5BC��I(�ΚKBZSP�y��������*u;ԗ����]8�H&�b�#e'R(���}Ll�����D��z��vlC�{0S?c��0�ꄆpκ�iivfJ�W�:�5�2�̖:��;�X6��kF듴�&�T�]�w��=����/��,��7z�i=S�CkO���Z,�(�-�JGF���~�v�����+v01h#2Q��Q��D�Нr�l�I����J�mb`s��z����"J�_<E���p�m�=���n^��5�=��ﲆ��A#F����͚�D[��WԍutQ�2V�Ӳ��_�mDs�X{��f&�XD�M�w%�\�לzPY}p�[ҧz���M�_���{!�� W�-fk�Z��"��~��DO�|��TE~ɹ�(Ѓ���`�(����%��c9!�ARq�G*0��Fr9C�8�M�<�=2pz��l�Q���TX�]��P�T��Ǉ�ĵ������P�P��Ѳ����a��u?+�2z~���O�B���E��$�GuC�"A0e�v`�d��Ua���Y�i���.��C��]�5Cͦ�Q/z����L� aC���QW�1�{�ڨv���S�hbU��)�'fص��|�-�'\�'I�O�KM%MԞ��כ��s�תX6m�xPAtj�߃����K�:U�l���$�C��J�������m�N�ܕ6ߚ��h{ȍg���UL���b!�%��w(�7�n�֙�s<�=.�"���"]�Z�w>^=�W+��pw�Qrɏ?Pc��	�Bc�"#�X̸���L�,��>�J�l�jC��vh�{�q��SM�[Y.H�`�(W3�ʿ�������lZ
�&�j��yi��8M�7���Y�Us�_C��d���"o�שy�}:�����iٺ3?�2c@�ڻ�wjV8 8���\$��M��B��g��ozд��h���2��_+!��lNm0�]�ȍ�M8W>��yVd�pĪ�KC�v�z�V;�2�������⯉����J��[����+�8�h��K��������;���w=˵�6-K�k�u*�]���vY*���>�v��,Վ���a�fΫ�?��ҢDi�f�V6��Yd�M��<��/3�K[���T9n�Vl����p�6Ů�Ҹ��T�W���xN�O ��M�sqI���l*@���.~�-޷d���bf���Kv	��:'��'�L�2jI=k�(��)�7��xB�j���<b�	��C�b)?t�WsEL��xC<L=�2�;��x8� m�$g`�]31P���=���ӵ�eA�/��I�ϵ"�;�
�;�K��x��G�ō���(p�v���Թ��ڼW��@�nЪM�#w�_�F�c<�v��61+]��|���3WR�=n�� Ln�f����1x\���d��	:��0���GK5���Co��l"۴^�,�H��\���pi����\�E��*p/$�L�� �)<�RY�I.����| Y��N;��H�}���T˾�M�^�"�ܘ~�|�}
 c5�ELt�k���B+���C��C�ݓ��8�n̰��S��8�����+A┄!c��f3r�kf<����
� �?HɹsSc�J׾�����}��@�����:�X��Շ@�L�g���Hq�u��+��p�����D���#���J�;N�����N����V�:!�˿��puWon}��(���G���sWNk/�z|*�b���b[�������wIa���R��I���/�\���")��K�}��8�l��K��ּ�~�/9���}�e��D��A��!�>0�8T�t�-��뭃��m�������b�hP���U��(0�يdu���|�d�5�C�1��c��]uvv��=�U��\-��ڬ�9ҁ�$��خ�m�T��osՕ8+�L��"���X���N�2=L,xP�ק��v>+WP�U����ۯ�[��������w��o)�Ƴ���{c$bR$YY1;	U���9���)g�0_�`w��>��e�ڪ]Ŏ=��1(9�`Aꪬ�k�Z���y
	�~����=V�I�?���,���Y~��I�ޭ���{�u�����f2�h�� iX�B�d׮	tI�8�W�%%̉H�t��E�ل)��c��$�f��۴;��]|�l�ٻi��y��!/��k�A�����"sDd���'F{�q'�)���&gB�T�Ϊ¶�f5M�:Ǥ�89��D�vu�6'���k�.�gF����P\�A�@%��Ӯ����DT9i�|}�H\�~B&<[��7�xh��&m{ܬ��~����������v����\L�ː�<zy�^j�g�`.��s=yu�7�@����^qW4��d�2�+x:�D��B��o�tz)ޟuؚ|���e�:g4]��9'���;Ք��u:B����L�r�5T��S�F�.8��ꖸw��]y,��X�v'����͑;.���.8��!�C�}�N�1<�J+VghRA:�T�#WgG��A��~�����qy��.���-���z��P�����~Z�����-�����˄3U������B�T�*��2���
UuW4͘n޸�rL�R�Q�Tņ����)ϰ�t�̵A�\�ülS���qc� yv��=�8�����iz{�6��V�����5�U��������TP��ż�Q8����kģ�H��=`��(�[���s�]��-|�h���d�k�MP�;Ǿ��ә=�.��������a�
��M�f�k���s�_f���
����$���\��`�!��=��0ߩw���r"{�Ő���y��b��.ggM��$[�T�����r���B�qG��b����#���A&�S��[�i�mN@g�<�x��F��~�Fq�k�u�?�=ʥ����� �n�m�xC��+N��r�#.�3�)�o���%�ڣ�m8�(��L��ިb��>��\��Y�z������Gf�A���{މY��Cs2~�g�`<�{�ts̈́�I\E���o{�Փ	gkdE;�ȊO���3	Zp�I~#Q���UT�S�x�{0*k��q!"f�}'w�d]����xb���q���6�ݹ>�)�B5Ǝ�y�=���F'��ѩj�fx x�xv�~y��`��._�N��V�A礂�_Qe�O��D%��r���8��V+�4_t��DQ�`���ߢh/�!����%$%�*a���9�2��J��A ����g*�������b��V�!W��[�wU*�W,0N�f��Uc@|��p&��9X?{%�&ƎT�	����!��T�͎����h����6�Gw[*��s(f��;��N�n�iC}ufump��A�N֜�U�^u���vq(R�)���΂���8֚\�0�ϟ�������g
�K2;�64�q�x}�r<�PM�3����^*.'�iM ����tD����3!�ՒY���8S;�G��}E��<ب����7��w)/b�Bf���塨��:ޒf!M��H�]��!���
f�]�/�#�C
�j�u���dޕx1�f�NL����	;z]q`������;,<6��O	�ݼ�V�fQ(����k�Ԫ�"���v�*�JA`B�B-������QE Q@���Y����䳅��͡����c�YvҠ8a�@�&��*tO����z`n0��@vS�J�7E�b��	$������d?;��x3jT�e���+������>P���(`r�8�l���[��ǣ9fV�*���!�i�� �Hd�R(b��0i�%X�)���T;�
���*��j�����x1^L�R��\/5��T��q8�;��:�ٲ��E;7jb:�²|b���F��)V�4��T�Zw�AG�;���w�����_A�H�2Fnb���	2λ7&�a�xq��%[�Y�4�Hr�wF���0�'r؏H���s
�[c��u[�V�n�c�¶ɔ# #m����#&���b�n�f�����U�/�)����Y�M����ב�$�D9uШ��C��H[�RgMͳf���0��Y���ۂ��(IK'Y"�-�ra���,j{5����,~���m�I;�I��\��󾣏&�<`pO����3����3���6]�M��d)lJ�)�G���T����ת�8jP��!���u"��E�z(<Z�Ո��>�&�p��s3�m�D��γ4���ønq���S[e֒�[D�DZ�������
=��.���l�[����˙{9D1����Nd�)ٹ��=����=�w�1�D�|�e�Ԃ�,
��7g�z��y����:��"��K`���\��
~�7wYe�DM�Z�M��kP��A��	��5�&-�.C5Q�9(�)�w]κ��f�\5�Y�'�)�Z�x��Pq�z�&.H�uҡ�-��Ubr�k5%���4��8y.UƄ̼�L�|��/{Q�=�B��r;�+�K�?�3��t���b�{��Ā��+��9װ�k��S
�&^����,}�¦X:u�[Bq�4e��aV�e];c2�#����!���`����t�;�X��Pi�5Vb��v0��6��8��9Q�5X�NN�E�8U����Eϳ!�2�eGf�V�=vbaMҟJ���>,C� �s�~�̈́�g#E���^�P90tҖ�T����%��OwU���M�q_[�Y���+6�ڵj���24S{�I���Μj�s��n�,���}�d������8/iXz�괮���v���=�j�!Y3��Tt�ir���{� FKM��'sU���fJl�H��V��]���<|��WV�����.G:�u6��0Wp�Q�.e�3�epB��ͤ븳���O�#謉����F��)FZ8�j����Ğ1> �d��)Q	��x~t�a��U�].��荞W	H�ި��T�d%�ĺ�"h��w�U-̽t�A��`.'��0�'N�fm��[���n�xm�F�z.�J+%b�HI���f �#!"d�L 8k���2��h�m( ��Ξ�J�g���eC�j����5��k� �`�p��I����淤C�TTŎ=y
MĆ�����w��Q�Qx�j�݌�>@�RV*��d����G�k����va��1�I��~=��W� �8/H&�vC��Ս��7~ҽ�'s�W#�� '�7[q�`�-it����%tþ�P�
>��"�D�I�gpExz[C��][V���� �/�oT����'P�ZC(��(�EI�.�Ѣ{�P���-�R���E�r���|*��p|檷�Lm����Qx��$k���Z���u�k[�	�MhƝ�;��ki�߼�8��0)-�蔰��2�.����D�j3������Nj��J��çߌ��S\@�ɇ���0�M���*��}�3O�4C��̢F{�r�����2�$v=�x� � ?S�N���TQ�ail<e�>h�������cl�e?���0?e�"#A�D[�n�֦��B��`b��P����"$�!$����Xw!��IX�-����GPJ���f�Cݭu��lZ���ޔM�&v��%�X�)��f'Xr�8�5�V�>�[�Vc�Fړ���ݧ�&�C���ۓ/-��`��tF�TG9��O�1�w�aO��$8�z�i����&�_:b��#S�l��a*�g��F6�uP���H=���8ந���X����v�Æ��L[�8i )���g,��C�>����[�����as�cg���RkgC��z��Uj)��ʔ��E���28�~�W�ޒ��iWD��$����w�1�K4
�_�nz�׉y�Q���.�q.w�3�&�=3E×�q}�k!�D���3]F�A�擋G��qH��1_��XA5�3!��`C�v.	����h� ��z�m1�F���v%:o2�;��|m/�\����9�3�\)t4�*�v{͆�`�U��-�K��8�"G]yRo���p[�w{p')���&!�����у˽�����	WUH P_��TDUa�Ŷ�~��|����_�����$�\�o^m���t�~�U�o"��`�s�	��	ߪ��3�3�TFl*��(�#������r�;T�"/w�V�=J{�X`����NFVО[������ҥ��'���>�׍Y��dz�Q����;Ю"�# ��V�1�S�ºs:��_/�Ug�'�	10[k4�;�-#d�4	���7��t�T�!cI?O�m_��p��߈��VM��ɷ秡�٪�	]�wX�H$�)~����P���� ����m"��]1h�O�u�ORθ���v�s;]���Ln�ˆ.��]z�BF�Y�MF��}u�s>����6�f�!wׇ3�;ן����(@_ɀ�ػ�� !W�IΔ���T.��I�I�|��D
�Y3�؆<T5<��[T�m��u��p�6=���Ǐ�qz�2�^��6q��p�w�PIzn�I��7�z}�9���jم�Ƹ �B��`S�cB!=��y\�;n�ta|`�I@���ҥ0��	�Æ߷�~�r�#�F�>�l�0z����Mn�A�7h��j]Fqe2Q����CЇ|���nL�r�QH�땻]��-1�Ǿt{*�"�F�-b���G=B'C��6QQ	��?۫4�����]�����Z7�Bۊ�N{W�a;s���� i������}�o��!sv��f�:f��_�������|����t��;_L�忴e}�Q)��w�,���V��؅�זD�cأ�y15w�NߪG���r'��z۹��suFOw�u����Nn�L�8��V�$q� $x&�%3^p0��l�j2�����նO���B#!��Z��pUmdv��T��%=��2��Q������rk̼e'�HS�ҙ��C5wM�Gv�����o��	Y��}��/�l�;������E�����&)zO=���j�$��uA5��j^��v*�����[o.3pK��j��iB�a��s���Z֣��8�̐�v:1�fh�l)	Fn_��Ǯ���}��wu�/��?�I,��:ǞP�ɛy��}0�4bFU��ݡ���}�g�\;6C7��y;�<8�h�:���ߎ^+�U�ޮ��@^��C�g��b�efF%�_O�X���͸Lۏ;/���^��īF�RN�]���zzc�/�rb�SR�p/�ذ<�5���=h�V'ş��[���k���b=ޟ�Bbs��↬]/��q��ʻ�w/X�Jz�]�5�4z=��مr���v���� \��%�~3/�1m����%Ps�
��[� ��&Jj���I��f�hY>�s�˄�e����c˿yvZ�������b��t{L(���s퉉�(*�#���8��L�O"��P��$�B���>���S}u�6�5��먹V�D^EK�^G�>�Ck�Ә$����LmW�a�W2	:�k������� W�G	V3�N+���%��}ב���ܿlÏ��T��{>�����]ys]����������^Hkև��n'_Gi���Qn���'Y�.S-�%Mg��H_��z-�����F�rP��BR�w.}��\>)��^��Y�����+�!U!P��h�Zn��N1q����}G����$��D�c.3�>tIPQ+��[۷�c�"�j���N�yKd�n\1Ʀf1hV,�@YDi5����~.�{{;��F�0i���_[W-.�7��Z��[������U�[�����GVl�Vkt�=[تb�^g\d"z4���47]�vo9@՗�x�O;��he��y2P��h���+�א�s�c����~�����W�} ^�l�td�[Н�dIbMWmA␉+�T ��ݒ��H��Gb���{ЏA�<�D>����3��y=�����u��{e,�ac4=>�i�k�y~V2W-�/���f֡���\�trŨ���wV��W�e~����i�u�KѤpب�C���}�3���)`[6�k=�{�6h$V�͗	*�S��~�Z�ꬴ:c
蹃�d�������0,�D�`��g��p!��s��w-�A�Y�PEv�Шknt��
W�+��@�x��ɦ�\��j�O���8�I1�;ޏq謋�fxs�c�6�`5�f�mW6rv�^&$�%���!��0������{$U4,�eP�>��b��(X����zC����n�4h�j2.$w�\r���-�������_��U}�j_��~2w�J�i#+'��d���Z�B�f�ڰ{�H�>�dÎw����gW�'o�TM�+�9/7�-� #�~�ws�`�{�����7f%_2�>�V1c.�]��~�t� D��9v�����/�/�X�:O��]u�^J��^O���Ɇ�����mʄbLV��Aܮ�|��d�VwU�|�!z�`�ۭj�w9�<�<���	�u>�J=�c����<ҹ� .~;��B�G���{����rK^�Ut���[�n#����\J���z�j֋�4kɆl���J�pf�݅����*�Xk�h�GaP����@��0�<����T�]dLh���V Q���{!���5:��&����k�\Iqm�KL7\�,5׫�QDV7c��\�e���
�A�^צre�c����eU�ϙ?E�r�F���~� �w���/��^E)�sT� ��r�����2Ͻ�ju�v0�Ka���q\�O3H�����1hOX�m{ؒJݹOٙp�C�-T�Tq��Ǉ��K{�0�T�<�B�Ҡ=���b1�*�^�<H:���E����ݿ))QU{��T�Ec����28Dq�x�eE��Y�7R�s�6�a��ЃS^��q�zgq_�Yz �glw�E�kf�������/"������3��ߪ�����%ޖ|o#�>[ǘۜ��,{��=4�:�������a�6�/h�À�g�5�w��ꋷ/�p��K��Ҏo����ҟ^X�9���E��i�/C�}��]���?C�ފ��LB0%�t�Ơ�D�`4Ie ~G����JP뼪i��o�0��Xx�U����f�:���:����=Z���==�Q�o�Q�SZ�Q��%m��R#��j :�0���q�goe��4q����q�w;��~vv�'N��0�ấ�RnH��p��^��[#b0�L�d�2Dn��7��}}�~���� �XQ��A �>�T�<��I*��/~��FI#\�uN��L.��r��F�n�w���/`�tD
b�etF:B)ܜ|UU�J�*}�d)���C�����R�[Z�z�gj �;��{����e७%�����=6�1n�����"��'���~�]���:�v��1��ѻ�6</NH��L�/;ڮ��? "0[��wu�K�[�C���y>��}YM��~�������b�fZ����b�O,�7�F���i��B\��\W��uk�[j��U��.1���7��/t=���ӫ�{�	��h�TE=m��ϝz�bo�~>�7�K��,
gC<�g�Jy�ϕ)@p��l�D6��2k��D<�Q��>��5�~t�ޓqH��r�m�8G1��|Q��SJ�[��eR��!����^�Ջ� ��H�Ge�h53k4mt��帎������}y�N�����^����3�x��n�`m��%���2d2EK������K
��=��إ�y>��z�U���G��9���o7���堔��w�`<�ڴ��s?�����ߋ�����ve�I8��v��9��3���u�y��»��kyg�,b�n�/��k~�<�v�,�k4����ټ��u 哮SL�< ���[�t?K'y�>XOWNr�7rh���v��o%��UG=�(�GI�1 Vu\�[�p���3t���4M×�)'Q�gR�{�~�v!�q�G�=c�C���9����T
5��k{���qa�y�[y+v���gm�y��9�r��� ��������-�|�ڙ���t�*����{nzn�<ŸĴ������'��zu2}�"����VlH�dYSz�t��q�3���X�ٮ��ߓJ��{��at2B���������3,��L�ϥr�/y挻��Z �����d��@W}5w�^�5�Řg�=*�\)ɟ�V�9�At@�o��a/R�1 ����!�iMV����߾�:����",x�ԁtL�K�׈!�К��iOOyB�x���%�M�M*��ۗ�����=?�~L=��uޟ�$Qv�8�^$D��.G��h`���<�7�}��#
�M3A���1ڟ%^�-VO��Y0t�S���*8�5��Yy 3��	�K{����ʘ�J�y�yL{���]��3�"ɾ���Sd�+FJ���F�Θ_VFOd��n���8���<�Yh�^q���V�oi�7?֮zOwu���z?Q�0�;ү+����% ��"~���sK�7Ti�˟�E��=1iy\0��"����;u7��D�@��,���&"�z��(��Y�r���}4b�X�＃u��"f;�Kb�{ #\�������;n���{�lm̳��M�a�7�5etAКz"~�;�*�.,�(��uq5��q�o��b��6��K/>ъ.ġ+T��W�KY��S���� �H�&"|z'�r�D���ت.��:#.�@ /iwd�	j�b�UJFi/e2�U.۶#�VE�j8�qT��t�\V�A��3�pzsn^��q��RQ'Gh��Qr��m��m̞���>~����9sџi�*�H��n��ӏ6��.�t;8)U���[����������T��豇�Ѷg+P{��yF��3�����|�<<Xv_���"�Z�-{l��O��Ȑ��m������vc#OGT�qy��7�� �QJ'9֢�.ѓFnO��*\ko=}�ڳQ�1�:%!;u.չ �^| ;^=DD���()�
�Om$�ʏ�7��w��e5�9˭{�k�7�������B�ȅhϛ�S"�A�[,`�]3Ƿ4�5�d�i[��{��۰]���Px�v��h�,պ�k��WT�wfM4�
�H���ڔ��������t��ef��u��t0��ŧvw2mr��^�zh����KsV4�Cn����O>�xC�R�"L-Ys��쨰NƁ효s�5�b��"_e�Y1]�����5��h�±AT�b��"X�Ppd1)�iS�KW����U�Ų�#�'/��OI��H�r(�Y�5E3c���c.� ��륥�˺��u�xf��c���c��~�R����'�{##��1ǋ��D?���zI���Kz�B��}���?(��H�~݌TM��q0bj5���m��is�=�S���ǋ4�t+�xS��Ã�z�E���k��,u\W�Ӿ��Ú����H��ҩ�K�k�+�����xpe�)�4���Y�B����<w�[�k�ܾ�޽	�����{�6'���?C����"�]z�MOҴ8�/zQ-����;w��/[�^~z��$��<��&����s+�=S�?tj{�<�m]�
WW���$��}�� �	 ��%��vI����kLǜL5�3���mX��}���c�u
p�P5�a��|]]F&pT�0�\�� Έ��
�7)��n�ĕe*���:���u�x�Vq�mr�~5gb���v���n��WRt�M�x2��u��"���S����G�Op�Ikh]��Y&�vN+cCw/����� �1FX�{�4r�e������9�G��ګîh@�9����y������v���DmH�f�?�8�αu��ʗ��u;�s���'A�Nu��b��1qZ8u1�U<	A�x��*е�ΐ��������l]�t�Cc�v��ҿgMI`���Ï�*���m��E�:?;�˗�tU�4�v]p=� �v��j>�>O�G0��z�{��79�}�����Ysi��?�M\��h\�g0n�/r��m��N{�0��欫��DbPSkF��j?׹�����]b�q�7c����ھ�&K�#c>i��7hђeK31s5/�F}�����o��0D!���Y=sמ������U�:�[sl�{gS���8�$F!���hD�vTI��2ZJ�J� UF���ͨV!k��e�I�Pe��>i�Q�3��Mj�.�4���sM��+��L�R�K�ْS륧�K�����Y&X��8�v��T%䣜yZEE������gPå�m���4�혷w��=Ee����3��O�K�����y:��gS��-�2�(�T���T�cZ�o�O��٦��K0�N�#r;X7E��d7��p���:)��6�I үr��n�u�zz���A���}�,<��s�&�C��|��h3mcd^���ֶ�>U��4�	zyW*3r��f��HK.^q���F:��u�ys��䫜�7mI=�z���׹Wj�i4=��h������BƲէ�i�^U��T�2-��wP`���v��T�b/�!�8b�E^�\���S=��2��CB�a�\Ʃ�3�e�kG��ݫ�T��eٱ�e�G
����/1^��Fܝ���ym�6ԙ��zF��:w<��6f���#�̸V����;�X^��sb>�c(W%�q�C�o�m��.�r��1n�7L�s5���q|{sM8�ծ��4�"�k:����2)-�z$3�ö�ɖ���d�
�y�8�w�:��?P7��t
�J����T��t�+cCZ�w{��Z'�r�Ռ�/��P��	κ[�;��H7H�O5t�n�qv���G6:��{�g�Z�Kt���w�*��%ذ�@�Qrщ<X2��]X�Q�����j��Y7�÷g�ѱ+ZF3�-�ê5��&h�H,M�z�WY֧3��2��$�pna�pb�xz��*��oE� �o����nuf�C Y�o<���NH=�����Z;�co�mgKyw��7�T�Y>�_Y(\{:�4o6���M%(�Q񗢎�����M��������{�q�hE�i���g2���k7�D3�)8���X�����jP=w}�+�`;���v=���FFb�()MX�
����O�=:lM��:����L�4~$)
'�I����ץ�\ÜpKw�Q'��O�ջ]S!�ċ��M�mQ���`���nk�g����C�\ۼ�M7���A����g�c�TZ����\0����oiq��jN���p�4̔XT�Z����9���],d��w=�����U�.}>�6�R�:X2����bI\�c!w�m0�����>'�7sJ�WF8t�w��y���t^���j��	�i]�\M��YQR{3�ߠ�<��l͟eE7���Q�W3�5�f�K0�^�N6hiP��GA7�V�/��LԴ2�J���u��$���7�ʢ�Y��[q������p{�EJ�;/���C*B���Ӯ�O�\��V�{����l-�M�TNp�?����cU�y�
M�5]�n�(mX�G����T"G���0��+�S'Mg��]�D~��Cz�q�t}�Ҏ^�̟2�q���Q�5������x*��k��8π=�K��ѵSѱg<T��˭�����Y��b�t�����De}��r�Tz  ���9h ,
�f���{̽ۙ�5��I�\nH6gp��#Fm�ޙ����A���BÓ��㓊�����#�gZ�˶�p�����f\:�m����=}Y��Z�N�ݣ\=.T.e��os����ǹ0eE>��Y�9��!j�ݏ{cy�/a���!�Y�(m}�����b�1��qv�^蚄^={��D����}��ڢ�♢
.�b��X��͕���j�.����/����{��[:���:2w&�J*d[K| �܋���1���-D��&)A6*��[3�랛���h��B�e�ʲ�Bս��"0��|���w�ʇ(��i��R�1�ݚ�9����s�nC������l�5t{z�ϯ��.J*�rD0L�N�t�����V��B�8���Q �#4�Z����Z�`�/���v�X[�a�=��J�^}����.�t����w��=��0�]���ff�\�%�@�ZM!Q�N$+C+}ݘ}(������/�3q���ރ�<�j��e�I��wu�j����6 F�����!�VoW�B���s��ύ�.<O�=�jg��h9m~;���ŷ�0�����WI�16�Z�+P� �͊~���51��`Ó�(p� >�R���5M;!a������p�h��W2
����.d&[[��h��/�o~���ZFʎc�����wp�ٜ�)��ō�o�oF�V���0E;R2�����@�$��Wql��%�n��YL^��J��i:t�ّ)�j���m7w)�����Ӓ�@���t���;9$��;i�z�7[��#n�X��	�&89�Crg���V���w{	�C�~�(�)#��U���ߖƏ���#�,kH�<[X]�� ���Қz��<�D)�9S�d��
^���VJb���y[M��ڸ_���T��>�s���C�j�o����p��N�����Q��HTs���?}m��{��c�ҷ �L��C�.�E8�*C�0��f�A$T��e`�(eת���0r<�z�-hk���@ݶgJ�1�r$��l�s	�>7��j��K�����*�ם�e�<�i���C�T�̂I#�d��l�]o�޷9�9z]b�p8#7\9��H���Z]�c���.�A����y��y� h�n�}�7��t�\���I��S�R�9���⑂���oԑ�Ix��)PI.;���Q5��٨v���Q�ݦ�vg8�FEѧ"Fp򞰛�|� �@�=^E��^�*��C2U���3<%�ɉ���m	6B.��9A�mAJ��Mq�+)]jV.�]n]�H�l�$_�_����d��C�|L��Ew_����y��L`�X�54����&��\� �j�KF:Kɢ�A�QP�W�uje�\N �e���$-l���՛1Y�m.lu���3wע� '�zK�m�+�O��fX��=���J��U���#�7��
��昿k+8G���1g���3�L;���׃�����j=��f�NW����x���j�~]hZ-'�Z�K�<wϦ��T�ѣU�8K�K��s1R�:��Uib=��l���X5qOծ�y��`�A�Y9У+jO���\�	J�����\��5���Go���0Z_��}�����7��ٳ�6*>�u,eWC�ӭ����;qW�P�/���_Y�Ε��`�=)�����Ѯ'
����C�B���r�ϱ��s'ߺV�co�y��e�"�VM��{e��I �
#/�V���[#s�}S�oL�V_S.y�l�G\UM�ˎ�7&��;=3�?k�%s���S`��J}̇jZ�V�j��rc.m�dKƯ_�x01���48�'������ ���1똂g�i�-|SЩ���ib�0x�)�B�j�&]���ӓpr#3r$N�����ůj���]'�k�6D�$]m�>v��r^-\�(�r#��6 ����m�a���i���Uv|7�iά	z�a���y��������9,%�z��� D7� HJ��/��ܝ��7/�=#v�z��3˵�NIG!ac鴦�mt�Z�x�j�n�^T��2����u]E���m���C.�sdk=k_-�Fu57'wt�����2=�v����<16k���)Gʃ��E�|=��^�:��?�� l�;�
s�&7�w�rmx,_��*N�>qWtjpUKVm����	���xz)���}��w�)��mU���������6e�@S���x�t�DC@s]��ٻ	�VܻW�3'ofI��J��J*t��iI��yg���[�����0��T��H_VA���cZ���('��x�2~�'�p��7݃79Ak��ؗ�o������wuLL�{N��Ď�ue^�����8:�ۘ���oU�X�=��t���Aj�NI��߈'so,a쩵���� Y��!S%/{�� DZ����]fX2=T�D������L������#%r�-�ׄ����-k������7ǧ�r6X�����A����߂ x�O��1�]����˳�:ݙ���(/����۾Ε?��2�t�w7�[���X�� ����O�B�[�;�#mGEG��x�̀�(�^�q"맨Nu�I��\%��ޫ"V>�7�RoԼzㅀ�R�+�TU"��|�����y;�az�a��Zrb�O��7��5��,�Aj�ID��D��	��;�u+N�q{��*��UI�#Õ�]Ĝ�6���9G�`��β�}�d'���T�k��?W�ѻ�@֫���R�.��NM��uT�dǔ�5:v���=�q,���OQ�dʁ�u�f�d�t��T�Ӧ{��t�>�h	�^�E���z�^�Zx�����.�F�=>��z�"�z14�7��'vT�½�-�G�^�i�)�����NK���3�/%Ը�8�z.�{/�@���"�;�=}�*q�o"L��	�/Ԫ�Y� �����zg��ܔ����;r[�����6�Z<��v�ڒ��@��{0��R��?�p$��͉�����B���$|	�8�������֌\Z�� ���~Z�zV��w�7|�5&z�Fve�a�$�a��t)�=��=���ass`�Nܪ��n2´ǲn֊�1�z�[� ����}�r}�s,�Έ���6G;&�t0�����g�a�	���}8X�!����w[�~fy�~P}�����z�#I�߇�-���33h{���u�疾n���^�Zضn�d�v�i]zXCw6s\���T�H=�8�F ٳ��a%P�$���z	)�9�~�A	P 2�ܖپ��]��W�������� (�Z�'wiá���8a�®�����.V��vd�r�\�٣��o.=�Xv[��/��i�sj�v�WD�lz���!YA�Sci����l73W�ߗ��˒y����6���r76�λ���_s�r���\MyOt0#���Wvy�ш��wusr�D��d�zh�UI^1�:D�K��Qj����	�)U-��B�<;�"5�2�5� �����떜���`m�qp�������!�����q̴jZ�/��,(r��UM�Ӣ����%��&�a������&��p=�~DN��5O�i�M�A��V�u��Bv�\�˃�0�F2�9�n�h����2u�Ӈl2����|�2u,�~+[������)�w_�k�6B�=��[���E3�6Q����":�u����;}�!��jKE��@�p��6�N�P��)䘺3������)�n������Ͷ-�{�C��M˄E�K��n"f� ���':�+�yx!��1�8�)V�.\˫&:h^�' V�VrR3c�9k�ͯ+yv:D�HLy/
,�9+���8���
�����WK�����au�D���_�O�Wƶ�M���z��Yc��"^�m���\\��E.��JT��!x/98y>��M��˵@����B���-���9��$g.�3����gVsħ�F��E-�<��t+�,������.r-�V�Ԕ���8خ���ļ|�Pݜ8C�\>�X�*�h��o*�Ɖ[�C���[��=�|�]V���v����V�jcޑ��6*(�Z4���K�J�~���M��u��U�oĒ	?}4&r���p����k��T��k	�2m7�&����J��?tL+ޙ�7^K[N�\�:-��ļΊB"5i��wiZN��m�9u9K�v�߀�-���11Q�[�'1��ɲw��_����Ȫ)yf��Y瑩ʹ�T�M��z�D9d'������K�z�#�qVsIH11���$~܅��?}dk����A��YOjBf�c�*�ʖ�j�n��h��p����T>��+^Ū�fn�߉�}R[���*�94�C-� ��̫c}�(�W.��Eb��'�.��,N�]�މ<�`����.���'��B��6��~.�z �Ƒwr��A�WDc:#�i�k�W����U���V�3oN�7,�:`3숄��˔��
 ��>�C�k[��o���m����JfLص"���fl`�u�]�2оeJ����_CN& �`��X®���Z�gx
�cȎ�+��vv��
'���9Vf�D� ˹�R���z�;�2�c�2�<��Z��j�
\yϬz�^eچ��*ڪ�hvGcHҌy���uv�CA<%�?���� ob4jehœOz���֣�F�k��aP�#t9y��񑧫ն:z?�����ӳ}��ߔAy9p�i� ^Z�=�۷^H)���]д�e�5���*�h6H9�}�s��k�Z�w�'�c�������g�9Y�'�V�k�tz*A�H�=����׽n�O�v�F�k�9,VXK1�ܺ4�pV�K���~_W�pa{27L�\zV�=�Uq�����(1����$��5�pF�ϛ���g����_>�S�����/��烗y�<4��5��W��*���Dt*�ه�.��q�YtДƁ����ކ� �Ӝ�ҜZ����9��Z踡v8n���+#�;jq���
���/��r�j�7w�k��O[���y��>4`�crfQ˖�$�&0��_l��~�w33G��}������ú��
�ڜ�5�uf}�T�]�Q��fν٪:s����t+�(��E�u8��5`����P�̻�Xyqn=O�#���G������!���0��Z��~�xi���o���u��
�2)LF�}3�8L�=z��ڵ�6��w�u"��Z�7���E�n�d���m�D|2����^Z#Ϻ�gp��$h���w�k�g&���.�[&9e��k�;E<krGg��I���
ت���H�{�iYG��4��~<=�7�
iK��̴u	�B��dr#�,Q!U��Mf[���y��xޗ ���o�d�^�c������]:�{ճ6���3;���=9}ͯ��قM]�	��̰{l��p�tyU%X�u[X��S���z��f��ŵٳo�bF�x}������dg��]wqv��FEC��%�d�0���6�ILc_#ѧH��s5^��=�̮Տ����ݵ���)������S? G�,7fcш���d�m�S�i�����@�6�0�&�g�i�4+�ae�E����R��-��	b2�Wj�l+��Ўe��Wej�����/jլrrު�ÂUKZ$o�<��>��2��a8Z-Khe]Q�l�ZQ�O*���{r/� ˹�'r�`0�%�4{5������n:�ƥȢh����X��ܠ*WP��I��w�Tr}T��6��م�h8(Z���Z:kj��3[X��*�H���6^��ݩ����j��'Q}���7օ3
!`$������E	�eX�d�W��}�h-k��b�+�X$�D�������/Z�Qb���o��ז��A��ʱ7�
��p��=s�O+Ȱaq⩁]�ml�h9�p�+1���(���t++���@�TM�;ٔ 1��08oki��D�9��2�����.�
�k ��4N�>�Q9J�c˚a���<������h�-�-�/;��c;�:w��{R'��͝._�~�לּh��_#�g�8���rxn3v�;�5Q0�_abZz��T�vf��9�`��j�^����lV������ћ��{ǔ���s)�+�u��K����N�jw���3��z���*�N'{ VWm�^��A�Ւ���GqT�s�\α�s���c�����_,.�)���C��i������)&gp\����F�t�w7l�����z����d]:N~���G��y�!��s��t��㍲Z]�A<���Z����]�*�x�N��^] Iœ��<գ��ۻL�kM��/�V�o�W�U��s/�b3�����4���r�R�]�f�������ky��R�X�m��rß�>�S���p)��+��,w�P՜_\��ј+j���Wlz������m��M���MS�33X����nDjZ�)���U����m�
�m�	��x����&;��5�ugi<'t����������{������x���5:m@��C�e��%�SE�x�X ZY=��wv;�&t��2oc2X��h������M��
����s++h�\�R���X9Zt�5�N�f����ڐ����1Uٕ#+	J��k�O��L �+5�l��Ҝ�Sga�������X�x't΃����ʖ��.�U8;�	���8n�,ί�wJ��zK� �]��Z��������c.��V�NP;˙�
u����A�ڻl{�q�on�F�$�L��R�4-��w8�fZy}6*a����ʜ��dǙ�y}GL6%�H�3vv����쒛������C��Ԣ��� >4�p.�v��H�������=_:�\�su�X�%�0�HW��Sw����XN��W(qY�l�*�^}S���{c������˼�Q�ܦ	,^��*��_pT��#皹g2�
�lT��/�f�\����xy��1&�6�LK;�E�A�k�����]WK��[���`�'uS��ggW
t]<5�Z�=u�Xl���
��r);5��B	5�tŴg\��1��dd��]��\��}^u'VWxe�����}���}�kY�m=�z}
�I�� u�h~�䗄�(���x�v�ͪo1�,w��V"#�*fT����+՝<����R��@���G�=Ƴ].��/�w�]2�����S��g,,gtE�'�W��v��s�x\���q�'}>sĔ��y˾���sJ��N����s��^�o�?wǺeM`�����.��'0��VWֻ�����]�z����9��r��LOܦ^���y	�������pi�M�,D�u �k�6Wf=zd�:�bæ�
���D;j����"���5;�ʨ�Q�!�޺ԅy`�?i�u��M��8�r�ڂ3�w�w�������l\G�6d�|q�\��k�ʖ^K����v���^�%����r��OUC�(f���tT��Lz��>V������9�޸tBQ���Y$v�T���rQ����9O�Σ�N�|v���1�$f��dj3WM��3,�V��e��Ӻu��Jm��w6�t�1��Wk��8h>�}sjp��l_�)q�c/ϗ�h���\=�Ē~�]����"�Qr�/o�l��%ۧ�s[=�^VNSD��pm���K~l}O�݌Dخs:�Ņ{����՚��-��.�g@a�^����̟��z"�U0��0}�N�\@Fv߉׷G��ԅV�����*��������WИq���xrǸ����5�
�C�\��x�Y�e��m]HWRh7�]�Ԏ*o��Y�{5��"��E�r����5v����a���|k�߾��<.�.��d�x;�>hf�Iy�3򹯝����]�7Ck%�3R4�\�!Y%�6���]g1��"$0����x��q�����u�wra���SMQ���Y�!�$���'�}������yU���vb���q ����1����4������7�l]1�%Y�=�J��hg�Y�g�`�UW.Vi3sZ��hk&�^�1̳B�~�ٷÐV�YheQ�LuWHJ\��L��m��t�Y�ՙݮ�w3L��ã�w.��2�E�̄�+�Ը�̀vG�(�oWv�w3�����8s��Q5o�C�y�A���A=l��;�������|�����S�2��ݪ���J`�Z��U�Lm0�4Fk'�e����sO�_�4��zN�y���� p_��ay�.j���t��y�q�I��`�B-Ol�	��
�U��.9qY�x�
\?}�Vt˒����J���}��2!%�j��<��Iڝ~��.�G_��a���xDP��[���(�e���s��t[���_>�U�6��}���_����׎�΁���{<lߣ~#��ǎ�1u�	^��8š���ૄahr�<���u������FƊ����{�_p͝��̌��S3N�a�{�#��vP���S��'Ol�l��;&d=A;&�y�9w�p}a�E֦�u��MQ-=�M���UL=Ͼ~�o�o�E�2ް܊��⼣i�ǿ~��������}�V)��[iO��>�Y-������N�I���w˙�8)�9];P��;�@�����;��sy1)��mA�w�3Rj����&�.�b��'fZF�<9�x�m��)ͽ� �29O��E�#����z��ۭ&������5���.H���ò
z3�����V�V;����ѕ��C�.$;1&	�� 1V �6��q+=>��G�"%V�ĭ��,���]ԹˎG��Cx{���sJr�<#�
[����%o�g��ɾd�O*�ǭt�NP�����
�1J�<.��Ҍ��[.�,Q�tD���]6��(�UFX�誱�R���!���j8��my�K�>0=�$l}<�s�Y�W���ŉ��o_+.�f,�e���Ҫ��')f���-�N�u�ѭS�^�m������g��+>��!0Q��[�����V�w*�bW�࿸���/r}���������b��9N�w������J;�o~�s4��z�N��b�G<;���|�b�d���a^�4��e���9�{��n��(���}~�1SbTN{�M\C��
ə�kw5{����1	�@{&�̺�1ud�ȕVO�k�w�h�ȩ����f�ы�o���Q3��"嵷���[)�Eɽ��-�Cf�㇒9c���N�60�k����z%��3+ON��)L���.�se���V��v����	 ��9�+��M���I�����S.�uut([19�'��,޻�^�V��Z���vGyH]Pn1[g=E�Ѳ�*�i����:��%���)�|k6�ݵc��r/��xM�6�t�S�=������j�>��bO��%�c7��;ǈ��F{zD=����|~�7=���:�-�x�۲�m;�9PKo+:( �}uMP�<5fUp��M��	��hY�.�U������\hi��m�;j��n���wB��ʹJ�Z�Y/������u�"*l)Nr�D�g�2�\�����""�)߯Yva�d���v�4�+���;��#R�cn�bGgU ���t1@�yM��~E�ʧ�ϊw3u��kǔ�u��=m�i���@�z���b��)�6T���^��7ҽ0mr��x�1<-(��Mt�'r�Ӛ30I���?{�5�s��&���}ח�%]����<����9(��պ*��'pv����s9��#U�$����Ѹ��&��3m�L�/^r����V�������I������{jb[��X�{.�!DE*ɲ������g��ڜ���+<}wN���	~���8�񢞘��R��:g�3}g�o������{_�!���V���F]wl�L����0ya&�e����S��~e��24���;���@�H��[?�t��l���7�y~0����3Fow���O����C%�eN�g���)K����k � ��͙=w�cU3'ս��)6��TRg�cE0y���ȅrwE? O7T�s����8���<:7��.C����U�Y��^y�x���K�uN������ �4L��>���H�pr�����3��.��3����s$�7C aEƒs���.��<!B��ܺ�-o�EE�^�}��O@�fSVU��~lք{=)E�5���������R�wdRѰ��ۭ��^���}tJr� TC�O:}Y��Ǖ|��=ܑ�z�������Y����j���qX�vF�JA`N�1����.n�.W�8�/�t�~��a��ou���:�&v]
u�|�U�Pj�l���ؠ��6���Dj膽���4�EA�z��0a�N�am��n���d��t����bo�g�D��eS{�fWl�(�r6}�'�O���j�B��d�1���W��UTpE��O�&gmv^�G��vp,�	t��ϴm������_�R9�
	��o`i����*1a�} Zn��5�#b�����&�;zv�;�~��"8B����r>�Z��Z"�)7�М�@�5�v�ny�"-�Ld_���| {�$0ߩ���/Y�W���M�w�ӓv��>\��s=]����� ��r���zf��5ex<�:�������p����_���u辥���o�u]�I�\{�����;#f�?��BtT\>��W�l60���R�nͤ1����]��u�^�����۸�l�A $ &�j+���9vp�[o�_�\1��[��wS2^�Mb.��N�8��Md)_=�j�;�D�<�Z�y^����n��g��j���p����7hG�Ϋ�J����i���4Bi�{ �WX���u���jS��O�7&8g�Y�~��{	�����r��e�r`�#��Ves�n	)^^����n���2��s���Tvs|:{vM��E^p7�Hm��n,�e�yJ�����5N8ݛ��A��6���T���Ϧ���^5/��!h���=�7Z�GF<)oob1�n#R��[�Jlt�G�� �9u`T}�\c<t�kQ���;�u'oL�8�4 $oUD�c�/� �mZKpõ���@����fV�$>U�.p��SB�w�T�k�c�K*P��y��Y4�ֆ�h�-��-[]�A��V��JN�=9�ʜ�Za4�,i�uSJ��KG<��5^��풸qxˤ9:ӌ�t�V�>�G'"�B��W��v�>?Ff��Ѹ�V��d>�Wֲ�s��[5o�-�RWI�O}�}��Z��}���}�����JĈ��d
�G�7��:�:&�G��ak��8��w=H�ؚXC�R`ZT�����j

_B5�G3y��!���0��m�_�Q��_�:�93vZ{��K�c��{��֚��9pQ��غ�ݒ5����y��}�ޙSV}[��K6��_I |ZIb���'U�,�x`�c����9jmf��v�/o|C����ﰅ#އ�
�L��ł��tay���֭�n���x��&]ԜJe�ˠ��]P@cz��z,jN���oyExYǴu��9���z�}�
�5��[��]��(�!=�*j-8b��7�O�~z����V��ࠋ��D��ۇa��ׁ��a`��!�f<;0)�C[ǯN���E:��;(:N��Z_��θ4��r8��<f� qb;&�awS_m�S����Fd�Je��⮊]\��-.�� u��p��e�s񎾟+���]�V�C2��7p�[�=����Q���|�ٮ�|z��d��Cܗn�v�Td��F�l��=xɏ��������$���>�v���Pt��#���y���?-p�Y��z�;�����hf�en�E5r������6'}[����Y�-O�MfMoF�P_%�6F����yF�A��u�Z��ëkz�`\wt��ib�ՙ5kA��*qH�}�߬f�e�w\8;"3*��>
��T��\ �x+cm���=�}����,~��ȿ!;.�ϬD�{��g9J�ODrȽB��w�L�#��էu����������Ź�c��3Vr���tqU#2f�Mdcqn��j|�;iC��Kގ�m߮}��w��cjm�7�a�a�{�м�\wG�b�\A��>Sx�9~w��6+�=0��ȼ��j�i���=3pm�|&�cjw,y3쪔�����ޤ��~-� ��٩�ց/�b��'��a�+�b�%�DĿ)�7��ߓ5���~T���Z�^��-/~��ͅYo�x͐0_��5��s�g�]x�T���"���݇�8���*��q.��9
�]x���ܧ���e�;=��`Np�#�d����,�Q5��3��@	W�����m�%v+��Ջ�~�B�����q
pk�yx ���sLGwF�ۼ_��}��2'b��Vn��WX��NtW<n�1���s�%A��-ͼ}7;li��=�`ޠ�Z����9o/�6�JI�]�+]��!HͲ3��I9�� �k��!�U�R��΁=�k/WR�3�k��<��&_���O{>���]���t��wL�yW.�ʪWsh�8]�yٹw��9 }�4HeL�ϡFv���7�v5f�
Be��WG�Uݟ��-"WV��y�^E��X} b2��:ί�E����P�=�u����^�\׏}���|�w�@��&�d��a�}�6��$	P�}�3e�����6�>���ݳϕ����X���(dB:��u�PB.�RՊ"+1���
��i��k����T�d�\r�'P�q4C�D��UwN�k-�9��P��
�7"�'�������3l�����/7���Ԁ�������(F'���,��N彶�vo��N�8v�|D��a����5̦�L��:�"ϝ��^L��&Цc�5�`U�$�)��h�f���:���;5@�]4=$1���Y��c&�����ϊ�ػ�㻼c���I��GE�zQef}��X?|����@���Ԝd��P�s���gfb�͡/�x�7cnGö�2��Kh�$#>�_n�T������Q��IkY��<5������M���YzG���̭���:�fc�c+�!�%�sn�W�"�9\�T��P'(��:4��|KRmkw�l�N�Q�W��_VS�V�:���Ta�W���*���X�w������6�H�G}��vX���}H�����c�Z� �B�M��{���E���:傲
�{��]��60�;�@��d#�R{%v��zh���g
Pd�Q
����-�M34���$,Cr����]5֍�gT�oMvM�\n������B�s��[�n�c-I�ٰef\�\���NA�/@xE�&��[��v�u# �|�\�<�j���Z8a������n�mփܐ�['���;Ǜӫ���,���֔�b���Ɍ{��++���[�)�C4������zQ�D�[&ƾ=gLj�����ވu~[�0e�`%Ѽp.��wn�	�KW;�o���3��$��gj�:4�ܾ�=(w��[�mŪ>�2f��e�uF�U��I�mX���o�3�;�Wuq�ŧ9�E�z�n��&0�ۦ+�XKOP�u��4�)t.N��Mb����b��k<����
�83��*��m�Mʬ����Ή�q\��s���r�R!Vr!V��hM��]�#�J���_J*�"h��\[Q�2�oE�gpPƅb��pڗ���%('�V:��UB��E�pWYWf�@�*����h�ݺ�OF�ٗ@�[�׎��!w	G��m�e�
he�С�c���K�M�W-ۀ�w���.�]�ޣ3������s7x���N��f����WNә�2��(bfɽ_������ʿW���&4�T�U��Q]|�f�����i>|G]��]��]�)�M��o3��^�2�GfF*J8٬ӈU���v�˒�2WjQ�ٱ�>�ٞ`dU�|kx�[SO�ꖳ�A<���+�ni���ͱmʛ9#%�S�С�Ͳ�10�3#���k�����C����G����'�`_����[��z���2u�ymGVE��ޱ�y�rԯ��+�:�]���Obf�
�U�g��]*�j�a��=�����&b,F�vt%������yC[��W\���:�=,pa��.f'iU�@��a<sgޔ�o���p����s"nfӎ��Y=��H+���[�{|�f\Ae=�5������� ^?z���*��4iϏE'��R�8u]7i>�ey��;����If���+m���nw|��[�d���1e+��,it��v��gY���Fa_�\o^�u�QWa�+��d�V:�m�]lEz<�_�u�.�x� {�DF<iΉ�u�K��F�i���z�B���J���U�[}�Ɖ�.���?\y]����X�����X3gqF��������Ҋt�%5kB��Xz�\Fh�y|"�J�>(_������=S몹-,(p�4��{n���F�h�V�6��74��<b�Z�9����wX(�.�nh�s��y9r��cXqx��}�^/��	���]�Osj�Y0jᣭۇ������MՉ���#��mш�'�79_�r_������Ót�K��J"A�ޣ�p{Е�p�F�����9�t1qck�䇙�φƋu�2-mM֌"l�����3�������_������ ��+����[�����+���o�Y�J�y�����X������o�\��A��B��M�{�'�hv�o��/�-V]W�o)��Ҧ�)�/�����vuz���e�<:�*^n�+O/X��0�>�+%��51*��^�%`&�.�94�+p�)�{��[5C3#'*�l���y��zl%+��]�=��9tx=O�V^�g���3�5}Yi+Ӛyw��N"�� _fL�3!��h#/ɝ9.br��E|���J�a�ͻ��QTXț�c(�ʻ��V��[7�gR��Q�p��E�bvp�:�nG�qYaН�ci=��*Th�E5ܧc�;�خ�����x��z�ϴظ�*�pvhi{1W)'��ml�]3�%���/j�������sެ`��m�z&2Z��<�7p�?}�>�����ʫ�h��Cm�%�Cj���GH��z앐�ǱӃ�
��j��hjHjm�9�<c'+@7_�)���W�/���u���H_�16T�z|�'tʋc��w��ە�
N��`�y�S����ܠ�z�:��x>4u�!�bx�\��]����5Ri�_�cO=it�8)}�]���O[Ϝ�{(���`'Zi�����Vwu�D�5�_rּ>�#������K:t��m�H}�D��(����9�U97����{i�n�{���nM+@Q���<���\0On�CF�o�ӗ�OOg�Z*0[X)��JױͣW�Oz���hj�KNA�uno@��ySl���> i����C.��\�YY���o�B��8�Yi�ky��8̜�ʾ�Ga��.q[�l�N��'+{o��L#��#:�S� ��%(��	%��y�xye�boCܟm4�*�;'1��A���}�q��ꞽ�.ŧ���=��B
��-f�1��p1�%�m[����w�oL��Wz�I{���.�F;�C����i��[f�p�BEm����@a��lg��洪���\R�YG�rR�pF��j����g�+���4����������{S�=�Qj��
~�w3��DZ�[��X8�o����V�F��ȋT���ꛫ��^�1�6�qe���[��F.6�վva���/��&6K��%�l�nn∹��f�Ԧ�$�˨L�;n�XP�r��Y�o��&�))|���C�
�[�s4��b�tI�;� }��n�[�T�;�����]�U/.:�w�ڻ�d�S�j2hTzj,t�]چO�Гd����q
U��3���ǙP���L ~�=�מJ�F��b���r�h��������FI��eL)!RX2=�w��ϳ����\wv��_^o���]d8��]['>��77�ov4d����#lVi���u.����n[MYo;v��ړ�VT��v��m����l��~����R��*?{�A�f��]A�wo�Xg�r��W	�e������}4`���Zr5��^��w�S�!���:@vɳ�Ω�3�=0y��MNCu����wD�	���-LTZq��w|i��*��A���^�=#��㧆�u];t�8����##�>�W����7���v�S.���l����~�:�h[V��U�uUUH�]��;��[�Yq�}�>��$���C�!p[�g��A�����3!�:A4lɃ�V�u�/M�������֏���N>~S���}�̘�.��>�0��;Q�zw��8ҍ��=�yEObO�rϖV���fn�݊q͜s���/P��!��q���=�7������ܨ�n�s3��4�D��Qou�]�mkS<�*���	�82�|֊뷸N˘����ƥ\��˷F�;�[2�@$Њ�tyB��@S�{[[��7Ѓ\�Y�ƴ��u��>/cu�m��n4�2���}��F1�X�o����DЬl��t4�a���yֲ�pr�3$�G��>G�n��ѹ��f�"3+\Ac�?��.G�:8ཥ�s�W�@��i��W�;E�����5�~�����r�)�T�m���-d�q5���f|���j��Ll&���o7���5־֫1���!���W���?�3�x�Ҙ�%4��^9���1����[���Ԯ���1|���e
p^�|+��myv����aܜ[�����[>�Q9�4�:�8[r��F�s���ǿ=�6.���2V��Eȭ���Q7���ۤ�TW��|֜���~�{�}76:�z��R*0��ж����>�zZO�iS���f������싹ia���u���LaC�Cv`���V�[�1<�j�Ynogk[9}��L�ĊV�:��ʠp�2�'�L2���!�Jd��pfo5��ܶ}��߽���f���r�ך�E�\޹�rԮ��5�o8cA.�dTH�}��:�F�U!`�DL�WAl.���73>�W���N��F�E���I �d����Ŋ���7z���]R�UK�����g?d�\�L�e�#�s�i���8��f%.<�$b��������W�sw1+Ѧ��la��Yg���9���z��#�+{\l#�r����ppV�eL���v�E��Y~q� ��嬊���N�L�̥�\��1���n��VgU�OF\jͦ��rC��mԯx3]I�Q�}a�F�&�ƴؔ�&M�&�������c���?�[fp�}�.���FU -��^��:����t��~38̄���.�����;�WW�|'��>���k�����צ8��*��]$ח�<�dNkgK����J���7�!]�v�1�B7���=��Ն�E��_��1~e��sH�[~7����8B��'>�x=ؔ��Y�s
�'�9� ��C�e�J���t����97!`���Vy����['�'t�۠C�7S��6�G-�R�αԧ�d�xT�,�v�Ic27jX�'�C��/�� �d(���QKke�􏸷�Y{UK���.��b�]߬�'�/67y+�[�rԒ�r���sDFo�C`�L��T���vd�u� ��M�5�+2|.��%{�RLLռ�q�;�� 
щ��8������}���?W�5_j?�%Z���e�7�0W��<�׬�������_  ��}�2tz��uJO���eN^8�G.z�V3Z�27�������ΉT���WW.�k6��y�3��w��ԯ-9�2O�� ����!��$�Ym��ޖ���7�$�MUE����m��s$y�ߵ��5�~V�`��3rZ-��~ �D�`��W�Męm��ރ��J�C �%T�]��zl�Ǽ��ź@�۷�|oI�.|	-�)?xc�$�W2��vD.������V�Z�s^��TVT;Bk�u5���c�y�J��Q�{�w�vXXcQ86�e�\�h,jA�����e�N��Ò�\���]:Oq���G=ԞK�[D
��2�s��d᣶��s�.�e��!��)5�i�%�4e�Q��4ǧZ�N�&fu�w���ݴ�x0Y�֍dz�vU��^%u܈��SÌX�{��K�v�|�7n��bK�{6�M��`�<S�ة��M9����V���C,��u	֕�z��pQeeGԴ�Fk'm��=�� ��� Q5[����v}g��u�'�7�dZ�0�܉���E٭����wA1�\��eb�d�jD=kf���}�T���r���[��U�Ȩ���b��]}�W͇��w2�0�Ճ�u�f�o �˥{Ufd��V!���<���Ia����&��~�cF���[7~���'A�V*ڼ���/ :Z�!ϵm,���aV��UD.\�}ܪ��/#D���������m�d_��� �}l��ܳC��~6.7Wy�q�Al��2$_��8�a���W=�mj6"�Y6��ٝ���m�n����P��jD���ul_;�:E���w�oҚb_�u�˙�=����I�O!̻T!P�T(�v��V�r��W�]��H��U�AW�M����z�˵�Ѧe��0���qWt�}�]_�&HM���*����EM/c���#:(�΢��F�2p�.�f2K���׼t�����A+B9��Q��9�.y|8mg9Ukoip��]a ����
&�J�Y���sl�yݮ�&_�W�3zFD����۠V�nn��#R�l��ċ�zG�i���z9�^��{�y����O���l�3V�P��ݨ`s��;2�Y���T�����]��\U\E��~���*]�����̈�M�]�C� >S���X�/*0/L���[ܩ��M���&9VӢ�$��Ò���e��ٸbwS�آ���6& �L=w�Զk<���=Ăb�Ld��sO��xN�����~�l?t=~b˚����.�O��$*�g|ιlY�?��Q���,���{�'%��ͯ�qp[b��h*ed��n!v�+�V�w���77��d��M}��Y}^��=T�xJzz�n|I%aW&�(�j�����:܅�5cxz�l��z�P�^}����,� �����
�^^<*ͷ�ug�V(7e��BVM���%�6^t�2�E:�2�x��ܧJ��+�\�^M�����[�lc�A^�t�c��)QE��s1�֥�I�����X�[w0�J��ᗕ�k��2��[�"N��Z�9U�:��5o`�2rjέ��xA�_�OE��I��w���9�i7�^���'�Ρ����������W\�%q���gVT��)�Ӵ�A�vm�[X�r(X|X�F�=b��n!C����z�r���H|�J�1�}���e�$�߻b�ʬidYDgZ�����3.��P�xQ�(@�6��I� R@� i �H(B
m���������9~yǽ�k~�kNal�S�Ɨ���P� &��C���S�>��et<�FM.�(�����Fr�Ŕ�E���7������R�lrv�,OݗaNTsÝ]��$�'K�gt�cYm��
֝�Ø(����i��HaHS���8˗��[�z����{f��`Vq6����uYY�cRV�-�k�CY��iS·����gx]�����`�!��6�%���0�	�(R0f'��.�e���������~;S���쾹�}����z� i$�;v ��.B�qli�������W z��K�\�H���%LK�Mȳ5,'>��Z��iq���eI}�eҭս�8B�;t0�;&���l3f�lN�Z~�ᙐu��
��Hm�����5�Y$B�$7a��E<듥Eq�]�y�8ŗ�FhY��\�f�V\ŶQ�J���ܨ7���t��rI;�Io���-T���孢��;��w�{T�I�3���2��Hr'�æZ�GE�c�:�i����O
��5uf,�y�j�Z�X��s�Ls:%qڇ���&���![Ɩp챜�rv�n@���u��'{n�Wma
�ԬN�<+*D�)�"£K��]�}�vX��u�틏u@�n��l�d�[v�9�loEg4yx��FP���Q���N-]��\(�u���on��l�X:��e|�E�ф�G�.�.��-d}�9f67O:6S�w�/S�Պ����̊%˸���7���P�e�B����0*�6��<��4ɣsQ뷝����ЫS�ۺ񫶸��]��x�̀�(O�f<�[��U)`F(��w5W��͌�/�����~GC��Ұߜ�W�:T���8�@��9u�.�]]�ȗ]I��L�D���bA�i�P��96^s]7n�7��a��w���D���\ڵ���Y��f�)K��zz'}�E�H��|ɓw+	����KN��*�P��4*�*Go�0��⩼�Fw.��(`�����N�ӳ���NnآqD�Ӝ�u�CEǤ��f��􀍴��W�J�t�v
��ta{4U���*���eN-��p4ˠ؛S�Eiqm�I�9�����[Q���Q@����:fܹ������h"���b�\A�뫻��a�:!:�o�/ �"�K�ˊ�(���o ����9��R�XTew�qF�*S�|:��o1Sӝ�����Ÿ�Ie�2�d��;P�5�S@�7{����ѻݙ��C�̓"���Ԑ{��_��
��j�K�ܻ����_�����#A����m�N2��㡛X�SrFK�˪�s�\��������&W�����@I�UV���q�w���T��ܢ(Pg�����|�sQ�����c|hF�SXr���|^̾����h�o�iv������1wS��G%�¬�Yvۑ��VS�+|�!����6�m�v���lmvȫ����3<�x.	�W�VӐ�_|�s+������v"c����B6o��4���Ϗ���Wƫ�kh}�!��Z��纡�e���F�|��T8�lջ�QO\;//٘�D�kuϬ�z~'����ey���q�2�~=@�C~ħ$R�R�YvrM�3Ň�* �I�/;g��j�߅{��S�in�i�}��W�fV�'���I�ԃB���{�?����?�s<�u��^ip,,���3c��ߥ]
�r�$�[`\�Gsݣ{J"��U�.�z���pYqMl�vz�r��2P�\:r�O2��ݫW,��sou;<�|WgK���$h��IL�K�9ذ��^{w]R|կ��G0T�L�՝b��U6R���:^FI�%��{������c���h	٣���M�'�m�{����>~w3��[~d[�}v�OgAݻ���3��s���_!��߅ʁ&|��D��+��mv}�[���	��mOj0�xH�22�1=�qXnK�h�l�6[��m�x���l��n��iE����Aa�k{���5uĴ79�d157�Y�׺ޱÅ�e9���\.�,6����Ϡ:�I���k�L�<<-�xnܤδ4ni�Ĺ�]�Naŷs�r��P��d�W~�WU��j`�+e<�SM2/z�͖^!xKn%�q��|~�d��	��}}Z'���V��2��̄6��VBVG�c*��gߵq�rH�ǫ������i�Z��ϫ/����[h�O��܄���f.�_�ֹ�w�7�}� �@^�0��Yj)-b��TYEc.(½�ʺ�{�(��n7[sP�y5���3����ISl�gu��H�ا.7��Ʋ����W�����M�Zwyh�� ��WR�b���]J�pԺx����&��&�n�H�\X� u-���ǥvb߯7�ܠ���tTк��c�����`+�NA/�c(N]��p�ҫ}�њ�b��~y�g�_r��f��#en�v���00 ����7$|1����d�Fu�r�Zhj1�"��h�1���Tڥ�eTu3AFD�*���NPݯy1¶5�1� �op�㞼�9[;D�o(�DU���y%9�?�����x|�c�&dzNג~�_M�U1�5\����Ì��׺�����+�����z�|���+͹6��^� %V�s��d�"W��:sN�c������޴�]�ݗ~鮏Kt�i��,浝�W�@�V�~["SҾ�i�,��t X����x��!�� d|��=;�}*�8�ܩ�����-��5�[���I;�����ءr�ȯ@��Mc)�	�y��@�׮j�T2 ��z�v�6�5.����r��p>}���E�E�v�3vbߴX��5�S�܃&�zk�D���B�h��<�[�&�N���b�U�-b X�1/'=��('B��,^��^D׵����E��%4\sP7���/=�	�TTՙ��[ܦ��j�"ǻ~�U��ͣ�g��T��_�{\=���9/���X�����݃d�Cy��̏*jI�d�i�]J�+�~��3� ��ۮ��oD|��N����"�����/D�J���yC�A@b|og�������{�T��UC�%�?f�j����}c@4H՗�^�^��4��^���Foe��ϻzU���g���"�2�=r�ؗ��Fn5mL$���1����>���tx��J�;H��\�1�={�Ł�� ������O'w��:��T��6��60�e�YX����/�ެ1*ao����cw��wX��)t:d�l�E��)��D����?|>}��K"OGv�0��-\��0sU�E߷���񕶞ǜ��o���_"L�]}��q��u,�)��[��]�G#x�42l�DA(�W����Ro�3eG ��������0��W1x�]*y��G����%��>�rNE���Y�v�m���u}o�T�iҸ����Dʳ���7�?J �ƿv�G.[އ�7c�� ����S�N4]�f;��Y�{8�_��x1�~4�Ê2+a��*7�kf'����5�y}��g�~�ՙȭY5K�r���0���~�Cgե�0[��ԑ=v�
�Q�����o�+6��>�i���-s���v����N��j�L7`:�'__�C��^�b��H�>_V�p�p��/���ǟ�ض^��h���a� �?��Kꝍ����wp�� <� ���k(�J�䵂&�Κ45V��mǷr��wVu�-ieO/r��nU��{��d���ڧ+@ ��R�B��nX�G�wC~�gr��|�r��`�����X�o�|_gRg�^/��8�25a�?���W<�,�M��Lη�mF���{_u��9Je�,-����jر
�Q�)E������Ƶ����y1��>̋j�4Z�I=��)q7
�*�o��/wrt·��D�f�5H(��}��J8� �4�];�ʏ/�ӭ(ՙ����{��믿f$����Xk�J��!�˧�V���dF�&�]JO��n���DmW��|2�/�j�勜��yN�5~ _�}�zmNf�A��̞�O^���ET��0�s��MFa���A}��t{���*f�ģ���d
��/[�fOW��)�-���uI���[�� Y����V,�ʃ���|��hd��V���B��m�ú�K#�ʍ#3e��f�N�0F�x>o�:��N1��kJ�}e0"��|�mg�Y��^j�mc3e��:�xǥ÷H��� �'9UxKj�ɮ�p?G��>��{��ܞգ��g|�1��%�o��]ߨWLi��sr{/�Z
�{.Eɭ�I�x�Fց;^�}C��e���s)�E�˒�e^*2~W\�}� ��ۚ{�>�y�I�������;���5~����uU&��)lCs{������=����� �]����'JK;yp��7�ݡ6Wq{I��ayӪ��w���o��S��wc.a;���/o���׆f��|��3��m��x�>�gbW�/s!vi���U�_���G"sg��y ����ֵ̈r �g��ɟa�ݟ���뻍����z�|�\����F����kx�/6���G��([�����"��h����r����X*�-R�0\��ٚ
�/fSE�Rʊ��]�+F����ה�n�k�4��.Y���u��|~$�������
]O���n��2r���tf&��O����_PN�#ۋ�[����Ć� ��.���S=�Q��~�F��Li�tsk��E�w����4��	���A�}�7����+��J[]2V�C{܂eN�Pf3zM��|
b�<�Vm��V���կ���<1t\����q�T��;Vd�Z��u��M؎��#��X���'�r��잋n���ʦ���ً�$̇z.������|[�R�SVSQ�(L�4�\�D!@�
�[V��8�ū��Bmf�pLu����g��7K�n��J�/2�S�
�c������R�ޗLN���Ӱi�֨2�w!�_D����'�;�gM�n�G:��<,H��\��8��߭?e��Mb�L�-�D	�}x�H�,�W1�{w+��U�dX�댔&tХ9�s�y�=77�CX�������V%�̕y^F^��dX$�!�����v�{.�qڪ_�������-���S���w:�H����M4z����&M7�9>lC���8���,f�%�Q��J�"�O1�A����[:�U���N� 8O��ٱGl ��櫉&Y��}� �a��L81��R�_����A���^�2�;���5G
��c��āM�W����a��i���2�ğ�N}����,��o���,��o�����.���^?Ea=X}C�ٻ*���;dQ����ѥ7�Q���(��~��9�F'�!����wl0n,b��sw{F��ͮ�%V�B���f.kkՎ3���S��hu��}�̷S�.�_t��ǬOt���͎�mf�C:<e��*)M%є.���$�TN]-B�s���걽Y���:����q�j͖@�U��J��t�0�w?Φ���l�ꎭڭE�g�Jb�扵��Gr��}�F˼p�/��ku�Y�l�����oo���>�xդ��c���j�i��ޣ�#ķPb�m�J{��=9�=X��Jn�|��߀>sW+f����O{�.��i��!EN�n���ZwAm�=z'�bzݢ����^���j0���!�K_������c�
92>���;I��@P<�2��%���\�kV��vJ������꬈�W�\ms�#ܠ/ȧ��^-��]�pU�3/T�Bf�{��u�Y;Yt���z��:oRVz�ޚ+&s	b�슝�)i���o�,��[��DM�Q:ӭ�,Y�În�"�C*�*��4_����0���Fsu?q�ʟ �	7F�F��̪56N�T�#f�3)�P!wF[S��v��O�_dfޯ�|���U؋gi!l��l\��;��E���ܘ�����V6����kED��\���"N	�ҡ[��np��bd`���OD'u�x����#��:��;CS˚]�s�v\�1�(��0�Ʈ������b.��[�*��A�Ɵ����虽bT��[�Vb��ǰ�K���/��J-�(r�~����O֟�;é�aٸ`G��x<bŇ��ꤤ͛�@��y��ıl�ve��ݱ���F��E
�خ�!�MD
�B��c��!w�`ݝ��i��#*_����xy��M��"ܭ돾���������3�G5x���zi2/;�R�~��wH+N`o������:���+Z��[���n8{ �v�D�p@�k�ԓvt��U<�]��쪡2J�5񼦑�%���`ٷ{+����< %f�NJ��DG�`��O���p�ڱt(���[V�cs��w��RYwN�NY�5�8�c<oa>�[UI`q߻fl�@X%1���7�d����V0��*:��A�mm�s��R'��%��e]�.�NP����R����X:-�U��	�\>~7��;�BFhi\�bI�he����}�F��$厭����19�gv�t;����݆��b�ﻦe������kfd�+^i:�3G]�yWɑ��9���� ���-j�n�
a�'��[���uҗiM��������zls�Y�E�/~y�����r�Às{ė�\]��.��ܲ��k�n-L�)�GX���YǙ��g0�;���ܻC4�W.�hQ%�vԝ+��3s�{�~�Ю�	����3��/��޹����'n<��w�������X{Y)`s��3�bUog-mX����{��6h�r�Mi��5��N�k	΂8�rt6�sN�F�(�5W�qn�!]�j�'EHL$'P� !�� A{#7mqn8�M9��������y��2E�Ҁ��+l��+<�	o-
.�'��5sA�}�].ۻ���#Y�����El���F�|��i�d���p��VV�(���ŗVp�4i���c\O����+��s冷�̅�沺�n��h�˧����A�9:�lPKD͏ְ���.�pĪ6�Vv�X@��4Wn䶷1�j΁�W	��,CF�W�4�?��G���v)�m�)s��(�^���������-*\�Fռ&�<�KZzTh&�,[��{�� �eܨ'n�[/����2���Vr捅�wqޞ��,�2U�,�f��N�Ӭ�S�'!:����9��Q&.pƣ����kG!�s��B̕{Br?Q��ݓ��3�h�jњ�+�����'t��m�ےee���{SH�/t�L<!޲Oe�]er,[n57��j�G��c	�"ꠞ�Ŗ�\Û
~{�әE�}�r���Q�2Tʌgr�c)uw�8��0S㏮��Ӫ���8��Su�y2͒qI�#A|��ˈP��z3(��F<��
ctvr'�C�q�'�KU�Y�FZ��׍R�R6�&�ə�/s���k�F�E1�5Z�u�{����X\|�p�_F�k���"�hW�QMڅ�}O��@����	a;��D͡It�/ql�����37����:+�7��5¸�ve6�#gn�os�a�j�O.�u�]j59p^h�X�yv���J��B�{v�e��U�d��W}�6V:K99AV�
Z'e=��:�w�od��:]S����N�&�4��qw	{א.���V͋ݞJn��+�� f���vu�S������I�y6Tk!�2��gݹuj�d�\Ar[@^u5Tۛ����K�!e��X�!\������+J�Ƹ��y�c�5w�D���L��֩��D�ԭ�����N��?��X�FbU�1qY6��y�ٴ�t�k�S-2a�f�e�ŕ���ڰ��ml;w�.�Ñs�Q�jlnp��S/�ݳM�~s�gN2���N�t�l�dN����bi�HK�����䵶낸Ͷ�t������w���aY�f��*Ԛ!Ѧ�&匚c����P�KP�z����qU�0G���&�	�[6j��PS��n!� 2���)�N���olJ��u�E�^q�拼�Ք���~h���Q�|l�qc�+_�/o}�b����j�G��9����m����? GU��
��'25hk��c��&�U�8�`c�,n�Hٕu�.̬t�ԆtJh�i���(L.!)z���(xx\�tl�=��C�|��iV�oIGxQ����uk�zL�r�B�_����gJ
�ᯗ����T�=p&�xsW������W�oX�^���d�G�6��>� YȿQ��g���8Ϋ]���&��G\�wj�MA��.}���&0��XS<�l�]Tc%�@���k��t�E�X'z�p�^�������.ws+��ni�:���d��LL6��d���᭑�Hc�1�L�.gv�9KTV^f\()���-#S)Mm"�XA���5uc!�Rs�s߷�����J���4��y�����9�w��/?t*����=�e�5�;?>��ʐ��k(�s�lvye�w;�3qD����#�*G��%�:˵S8�q'�*�ԝ	�eK��=���^,� p$��Y�����^
��3|1\������zLS��[4N�R�,����gRi0� x��ΎM��(��bO��k.{�p���^4�]y
�\�廉���]緻��r��v;s�ךq�7圼g��/�e�}��z��ߪ]~�'?v�0��_�~������>�>0X�5�R����p����bZqd��I~X�%���ꫪ����w�9M��=���� �A���? ��������L�ݜ��6��m;��@tLz�G�]�A���2mS�b~�}<�/E�]��Df��|�<.� ͽ,����;/8K9����/������صY���ʾ��Ʀ)����pUR���&  �Oj��F�C�Շx��B՞��E|��6E�ׇ+�Vu�ygv��"\����/��T}�}✤R�S�Z8Ԭ+$#�`�`�P6���˭sZݼ���;��f�#f��g�.\R�v]@{��y;��Uu1-����d�D<4c.ASe�{uό�yV�s/251�rv���/F<�wZ9�w@T��4�VX��)���g7�F��k�3�-���2�Ļ4�v��S�v���6��)y���m]b�j�e����p��T�󱕻�+휷���.�Y���^aJ��ek�{�]�
��C(�����fv�=�I	M��Yi�5`y[�kkyL?Gm]�#zb�%�ۗnڀ�w�؂ϱ����]�W�F����O6�+�6��J��Ʀ�䩲�����oK���=>]W�N��2�[�� 9�74Cd�4�0S5w,Z��¬t�=�R��&q���z�כ��3R���z��BT�.g�͎,��zw�&P���T��pj��Y)u��f�̯ X\ͽ���QIe#A�>����,�7����Dx�٣�%=�뱑�9�C�������Q�*5^��U�����ą�{M@���U5C:��^ύ�x`ׇ�ho��o���SJ��{����r�,��f@b���o+����C��R��C�p�&:�s=�1��"�_K9���n�kC��@�%Բ��ȭʤ�Unh&l�LH�R�9�K��8{Ef�)/�bn��5	W��0M��T҄Ѱ#^����c�Ū3�vRzݸ������{[�E�v7k�3�]�
�`-���F���M�2����x�IՃ`?%u�coJ��̠�F��*���/���Ό�՚Z���[G1���kL�=r߫�<3f}�\<�J�du�hH�N'u.����������잱<�Pe��I���+��c�WOmI�����B�>J�%�z�{7{�}Z�-��P�~�=w�9�+,�D�d�A��=q�m��HT
|�3�ԛu��D(�a�lEȵ�
ec���C�ೱ/'�DL\(���i��C���M��p�e�s�M���{��Rj�,+���g��[oW��\ס-@f*��a�݊��7���v.�e�d�9/cp�t�
�����\��]m��zk7�ɦ��X/nZ�Kۆ
&b5Dq�(��s����ok]��V�-�����Y�V���*�s�v���+5����uwF�Ж����˩*���˜�qb���y�ݘ �VG`2�v0�(�_o`3t+ݬ��_�0�
|���М�߅ސ�ѱJ�zn`*����+�kNTf3�5J�����X+m�����Ndku/���oz��|9�éJ��A�R3ӥH;����y����F�vc���=�L������ǯU19?k�k%���S?QL���t��6�`g(��ay����>�Zi�)�O|�����$��w������}��k\Շ�xͫ3H��p�9V�3[w������B����`����=X7�I}����o3Clc��gR�5Ff���
Os�2bZݙ����d�WI���"��S�#�r�L\���"�4�� ��g��YѰ9�Nxs������	5߀�,[�CԊ,����KΡu����¯�0WE-Y�����$�Q���!�����ނ��da����;�;O����8�yu6�O�h��l��kPГ��,�O!���9��2�!FH{5����]��Ҡ\ŒLN�պц�tB��$)ɛN��T�Ջk��C��0����u�!���|$ޤ�b��w�ۉ��3׌�	�k��{"/���w���1�ك=�R�gk�_{PY֠��uz�1�K�c�}[3�tf�.J���Q��+ks�h��@=`D�B��Ȫy}Z{��+v��VGj#�l��+Ύ�ayQ7�)��Z�~L�,�cW	:�%�Bee����u�G\;�E�wQ�d�+���,�T���0+��VH�e���37j,��ж(]��������7Γ�3xO��mN�k�w�E�0�dxE�������'��J"���m���c��i��k�~�t��/�^�^.׭W�����L;�1��4<�(�yf��_-�[��Y�f.��o�ۓ��!q�k��Y2�7��W<�U_�{_N;
ۺv�G&n0��O� b��w�"g�=!��G�[����}��	E�m?xa�r�B�б�������<d���FOvv����e�/���5,e"Nd�K\�\�����x`��h҉k\�>��Wڷ3�nM�gw]�޼D��Ka��{Vv����f8S]�UC6salcFb:_"��W��j�؏n�O��wO6�N��h
[)`�ˌ����S�_f+�ȕ� �V��q����øg�}�sI���
����B����>��[�Q%��DE�u��v֬^�3�'tN�U]Y�*=N��Ë�nf��w�/r��BB6{^���N��G#}%Q��`>ذ�lw��nQ4-���W���c���NCx ���=�[CT��RD˺�>��=o�C~���J"��<ߐ�>��bL���A��箶I�%�Y�x,h��������u�|�~ǕrKv���_T��=^zb^W��5�+0k���>ۋ����U�Ƙ���G�`�՚�k���1T�X�4���%�`L��*6�Q�;�r�>��UL$DH3y�j�qX���e�b�S"{G���r^c�����qy�a'#DP��t�MH@�WuӚ��I�:�#��{����5r�ٓsV��;t�iڢ��4"�A~L���S�qW_�(��Qv��tKg����E�hB��X�!�f�W*�,0d��M�Mj�JR��˵�av�9�C6
{�j��˧V�C�L�\�j=1d�ʔ����Vs����]�6:����Xp����qS.��ݶlߥ� 7泴N$�ݨv��\���1G�������C�%��Cg�x��O�
�:���`S�u]f��P�o^�HΖӗ�1V��� ��o�dS�`�6#�#�1<ac\���Nf�]Q�_g�zu�v��sݙ�=��0<5�{���E�ޓh���H�|t�V��ނu�G\��*��gGH��z-
��5�da-�)��Y"��v�Y�V�����N������>����؁�>w*_W۩wO�eү9��c�C\�k�-!5S>K��7y�˧v�Ul�����zX����T��`��R����D�i��ff[Ma��K
y^�sX�)4M��-d(��<3k��'���=˧�,��N�A��xʰ�T��Ɯ����|�{�S
��vK�T�uRCa|��u��g����CUaDm�ܭWwO;��T��~-o�E&>��Z�}�Cʎչ� QeZN�ڛ��L�1U�kc9V�����[�k/��-��ʙ�g�t�\�q;�uv9Aqm���|��x��DӖ��'�^\B.K[����v�^��#���A����_�
�I���-�댺��D��q��t�>��@�H[��㗁}eL���WgĀ>��v,)����������KSMU�����'y-�"�>�$q�O�6K:����eO2��:*p>Q}��Lԭ=��9P�Mg�j������ �Z����U.k��'�K���<x�� �������a`�?]��co4.y�;涑�y+ӂ���wh�]��C<b�?ߵAzL��������H0�����2*s:��xSE%�����9J^;�����k`�{�3zN��]�մ+�ժ^97�V<5,`��/8�~� x��/����3�v��~��$}�{ӗ5ܯk��Wd��<a7�����U��|S���C�a�Wgon�L
q5��h��_GT����:��u���՟���?����q -]iX���ڬ����jk@�U,fy�Y�u����{�S�q7]��y�V��4L�9nv�Poe��G���S!�}6�����O��{�B�z���]n�S��D'>*������.���1I��C���ݻn�9�NG�{9����C�
�p�k_[��H���j�s��L�9&4MwH#h,�!����ߧ�牠��".��]u��b\��^^Mף�c�jݳ�I��Y��΀`a��Jޢr�x�ۃ�V�S�E�n��xfJ���dBkGc��F�ZLl�̯6��y��;�vt������t,~�@oa��������e�O�����?�\�v�n,W�� ��so���M)����b�$].�j�F�dz�Z�Z�}	��^�LH5`-y��c���sE_�����)�\����{��7C�l���}f/�.LuG.��	H�'�c���_kl���QJe���o��T��.]Q�$]G[2u����G._���G�,}AW���P���67*�_jY
��u���������5�d�j�"5'�-Z#
MDĝr���D��gmvs&f^.�i֮"��[�dc{��o���;p��(^�2�Lܷ�����|?
h�UB��T�[W���Gq�.�����;u�Z8R胑���ۖh�w`U��
�\�qP]}R�c�#B�2\�U�E�f�*��P��M�
�k/U�x�M����x�H]��(�Rm�;s��s�m|r�����g�VT����Nm=��6o��2u���ߝ��K
���X5�邕jN�00ٻ�p$����#�^���Q!�EK�qP$�R�`ŵSs�)�}0��� C�ᤰ����t���k`�2�yҳ_'w�P�OcXi��űn곡�3Y$�"�hE� Tg2{�[l�1�8u�R�k�7��i��@1���Z�0�Ի���e%͓��U<?c|��)���*�kA־@�0���� aA�x��ov�ob*������t*;{(Px��sI��s۽T�[W�����6w�u�����nvW::�k�v�j�vK^�Q�h>xX� ��s��L\�7���F���ǲ엽�r,Jx�Z5`Eʙ0j�p�h��9��'zS���+m{dt��v�}N����o�c.��o�g�M÷�H���Rr�u��w��f,Y�=�q�2��@��\��Ѽӳ�����I;�@�Ot:	J�rV<x;$��7K<�	�-����/�����O7rZ�[��2�C��S��n��ґ�%�j{f�f<v��]3�K�ܶr��]\K �)}#��:󒅥w
�t&���s��2����5��2���\����{NQ�c	�+S��]��]fH�ۖ��v�!tS���R�3	3����L��K
NE�[rK;���6 [˛C��3]��Wٙ�GLqf˾����s��ol	e�[�.f�ӫx�KI \���u�2Ů�t�;Mw6sJ�+�Ej"/:��F$�$�tn>D�1=����oI�o��th����wN�{������Ѳ�o*�P�eNʢ����48���;4��6��ޣŬ/�Vg'�*'t�����tT��T�����uU��^ْ�lv�����VXy�A������7ϗq�ۨ�n����c���G���9�rŚp�Q���5�R�^�Z��e���J�$u\x�m	�j҉7o3����U����&^!O�#s,�S`���� ��a��N��H<�WR�mZp�-�"����f�=��д0�_Q���< �ԺVMyC��4q�]Ne�q��U�r�.ԣ�9���[]�ZN�5��䮗Q��b��$YY���4k��0�������yãNh�)�6��=����o�(V�Z�N5pp�M�[�)��G�>  j\�QL��,��aJ��O��c��&���.�.v�X㮼��s�T��Xz����s��`�c��f�;4��X�\3���^Ԑl5�:ϧ9�n�j��W��������W�:�4��x�9X�v��1�.��5�y�= ��Pz�R�Rҿ-US�c���v���m��R��߷��4�h��h�g��4a��:���i�y��q�oS�@<̑��?k��h�9��t�9���B�龈<N���{T�aX2�����i����۝*J���=\�18�e�<�<K>�\�U���n5�/��G��S��b��R���Z���U赟�Z�Q&�@]V�������dd���m:W�sW�Ä��>�y�l�ص���k�;����R��ޞ��[h׌E�P�y[Vs\c���y�ٽ��bY9�#HO�+��d�Wa�0��w/2zn�ʝ@�ɉ�J�����U�����?]g��:k�Ss�zn�����;�윕Bt�i��X����k���ǰ��+�)A�ǯ�zr��;�̘ޟIGyq��]����ْ���)eD�Uyun�a��W0F��Qj+������s8�FVuY��,X�r�"WL"&���1+��'z�fǯ��Ӆ���]�de��(�|"8a�����c��Ӣ�������FB�N��:K�u{���S�ë���ûf�����4g_� m-/kN���~~v7��TA��Sa�3ՙ�ߣ�ƍ�/�$2,��'ވ�Ȇs��־;�~�&O�>m�m��^���'��dF�޽v\�en��&�����!��(����0>#��C~¶�Z�,fY�7״��E���7��66Y��]Q=�"� �p�NVu�(�.`R
����k&���7l����05Q��1tD���.�u:�.�k2N�F�����˼r@��0[:�9��4DI6`A�ȞaO��+�d��٬�x~��HL+u;H��;Ί�5v��i���ϥ5���_T,��աخ���4��F�k7��q4*cT�&�s��v��.oM�C�����$�=�G�a��/L���t���T���u���&�3�Y`x�.X�?$̡N��{*8�˟���+�_�]��Ћ��q
м�Ol9�〩��JEd.��oՂ��ff��[۸���|gA�.��fF$4�{��n�MM�����ϫ��|�Vi����"���tN�n��wi�]�5B���V�d��8N���={��D��\�3v�9���־3�3��u�{�[Kx_o�̢n���|�ff(��T0$��������׉�M����G^[�Q��7�ɱ&Yde12�.���uʊ+]�Vl���DS�f��E՛rW&��E9��wÐ&.�jNX�H�2�kq�mn�R�F�����w�������p�z,"��P��$������:�N�Dĸ���Y�簐�S��M�(Q�������R���|Sq��!,��-z����X�Ub��:%��F�A�uD&��Y�fn�׵�.���Ԙ!R����]�@ӦK]Wq�ݣ��R[lSkו3z����ֱYO��͑����}�է�ǰVF�w��R�/a2]��I�8�g�=���LbC5(M)�glf݄:D�>vc
}Y���vEι�!���V�Ff�4mx�{sS��9K���e������J����h������>�z%�eQ�5B$��+}s�,tH-gE�.��U)���Ht�.9�����7Ib����.��1�~�"�3ud�D�=�trԫ[�|Y(K�C7�<��ڰ3w�Q(d�:;����ؘ��x�Ok�����COY]���Y�ҺV�|K�:)Ղ>��v����a0�l��c�g??N�G{���]C���/GQ�wTH�ꥌ��2�q�I���=��8�:��z8��q��Fj�������vZ�|8���F;U��q�=�
��H#A�,����[�kǧ��͐��NXPO�|N^Ut��^o���-��ybր�S���T* 8L�m��o�'.�s�l`zsM0;���xzyɗ�h�S��c'�*Ry���3�������~1���n����&�v�]L!����{�=	�����'�CvPJ�JJiY��5��7��_M��'�.���D�W��b��iL/�y(2��&�h�@�X�����9ҭ0�ѼY�|�����b�+���0�ϰH�%z<KR��r�^�͈|�e
���r��i����$��Ԯ�*8�u��7m���#�0�Lb�Ԟ5W�&�]v�P4��Ch��F�ļ�t��p��t�����\k�9��BQ�����{vD���{bZE�[���5�S��,�V+v����ƘͧL�YCA��aJ�J�2`�2���{���8���_;oӞ^b缦��ĳ��%6^��t�<kiVLӦ�w�^X��\/�x����fm1[߱��m�tZ���1��8!�n��=�WCF�ow78��bn/Gqu��$�B
'���'��؉\^�"*-HV=nn�����ՂT��g]}镯S����x��-x����}��4/wR��/�2GN:�]���1�����h����PO`���;��gj
[��h)yol����V{�f�P9Y����7D��,�^r�φ'C>�SF��W��+Yݣ�f<#��j��k�ѕ�u�G+}�,��[��e����i�X`x�1\�cv��JY]�3Ϊ��dqT��/d��;\�!؞"c���]�V���>��n'�E���Hׂ���~M�q�yX���+�*�E�~g�"$�t��@��m�a���7��
Q�����Ý
�P�虾決����r����xs��~�D�-|6��&��-��v$�^>Û�8��~��(3�؎��dOA�����TDK��'���Ѧ�[���c�&Tuj��y�Eдf�x�6����>&�t-al��Q&�*訖���陰��4��$ ��
,��j�Q��Zk�l"ɍ��=��]�!a0VnR�gnh��+���ǌ�}�V���R{���P�ue��`��)N�;.�ۆ�Dm�������!�0��7O@M�H>����dz��05�*��C,6>vS�ƨ�X3���nZ�Qc[��D��A�}�Y�1e<^�^I�&\"L��-�⨎������Fj�)n�RC�u%y{ ���|�"r���'J}��͡rQ0\��N�L5�F���.�^�y�V���1�������t�WR�1�KZ8-�х�����(�!gn���@&�=,�,�N��u��f��;H�nl����_�E�Z��bqvDh�]��o�r�:�px�qD��%Mu�%d���.z�����k�]�x���7>��sc��y����3��Ow�'��6�nR�˱;B������d��2�B��s�~h���pj{��\�y�>��N�[ձN�[Oek�*��]J����Kٲ�c���?��u�{v����W��H$�;ʧ���K�}�{=G�FER�/&�[}�o�m��wT�'�$��G�����o�c6�T�Ly���U�	rI��%�Yu�c�өT�k�J�\�F1ŶF���������{��{��+Z^�@�K?����~���ff�O�R�,�j�ݛ�,`m��u<�;���\�t?�'L\R#OHy
T&��I��x���Y]"�~l��݌�y����'*u>'���y�)�W�_����|{d>Cu�^@��t9�)�����*a��ػ�E�Ey��mmx�Nvm���cc&�}־�n�%����ZuM���T��i"2e\��z��ߡ[(��^�=�$5���L�[����ڼ�����tl9�Wj�?A�e�%^�Ϥ��^x���]�l%��Yy!m���-��/	��}����Ѧw�S��Z�;a3��Ad�'�=ܤ�J�P�jĊN�۵�5F��Zu�+Y3����X_h��P������kU���q��v+�� f黪�R[q�+�G8]�8N_�E��!�k���"سd�hߌ\����P�����^�.�{%x�+5c�C�����_P�+��S1���@ӏ1�׉cA%��G���&Z5�XxZx�7I�=U�j3��}I�p��ƞ�V���:Ӽ~�����އݮj�<����c����ۃ�R�{.:J:+�J�X?���/q��.T7�N��M��D	\�6U7�差F��
]���d6���<��v�a6��V>wR8���ں�t�9�XGzuյ�C�jC���6L���W|>JK��k��b�1t��f��GM���[rm82{/F�:�����N`E�N����ٺC���ǂ���|.e9�xw��9k>F�iPȷ����3�x�+_'�7(ϋ�aap���ݬ���o��(yli�T�u\�F"��Uw\'yHEt�fq�mS���z��{�W�^��fd�w�"�*�w�؝���F&q7l众�f�᥺'l|0ׯ�`Z��>g�XZ3�`��:�f"�"#���O4�8v�x��w�z�N#e�֐�%�f5k��Y^�o �F�<�jk;��M����UA���~��A�i�z���}��B�{�0�eG�j7%Cd�I6e�5�{"s�o*m�	��E�僶��n�K7t)��xԷ����8n+j�?Eg���Y'�1�u��ݽX�;e�aI��`.��N���O�{�<��f��l�%#=���+�{Q��}�cy�	��]�=Ѓ#|�Z0����a_vv̗�є���q9��5���Z�����X���v-�F����.�]i��͉F���˺u�r����A@ڻ�:K������+�����C�$G� �ږ�]Z�lf�U���%�o_aχ���������Sݔ[#>'�������$;S��W�\b,Óf��z^]//7�ݻ̷�V9�ܺ�+�=`"1^U��y�Nj�>._��E쟿��J�뜚�5-_3�L�;7�R��A�+�d*1����D�{�k�My�gs��c&�f���}�#AZ��Fk��R��f*#���d
�6}>��d/�\����bz��p��s��)�:C�nQ�(���Ji���|�O=y�zN�t���s�v�OE�o��\��>(`�G�b�LոK\>���ꚱpHx.��y	3��zAU��5�w��4X�O�vRv�^�s`m©#v٥�0po =�q�ū�M)꼯��`����J��J�6�e�za|+��ެ��|ZΖ�Ol��������I�>HC��w\���Iu�P�_|6�L{w��>�F1�M4��A3rĈ�}�u�/
����n����i�Au�!I!�Y��%_���^�R�4�A�R/��+9k������^�,��%I��oM\&��sq�V�5	ptøtA����w]��LZ&b��]��r*�+\�g;����bwA�W��KJ�;;c��z:PƊt3Ou9�&�[�6���Y�ЏvVG�6�x�s��qޣ9��7���6�O�KKV:���N�?/�N�G�A,Mg�+ߒ���8�%e�d���YV�Gm��2�[es��q��w���[7����zX��ݟ��z?~�����Q�ϔ��n�*��t/%G~�m!��n�s0�@&��b���4�o�fuFGb��$�?X�b��߳Քg}�	��Բ�@ȫ�� 	�Ż���6"೫"N��,�7.|ђ��ګ*N�u^z׍�yV5Oܤ�g���)��ym�lVR���s)�W��3�YBp@�ʟd���)��]��t�Lz�x+%�٥-�΁�}��yu�7��򊶻�-��f��x�Ls�̃�ܩ�q��R��Df�w�A�J��=��G�T�����qzk#�ɵV��!��3q\���#�������POHK����w���C�����oY �,PJ��se��{�V���d�\)5t��k(����R���i�Ed�0���,�8�U�gD>�.����q���x��1���%���]B@�Y������w^���@�C�¯C!�����ݨ���֟]G��8<�A�^��0U�hl=��vt%f��WJh���;v��&�cE�wF����:�hC����g�"�e2���\Qni��m��0`c����^S��j}0����JλmAى�թ�{I���K��3#0[�f�S�|gÅc�Rjތ��p�6��e����@7��o|�|o>�N�.X��GQ����$���Vv|~��-H;�gWJ���\n��*jF��A\�䫨�&)��畻(��'�%�}z,vIQD�}�Ȏ[�ߩ�v����s�>�?o���iV7e~љK�|����s�ky�����3̅@Q��m��RѺL��f���%)R�E��,c%j8��f\]�f�S��7�t��,�^�p�c��A�ЂK���C�+�b�]��};��(L��#�����pZT�쒤wpb[��Ff36�>[�Zp�X�����˒nXb�.�ʺm�V{7��І�ޖ䮝XFn^b�ᒜ��e���U��mpL�v+Ļ�,�œz�}�XD5o{��3,6hP�OH-��2U��g�hV2Rʬ�X�ڵ"�W���*o<*=��}Wzc�]e�nmZ�h6N󫚻8�i��Ya��Ц�|�q䍷�>������Z3��;ˡˡ����7`�*;3Z	p�1d9�ǀ�^b�.0��گ{t~��b��e��qǲC�` Z3C��U��2w1l���}ۃ"�������WL��АxG\�Q��Nt�B��ѡG�݅�1�<��e�|M�Gp-&���0��*��%R�oz6EFTg�*��Y��j!��3dن�]���'G�"{�N���<+����Y��A �ZlJ1*89G����\�3�����(�bG,�q��h�r)|VLѽ9��B�Qކ�y��%�J��v���p�j!��W�:"ggU[�v3OF�d���
�pi����#������c�����u�ʳ;Eܽ�f�̨�t��ۑ+�s���u|�R���N&˰OD���Ƹ�S���X�!S`�)0,�=Iɕ%��8
�ƝΧ�uD$o�uɞw2��9W�7Nml?�l�q�E<�\�XT%��\�c�y�ֶ�WL�4��O�S&��L��.K��LUxJ\�ƶ�^� ��:���0kvd�9�	޾��Cj��](g+*�.�F})�`��T����q�-~v7HEʮ���f4��n�I%�஖bbj�U���P�x��-��o�H�[�y��H�x1�(l�COX��תe�ƮR�т.�r�j�\D*��|\[��sƍ��E�)赽X��Y����j��rwh��3ڍ�X�&�*b.���@�{� ����.����x�Xu�J8^��֞ld�ﳔ�E�iN��4��,���[����e��0׶6��}�U3��l
j�o��{����Fj}�ƨx�J9��:�;{�ZЂ�f{;��}��ͩE��{dY{�\wImlb�C�2n��l���G�]mCn~G8�V��ߝ�/�ٱ�d��6N�d�YYT0�^�j׬M2��V�*�]�s�/ު!�t��/K{o��iRCܙ��;ub����ڐ*�ci�N��.9�����~0K<�cǺv:��P%���S�ؕ,����MpPPVnd5����$�����e�le�
x`ٴF�Ӡ�S̓;f@��'gG2�1�]�C��	��*���D��vm�|2��5�-O�~ܤ��Y3
�(j��xދ�\Ԟ�(�����)�@������{�p����{��/��W��~���C�s��'v��(}����$6�;E4�+Ϥ�dp'�$�zqԘ�w���m����TTja>���Z��1��<�sA�&��X�S`Sj#�}v�_e���\u�2n3&��s
Z��1�����[��	
��[h�]F̋8u��.9S��c�y[SE��.��᳃�=Σ��;Kph=�l������t�Le�egL�TUl�����A�D������ �Պ^L��1�bpx��gտ}D˹�N�60�^�ʍ����"-��`�� ���Z�q����F#��,��尶�^1[���ЬSM�'�z��M�q�|��h5iħ��ɿ��|-��uCv�,*)��mq�窛��Ek�-䭡��9[��c�&څ�; �����u��D�/{��.4����6'D���.l�ǂܶ2П�)Y^B���VնM�<�@dD��W��cd��{�k=�N�Vb��Ǚ<�{$[V����<4j5o�Z��=c���w���*��D�j��s���rr�K����/8��,7���Z�6�#�cJ�ef ���\C�Ȥ���A�@��VG�N�[�k�>f��S�e�����19�mu�V_�o��6T���\'%/I������{x��_K������g�vC;���ޱ齧�%�b_�-���~!����}�f�HbϵѬ�9��j�6�-j2��x:O�6��A02[UU����X�5y�I2i���o{��|�k��Y���q�������:��B7����oi����UA�pX�wVfǸ+��-urY��ʇ��ֹ�$�]Z���bL��r�BN���;�m������Mu�{zO�x�1��Ų�g4S���oQ���i]Ԝ�X���
�����<���dDe��}j�U�}�6�4�ܓ5�RSx\�js&�{#nIo7ԍ��ߠS�v��ueH��K`2tDE*$�,.��99���,�b������r� �E����1�l'����3GE�a]�o�xN>ν�{��]1������ ��=�ǡ_8�U�sb��/��<)O�E�W�~��0�'wc�"뱟���C�vs*�����fv]N�Z���K�q/�{Z�5Z�>��_�X�/���_��R8$�|}�y�ݱ�Y��~(>�N�+:Ʈ��|N�'����_�����$i|.[�*�#�y�O���ʄy"��o	��º<1��T*ȓj��G)�W��웫ך�HR�c�A-\�j�x=O�����B�Xu��%6y���X��Ҡ��U���!5��>������u}M˻�LY��Z+�+4kY���3�]��B�J��.�	��3k�y�ɝ�8ų��I
��,:�/h�]�g{v�6 x2�ƻ���b�R��Q�da��s��k)��83貔�v�aɖ���ͫ�,7n�����t�U�'[8u����K� ���z7*�0�VW����oE�vT�L$���.vt�Dɮ�w6�޶'$V猓�鮺�k6��dCnr�'"^��-���{�^_}�{+�z�o�#fz�.��kH�@��sD�]��P̞���f�Ur^�%V��B{+��!���qE�zF`[�E�y�X�:�-4W��ʵ�Mr|G���M���-G�V�V���"�}��'O1�)��-N�.[��=�w�'�o�?N,�| H�h$T�yF­�g��7����5HӴ��k�|sU_,O�� ���t+�w��O�[�ϲ��u�A�"L�>�x�����n�I|�^5���c2KS�6g��}�"�G�2)���U��xa`S�~��b��և�z�K�q~&�,���R�]gA�#�kq���%w��򎗳�h�e:�:$��6S�#f���qQ]���.b	|���4|�d���|���)h�}�є��S�5���s[�i�
���y���� Vic#�j�+[7��j�qb�C�$�e(��Z���̭�c]����9Ѫ�h��l�t�L)����j�Lّγ����'����7��6�b��qګ�eO|��qWCd1��1�Gm~�=
�G�Zr�����r��/{^�J��Kj�<VT��G�>}�W�}��U�d���z��Vq����L'ٽ���U1'y�3{sn���*/&̻��!�jn��r1
��>�v��&D�is����D_��wg+���zy�啠�;�J���l��Ϊhʠ���!�8A*���p��������kt>���tf�����C&:gWd��d�r#H�^���n�.u�kR1gp���.�r�u)ia�ˏJ["2%�ިl`O]�I��g	�^���O��� �3�#���{��*�1A�����hzt���������������FO��{�/?{Ǳ}�A�Xv�⚮MrS�q��r���wo:^m��b��hcDF%�)�i�@w߿P���Yp:,n�b|q]Η��S�iK��QQ:b�5�hT����_W���s�qYo�fT��d�o@���E�]� �͋N�ʝ���{7v���`J�W�6�~��%E�tJ"�h(��~��?�f.��/���F�/��>�<���u�{.�r�!�����.��` ��;��pʔ�7�ݯ;����:�� ���{ۢv��(��i�s���ֳ�3}Q�^���Α�h���C���	�]��y�����W�����*��&sow�������|�\p�8hy�l~�Z}�z��T� (��qz�V%6��TW�C8;� Ed�.]Z�7fC{1ێ�OJ�l��U���p�\���뽪B$�������9'Uj���}����_ `�-��>MP�;� 9���K��{�6L�o!�>Q���O~�jmU�YG}���f~x����'��FI���oMF����ؘ6{�̯R��Z��ػ$���jB���_~��O���%����Y�1����z���!q�5�Y5q20���� =U�W������F�7˼ᝩ��[^��>��_��8�R�wV�>�#���5��{«VY��T| �9�u�,���.�$Y]��P]RM/����3�}�����{����	#ޠ��}����DƃȶY83�R�)a?�gY��M��o[�g0���7b@l�n�y�xw��7�|k��ﳨ'8�̶��,�U",�0bs6x�?/o~���˭յқ��3,&��WK�4M���.����;j�P���rd��N������uz�]ͦ�L9f!�eE�p3}��m��:��)7�9�;�"��v�Z����{���9��x6wB��IM�%:�<�x������p�O4�ɥ�J�9�������r,%�2�����0��s�p:��A�R�ma�|����z��1�'�YO�a
Ey�ûc�϶��)�i[���U����F?3���Zk�]�N���g���O.ciQ�)���	1�E�g�4y��r���9�S;4BK�*��~ޯ�;�_�hK���o��[��W�E����u�Q�liC�e���H쯣*ע��|>�?Z�c�����ՁH�a^���K��¦1ݯ��\�] �O���ڣ��sФ��ZuGXe�^�����c�6� �;��ikc���\�>�j�3���SϾs{����!sӪ
����h���Pm�<�M<B��ݹ�w���t��w�ywU7����.
j$Hg�q�I�s}J�	>�e-�"�1�&�)�<t���Pو�X���TK�N�^!:�0�;՛xb_�_���q7G�峗�-�VP4y��L�nWv9+�Y��X�H���"
��(*�ͱ��֓����Ӯ���P[�����I�˧�N�S����;��I˟cF0�m{T�s��t _zG
'c��A:nU��ĉ��CTb�nR�;��=�ՠ�ݔ��O��m̓��ڑQZ ��T��N�&����fcY����͗������S���=�`�SS8���W+yxw��MF��*��J���=���g��)��m���������K==���\�͂KX[���F�K�h����>�w�|��Ɉ�����`���T�'\�WV����m��晕t��z,ű��d��:����2]�^O�r��?~�(��^�nحi�޸����g��;�G���o���PP"��vd�������b��54��� ��v��S��؟F�~�T��5�2�Vu�]�l���4"�M6?B^v~Y1u2bf9�#�rw\�f��-����%�m��q��[�
fۋ���4��t�` ���K��٫�?ϖ�z�o���|�&�{��!��6��T� �r��{	��}A�!��P1�֞ }(��&�QGĄFC�ú�ժw˿�����։sjf@��ր�v0�ilY������W�,�LZp���5���VCD�^5J.S*d��-��;e]�9X�]���v�:vC&Ed,�uc�����i���@�w�ԅ
-�lxya�"[�&c1/�D�<jS{�YdWy��v!�j Fa�ÞK��p_�M���t��w�Q�G�*"vH��g%�U.�:���GY�Pک>�"h��6��8Rf%�.�)<S�Xke<L�\䯀��0�=�vM�e��T[�R�nK-Y���p�G�a�_ynԝ�~���o�Pu"S��BԌS1r��:���劓u��>!�zV��B��`�(��Ctw�����<��6��O%2��p��*�����nmf�oޘ���kXݏ�c�6[�`Ҕ����+X��)��uy�)�:3�i��E�JCNq^�X�نGtq�;U�vn2 ,���7's`��~F��ǆ�@owC�����d��M|��w8�c8�R�;fpƛ�0��GV�>5��tI^�/�g)_���'�2NZ��k���Fҋ/K�F��v�6������jM� K+N{5��,-P�Xԭ��vYr�J�,� /=~�>�s��!5l����Vv�h�­a]�bJ�������t����+&��'KdүM7}���c!+o5t�[��Tnu�Ix�u����2R75Z+J�9`�f�'UV�	���!��T8[�#��0�N-��z����Z�!u�y�O7De���SY�OQ�aԸM|������^�;�5�.^��Ty}f�ƞ��m�k]6��bڽ/>�ʬ����G�C�~;��Qv�<�6�4��n��,�j) �t<u�I�����#�|�������{��>ڪ2m
��P��x��9���� �'����&tS��t\�r:k&�U���U�5)֪���&ui�G��w��(5�y�]a� ��?n�-_{�3��J�"N���dZ��x�}�y���'�]k�W����J���$��Ro��-~�v�;5�CRy)�;Ϲ3��
��e|sյ��G�	#�6��U�3��N-���}��hoqlr|i_,���J���w�F��A�� O>s�!*�Ww�B���5��l�%�I�aq:E��$qpQ�N�h����e7x��:��2`Ք��:�����r��}�������6�όze�X�V���S�|5�qW�F���)��"�4�,�08lh��ө��[*Я��WgT\�{��Vr�p3�=�]eFV3�o~В��!$�������B	�kB�ݒ Bhd$$ 甐YHT$ B���!�&@$w���!$����M���!$����}���?χ�������a_�����#�����f�����?�Pr%/�ż�e���.)bik9����M����
��)"��X�Y?2�v��L��5NljV��؂���?;�$wbzh��f͸r��TM#�!e���h&�6p��fTm)u��e�y�:�rV֣mR�$&^!����u���Z6<�N�F�;����
�Yu�m�x��J��
bYvf�ƍ�H�^�;gU\�����T�P�e�Mʴ�<�W��TVb�92���ٌ�4SƎ���̺�U;܌��ʭ8�rcyW��G\�f���Eܫ�Xq�.�l���pe�v^��s �[+(�,(&VAL�N�{��z�y����`ƥ@D�U�Ue��٦���Ɖ���ȶ(�]I�d6+�����6�MS,�X+3Z��U�L'
l�B�xK:��VFP��
Pf8:��w-�%��4k�T)��b2��P�ʬ�nYX�f]+�t���-�vC(Y�3Idk��t��x�3��V�9�W�j��&\��~�{���BGfLӒ�E�)Tzd6���^b3v�bѭ�JŜ&���e@[l�`�2̲��fC�;�����݌[�G�Sq�4�u��]����wkf�Y6L�5<9�?ajE,9�6�*SIO&n�M%Z���m�������n-ni��N�]��ji�r&�X��9%3�RB�-U<slK�,Q������[�`������v��xr�V�39�uy���8k�_�[�64ٞ/�U��L�r��ؖY�uoD/ �R�*]$�i��'0�x��;�%�
TSc
��Y%ڽ�-EiӦո���"˯�ʢt�&�Q��E�<�LǙ �i���4�㗙6#�ہXv�S�׉���\/s08MPY�h<�]?��5���l��[���2��w�a�tv���@���i�������3����@�$�d�� F� $$�� 2�!�6I$�BBB!$�d 	� I! FBI ?�������$$��l���3?�B$$�����������		&�7��!BI�B�����@��w���!$��\��ߵ�٣P�		'��!BI������!BI�`�		'�������w4���!L6��������B����P�		'?�����d�Mg�t���f�A@��̟\��o�����@�CK5��j�R�G@7m�+M$�ڣ���i#]
�"TѮ�H-�J��T(H����U��
S`
��UTP���(Q!Ӯ(H�U	J��m`
#YTZ`Tт�P�UZʪ�T���I	�%JP�kh=1QBD�5-j�խ��1������=�Ү�ӧI;.꫽���ɥm�m�����j��u��]w��n�%���Os��O��wM{b�D�WM��@ � �� �P �GX�[����:�m��n���˳�wqŻ��Z��覚ݚ�L�pw+ik+Z��-`��p���*��Pۢ�w(u��]@׼�7��gN������@=A�dz-Y۹���ð�ޞl�Yx�h�8{�U$����=۞g�z�0�Y��)����Ҁ�OH]+��C��������׃�^� S��J� ���R�=��u�O\ �G��@z�׼ o\n��Q��V��su�A���]�t��W�{�������ӷg����(�J��G�vt���h$��h*���hG����p`7���cA�w. h\{{�
:�y��W�{�� m/P���&��+�B�c����xw�<u�4^���E޽�� ;ǽ״uK�<��Jn0�y���˃֊�溭�b�f�N݄QSVҥ
O��[��U���z��s��9������x���9� ��V��x{������@{�z����^XkO%TUu�P{���*^7OA�w�.^����=�g�hz�]G@շ�y8U	^������޼�/=��5�w�� �J�����SԠ��{�)���.���{����2ڮ�C��x�(����mu�=�p4��W�=�ˮC�ޞz�b����R�(4b�6�%* 2 ��&H�  E?5)J�����MU d 	4�$�*yL D�Z����b�%%h+$DTg@��}��{��[�����$I;�G��$� �I� �	$�X�I'� �	$d����{�'��p��s�7v��L�wD֛TnL���hژlA�c��h�e2ջ"���6�]fP"���.	wE�v
��]��>���--�Z�4+uxu�u c(��G�pna"6�1mc�ݚ�,e�2�O�"�+��[a�U�e0�ۻVM3R�Wp�e�X~P믯Y8��h,��M�5�cݱ��*��x����b�vq�Gt+ۗ�qEѹ�yOL$ޘe�t�ۺ۫���Q��;�D�f�V�2Ҧ\��G�74�2^�K��iP��*���f9VıD@'�Q�4�b��޷���w[���{mb۸��㵬��o�wiҲ�
�wh���n�x��4/,�˺�Ŵ/ui�U�0�zs�/L8r�^D��j��^B(X��k5��{r��:���:�(���.����^�C{w��� x��gl�[�k���:/�E�r��l�Cm��զ$h7z��z�B��ݛU���̫׆�a�+3t���+m�uI����,�o]��n���TӸ/K��Eϝ��-�uմj�6�v����>޽��v���n25�~�Sq~�UdSj�6�E����]B��Ĳ�\Pdui��а�F���* i/���\��wg7#�'�J7�0���E�Yw�����uF){N�7ds�m��x�&�h�t�jX3*��+7x��	Y�R2��/�GMV�S 87o2�)&(i(�*��n�P�V[5�Ku�p������.���kta8�"�5A���Pd����DU���A0n�2kP,��M�E*�0M@J�:Ir�@љZn������Z��d�퇲e��2��n��uF����˻ݻj^�겅�Rm�>�<��
�o[�����[�Q�%�$��W��˕������$y$��ȪZ��j���7PR���d ���x�*��_
�/�|�v��`���r�um3�Y+��j�F��KJ��\��=|mk[y�w��J���4+-�������7d5�V�Y�e�������>ެ[w�p�c`��G��9�����)��;vZ9D^Ϯ��5�� ���4������n�m�ط���"wl^u�/V9�̡@�wbP���y��f3n�M<���i+h`F����[U/-�M��߆S$n�cĨ[�3�J��S]p5m�c�+~�.�(�w��Z D��#7[���5�t�EK`Ц�]�
�w�
h[��MRON^�4�X.�d)�,��.V�!U��FZ�=�9ͬ�VVmƱ�f�[*�Ԃ5R0N�ω���!$B�AY+�Wj��n�D���+z�tPsl���b\�y/7���0��RH�ݫ�1fH\R��D�`9�	�zt(�Yl�E5u���8I���fb��-�tE��/�eɏe����X6�����Ŝ�/��]�����ui<V��)�4���Z�o�oL��ti�_Gf�W�"��7je ��՚����rgmн�'mSE�˰�9�7U!,��m��[{�OEB�+/�kkѡ4��.a���Q"to�5��N�]��j�����Лv���㩘+�$�����ت������·�"ӆ�$���z�Em]�׶@�GenW#�^U�mq�֭dkv����Z��;+U�9b����<���ލ:�6d��@��sI�]�)+8~�f��P�Q5���Ҹ�	�'̤�mfem2��*� �yB�O�,I����@�oC�� Bxغ
��k>�%e傦,���b��
�����yp*N��������īo9�a�)�*�aB	y���!��kH%"��Z[k\֛�����Ȼ8�ꯍ`�a|��A�����C�fb�ʼ��LH$QEDQO	��m�[ΉN���O��HLZZ.�LS{@�d���5ᕁU��� �P��$�ڧ4;*�C6��6(ݍr�V�km�̚�K(Z?�j��_l�	��-ب/�F������0�v6�ݫ7H��1;�v�q@��62Vճ{���Mݖ���b����6���l�We�_L�TU�5��@K���Y87h�L�T71����Z�")S]�%C(��K�"��U��k���+%�wu*��vs-��RpT#H�����ܿ����x�i�]�[�\�V�g��K3:��8U�i�kF��&��m����V��r���|W�1�$���z�]Ѥ�#�2�=�'�7o7�1�dت��_V�_�t��0�L���`Q�$�
sh8�����s�F�YQE%Jj/h����(lmT;Yi�%�5�,�sDe��uv��h�	��>}�|�vI��=����:�4z�������{u�PiawCN�#DTЬu_�;*��{w��[n��v���� ��[��B���0��:m�/E�ܯ����A	�ǔ��z�Y2� ^�Ѐ'�_$�b�Z:����0�2�+7FM�*����L���6��-��ӆ7[z�LZ�nZ@����S�Ӄ�����#�lz4�c��[L��:�
��x�<wx۲�-d� ��=E3��u����


˗t��l���6J�NM�n��b�Ue�,��i[��n����`_^�4�P�kSuƹ�t�k[��X�6�:t+�wxI�TjD�%�赹���4n�0Ȅjc�7uYyV�
�����Ǡ��0U�V�]`nK�aF�fAf���n�Rt���ub���kP�^ʎ��hd�b	`�,��GSKnm�r�1����T��J�e�-4�ch󱊮����1:�<�(�� ��$E6�'��*��`���TYlцw����
,,�͏z]sٺU�
��~����%e<��	�!9��lPR���#�76{���"�{G�뺥E�@��aK#�\0�`�=�δy#۾�y��8�+.�͵[l�Ru�˴lS�VnaZ��#A,̻�x���y�����滮u�ㆢE ��#8n�0]��4Q�C7.��m�]�7f��l�H$�Wsn� �~��C��a�W� k)PSv�}o>�v!�2��{V�����WP��m��p^AS!N�����sb��*6���1EqB���>f�v�+ת�� /7kM���Xm$��VŏUU��L�Vi�Y���H`�8F��\l ��Uwr����[�I��c$-^:�6<ߴ*�A"�j��P�H�Ak1�{�v6�g1e��;��f]ӊ�Y��S���[V�Qa���9�'�M((��k�/\��+n�Q��Q��8���h4	qd4�em�n�क�,�6�Z�^�}t�5�SGXmFAn����/.�Gϼ��3]7�nm���]f���K�v����٥L�m
2�� rmfA5���k4@&��T5�ç�
�pQ��Mp�#)I�_�u�CV�WJ��b�z6���ms�0S��rj0`�de^B�UZ�׻yu��5��m=��,ݻ/s�kB�`�:�:Q��,B���\6wJ�RTVY�4'�kL5�&��0)���ö,�$1C)U�Ò��b�Ѷ
0��J�M֬-[+4	�Թ�A�D�
�Ӣ�>n�V4�+�k�X׺9l����Цe�i��5Yuyh�Ģǳ\�u{w��n�""�*""�((��
((���(���(����((���(��(�� ���A{��݉Z�iUe@�(�H)"��y�\�bV�w ���O�TJ"�
�}�k�v�0K�w���w�;z�N��S7q����aRE���o80�͚�}�og]I[�0�E��͖5&�#�3���j�.6>h��1�f�[n�Q��E0�yGo�4ne7W440~ ���K
��wY�{٪��*1L�6R�����9��U��N��^5��Oz�xv���Nl�T�ͤ�m;��}oi���58YYS�i��{�mL��o,\E���ѳ��9�z�А�JA_��y�籽�T�1�?ww�x6�m�j©kz�o{ pBxb""(˾h�o�WZ�pY ���E��Cwy]f#��J�������|���D��c������QdFj�F")f�z(�|r��g%ٽ��(2��R�d�ܤa��i`��t����֥I�;/o;�j�|�Ĉ�0P�ȌFrf`��	teǙ�w����:��^n'kF4 �����/FS�V0�;m�ܽLnV3%��(����Z�u��c+�i��И�ї��"ܛTm����w�Rh7u��B�[��`I��ݺ���K�`�:���Yt�t��_E~F����2���l��r�4r�9�x�=�4����ٵ��s֎��̰�fZ���iàA$A���V��##�vܼ��IfeVkc�-���ld�M��u���鳨6C���m� h�b�3M3^݈�9¸��5'Z�{{b�/#�DQ=��]�����1w���.�Gu^Ri��U�}sZ�w!�).�QDExUl1�V�E!cE���`'	,`�f�@b7�w�9�y�S�G9˻y�^�w� �g����2��m}[Q�em�Z��v3+�&l���Y�`�Hg�o�vs�3͊�D&�JQA�ʶFmAe�
�D'P���oS�uz��oy�i����Z�+X�9�EL-Q�GO���XB���f�(g���an`��k"ܤ5��-�w�v��̺�^F˱;W��M���ｓ[V[g2!����Q��{�pjP���yb��5]�T���
��Rҗ5�B^sZ'<��5��m@� ܧ�i�S���zN��u5��Ɏ\ ��a1r���cRIM�F5+8ʨl�@�[v&�L��J@u��j�m�A���3m�e%��ܘP�!��^*�v��&H6�]UM5[�a"�or�]�i����&=��!�u�E��5r]�_�,X���n��ST�E�e��g5uWW�eﱏa����r��r]��C/(�O�5��h�7���IM_d��g��,њ������5�1���m�V(@�P�_|�_��
:~X���zT�LX&,Y/(��t4^���F�a�*�4-��$�/U[T��P(I�+7j�ٗz3Q�6�0&�5�V�� W'��f֕d��x"�����=���S�kn��J6/l"�����s\�����F.�|� s�V��h��Z�Ga&����@�sA���{�.�'GnX(V�;��Au�n�v�U��d(aX�3j�iR�}KU�Elc>v�)trS:��p�0(F	)
�W֟#���C.�,T;,���/v'fK�8v�V�.�X�����Q��y2���\���{f-�b��v[���7{�rJUZ*��Cj�x^��c���٭3gZJ��v Z2�a��K�F�U������6��:���t���l��N��|��@ɛ�e��B��vEh6��[�z �~��&��S������Iҥ*SX0n��In���� �A AXh��� �=�x3x/u�c����Pܱ�W+gY��N��j��ŷ�������Oo_;�7��c���cᖩ+tl�6�Y��*�-ͬÁ}AC�E��5��*ڌ©�*��.��TyrcWd���d�55��J��uv�ʣIdf���[R�e����r��d輾%���Z��*��k�l6A���"��;W�DљU_n?�_V��gn���Rq�Aꍜ�����%������B~��Z�azA ��4A����:��3Xq��Y����E^[6�-","��^��*;���
�����8hf։o�#:I���̪Ж�X��#��
���w^��.���Z��4�X���
`�h��$�&�8V�a��v�V��Vr�jC
v.��6��gH�nX�*��
b\7vkP�i<˕��q�sM�Ѭ���4������Mf
�k�7LJ���Gm��I�:&^-����%0�L�
�V�kt���xݜ{���h��0T�M��.�����*����#��$Y��ǎP�L��b������۠�|�m�����T���lM�-^�X�sY���4�%���JK(]K��ۡ��u��_j8���e���n�ىv�6d�L�َkE&��x"Ũ�3h�1f*�=c�/ݭx�4m��v��!��U��n��on�����)�P��q�(h��k��}�έ[����o��+=i]Y�^�� ��E���[�������n�r=c+�Aج�"5*�5���Jn=�n�*Ø$A���5w,�Rc���&��A���1�y�e���`��*X���E2�E�è�:	���YMk�=̬Ҭ��<�3�+ٔ~�tQ�KI��gB��Ē2��"�t�a%W(1/j����P�3>�<��$e�l�V�h�_U��wr�d4�H���؅��F%�Orڬ��anŋ��A�b�x�J���^���<�	F:�sfV�ƺ ޫl�]�m���+��h"^�b��uPI�҉j�LҎfXM6�ⴇ�7�,�f���`,���4d`I�ګу.��Q<��>!�qK<X��n���@�ʮ��y�Y;�r�V�^ц�ϙUu�n�R�AaFE���]iWz+s�oR�EY}��wh�W��4��ͧE���m������uGn�T�`��� ���&S���u�/f5doC#�(��Zrs�V+�����o ��o�fC�t=���p�%�<�s|�6u�>D�p��|����g_wwt��ˡ|ζu��들xNgu��qNs0źY%4���bQ(�$��Q�\��׺���;壇#�8���!{���e��6s<�I"N7B{v<'6ru�e�-N���aqy��2�	��v�ӱ���J=�6�m�Os&n�]��]�%&���L�aPV�ҵ!'y���*3LN;���Ges�����&�����w"L:�X{m��}6e�s��ý��_,xE��=�ZQwF�u��n��{�[��I�ͤ�r��v#|�Zx�W��� �w��٦�M׺gH{�|�P��������B�1�{�ۃ�-��tԖ�]���]�����J6ҍ�����G�<�YP������D�-K�Y��y��ř�S5�#�H��*�mi+�b-�ܺ�wa�������sz-\��o��p�\[Ԍ
�/;+�����gi%��nr�ĒT�ށ�k�LU�o{
�5��w\�9x��O�t�!��ӌ�� �V򚺭�]�ft<�-$y�%@�/����ǝݻ(f�x^�����	�i��=+�O��&�+R��,�{1cʒ�u[�b��Jxe�o8�9�@�,>�D�Ļ�2�u+9���`����)�sn�)ܖ��@M7e��v�ɫҼ�f̦$�w)��-���A���u��Q֫o��-��[���efb���ٴ�%'���ucxm��ͥ$\�άw`�Fk}�BB��m�^,]��\.^T�V�Vt�m�����ʇj�8�(�-G4�}�gXȤ�z3d:m*�硣S�`x�	*���g������3jcV��"3-�`L-�Zk�%^]s��<�^*������l��#�k����s���=_֖b����S����4C�7���:�mq���+�\!Q����(���Zm]O^�tf\�N�vu�:��]cN��k�h_-3$ k���{�&�	%v�ْ� ���E!���b�V��|k��%,G�����P�]z��rݝ}`�L'�/-����>=����4V��1�z{�+ m#Ʋ�XTkÙ�Տm$pؑy��혣�]�&�-�V:�y���q�f#�"I> tmku/ �kd���ub�e�)4Ik;��3C��V��@o]������I��ͶU��ew=�wf`�0��&���"]ùwo������d���.����Ry��)��Kgj�`�ֵ�XZ��)�V6!<ڝ2��v�1��!�8ꔰ,���Y�o���F�fov��(3en�=y��#�oX�k��{��i�ܶ��� w�
��	�I�I���z���d꺘�
}�_5�IZ�}��$�[��ݼ��gw"�nF�l哤�]�.�Z��I&�+�����V�mͻ�̝�X]o��it/8Ϸ���{�u�FFxW.��b�*�@��XZx������-6�_��|~�vr�F�J�#� `AgI�yRM��{i����=]���Gu�$���$�zk���L�5;r��ȱJ���b�$]�&꺿�ln�Z�o�9�rԺf2IIfM��K[�/��l��,��O^s��v&�֮˭�Ĺ6۾�R�����Q]*��Yȝ�v���Wr�2��j)\ �4���]ޥ�+��mg1���d�ߕe���t����z[�q�y&K�xL�����r�vJ��R �df:B����)b�V�N�{R��7~�:y|�u�-h���q{���n�dn$��*��pZ��_ݝ�ĒD��g3��1���=iMzq�a+n���M;��h�@$\��w{q�4�3�]�lU��P3;�K��w#�ڍ!e�=Ϻ=}+i���y��cV�g9\TGl�<n�"�G$n���ۑ7���e�Z�^�ufu ���P�]d&�m����p�4�����y[�7&�m��I�0��]��c���W�n�8���\3	K$�Ơ�/c�k�p��ֹ�FGv���Ӆ<l��׀���Wϓ�0�'h��PY�w�Dd�n��HtsN�g\]�_��ל:�����)�H����AyR�O7��j3,]�a�f�]`ӯ��ۺ"紱']�p��kk,��\k��x��mཬ]}��ǽ&�L���w�=����u[\��X����9�!з[Bz������+$S��z��R���dL2�f.��jrmR���8+��zN���:�Kq�hkMC�I>���5��{����ye��Z��p@��y
ua�FJ���z��	̥�b�P�w��:ט��ÚS��/n�7�����m�6ʤ��sY�;.m^�ـZ֒��|W
�v�d��+U��N:�8��B�s�8�NJP��(�瓔[�&#�^q<�Z�"jf�[jn�m,�J�+��k[c7 �/���`w�k1:Z���W�gZ�!ѽ��������a�)�#i�E�]�`��=�@��|��Nb����]37[][WI7y��ٜy���`�?�]]Ai�g����}oɤs^�m-I�ؑ=� )��t�To�Q�m����td|�&���fh��[�kP�[���ؕ�	
�������Hw�,r�	�{��)���]�Bt�n�)i哨$x�l��'�1M�m�R�<_#���]j|{�-0�M��5}uaH����zH�ը�ٚ�'�	�hε+��Zj��D���Z���̎-!ڵ&��8�Z3i��]�6O.wn�l�#*Y
��յĄ��|&�k	�RA�:G���䌛�r�샲�ȞF�Pa�v�^���Y��(q�\�����<��̬��-��Ɋ�b�R�3&��͛�hfvӝtKPKl���.�q�L:�f��s�]m�RɉN�u�C`)>̉���Hk���3w���I�^� X�FRt�����d_��a�Vcĉ�cf�&�5,�]����J
�7�r�V�-���C���g{��;j�+�Yiݍu�r�K��ځ���s�o��V�ZC�L�J�y�1�x�S�))�9>b�-*V��6��)�n,O�x���*�����f�m�@��T]V�Y,6w���f����\l�#}ø��� ���;�w;�{�a�����d������_u�k�7���*�VY;dN��9f8J��WVQ���؆
xVw:�uk٧D��U�,�WȘ	��N>�nʝV�E��Yv6y�w�!���U�H�Ta&���S��CRח�L�6��[b�y�����8�ż�J��r�PZ�lJ8������K�
�ї�iE���LC���|p��9:E��u����*) ��Z��ֈ1h'�a�RU8+����+h��-RƳ
�'k���mf�hx��[�,�wrL���l"��1R�};xc��}�L[�����u��k��>wX	!�f�:���8�vWSg7Yn��x����K��f-Ng:Ô��AA*��57��7�)�s�������/O,���kV`��
������N�w:2��SG ڑ�鍷y��
�+��[��-�ɻ�{�\5�/(j�]j�8,�b�}XYλ[ׁm�4[������7�tRXW�B=ƣML���Ǹa�gX�맥wns�G�n�.+mn /)��������ϷE�/�i�)�[Zb��M�B{���ǲ�Z�F)�I&][�R�X�ǯI3i#r��=.�+2�?`m�KE	�#�������[��+�{Y�M�*Q��}�L�����8��B��8j�>h�6w��o��/�nTڛ咲V���5e�ַ%=pε|�8N���[v)�wŤڦ�*ցw[ʜ�Oa����F�DV�*����},�#vf�������kX�0�_NB�Q1dI�u�:�h<T;5l I{�p��>�rXN>��^� ���7(���E��a������L(�z7s$Sgve���osY��S��L��m&������r�,QVR�c���Pd<�WE�ޙir�օ�Or��ǌ���nݔ��S���Xw����lpym�+8'A�-ɜmC��8�d �4+�ܕ�y��2{A�"��K�WSvtB޴����oR���v�O8
V�`tG3�}�����C#۾�I��ܽ��Z��_K��	-����Z�+K��-�X��5ޞ�������,�ݙ�d��7�<(����Hc����or�۽�g00��R_��d���۰�s�(e�a졦f�)����ه1�b�cV��`�ܢ��},[��u_u��^����l
�]Ȟ9o*���(u+C,w @�=f��&�1�4���p��8ݓs�1�w�6�^�yw�䳥��:��`�c�:��hvݬ��� �y�YӧVX��\�v�3U��W&����n�늯�&�^�����Ý63g^�غ��ӻ�3�q��i�ׯV7�1.��ow��ׅ`�.p�X��T)]$.t��Y�R�P�;Ut��+�&�#��v�VL�����+2R�ȵǸ�d�שfe�r��.Y�4��E��ٕ�7x��8�����[ q��݈Us�onIR��j)��d6��p��h��fըw|�P���⫴e��J]q���ps�#7��jݶs��Y�
��0�K���
��X��-��a+���V:;$6�V�)c]fgd����ܫ��wb��h`�}}�޶�r�IdV@�앶�b��q�`����ר�N���ip��̩�7nٖT�[�h�d�tբ���rʽ��˷/��fَ\]��yr���s��U�aBc�Nr�ovQ�V�V�ܛ-J�[]���_R6�r�7�G>mQ�ke^�X��� �`"��J�ꝛ
��Ѷ��s����z�2|Ȧ��8�ꜬeW@�,n���jgw!����{4������8[�v0���r�V���7�V��U� 
��� WM�r�%�h���Z37_<ˀ��Z:G�Xnb
����i�aX%�o���y��/�;���׈LȎ�΄�7)K8�I.�Q�5�u��L�*�l)(v���s:9�y+�`���k]N~��2�ڷ�eQ�2o��[�Z��=K]��L���\����e�Z5)
�W�������D�P�����r����ݧ�O� &�g[+u޵��yt�����ˤ�]s��y�E��îhݼ�oc�2�vޓ�H�!^�x�v��l��!ǹ=�K��3�:�u�4����g3�V��[����o@�v�ΰ!+I/.��d�n�Aǒ�CJ+x�<u��� u`�J��Qp#PW�@���U�f"���*�_@�l���� �Д��[2�;�\�+:��n�%zJt;#�B�'g/a�[{�KVE���Q)R���wv�0l8�� f��t��Wh����[<_\���c�}heL.ݫU;20��)��r�x̅h^Y}�Sw�\�K99��"5��>j�s��{���E�ڔY]�����`�6N%��Y�@" ��m&���v�PemLxxPcv&�I��C�[��y[��.�"�tn��[�zVu\��.����S/�[��ڡ�3*��I����h������6VӸ�5��6�-��k��;M�I�ʀ5wϬ���˹2����,B'����/L�(8*�8�:H�S����1n�* 6J�:F�������kg]�>�pWt��z����y#�`Y�upXiԩ]����-l�AX�H��1��x�'\op�uw{�[�� ��N:�uvW`���@�9���t�9��FB8��w�����ˡj��v��O0Õ��*���˼r,��g
��R�g5��\�*�@_5V�ΩN��R�B�7X�\;��e�,Xx$.�}����'�&�a���h�)�Ң없?Yݚ�u]�r�W�^�鴩�j�/��l��wlKۉQ�aU��+����씨hK��i�K]����ۀn��)3Y;,ǖT`:��!n���b����ݱk	gu�N;P��"�P��t:�+7�>�;xU�ާ���K�%L�;U�>�G��ٛ�U�41�
�d:9;1-#�I�;*�d���öҫu��bf��x܍Ƶ
�r5��f��4�ض��ʰv�/J����p8��|io=|$�����ޘ)��b��"�;���ݏkV�IԻ��6�$��z�$aN��ܑZ���0i��g*·I�ޠr�Վ�fv��ff�#�K,Rg�=�����XU��N�8z���wX�ٴ"K�p�>�w|.k�w����n�S�F�F��į�k�{���pN�UNѐ�t�YYEJ�n\^ח(a�'d@m�n������Ʊ.��Y8E��v��	t����|=(���aR>���H�]_L{�!�"�g�6\��I)�=K�㼾�n�SZ�w6Bz-���+:�ý���|�}�F�t�YN�i^=co����:u��&�w1VF��+��naw�\R��N��Ԏ��޵�
A�B�1���VIO3+�������['�N�B�Z�"reu�j\w�r�K��$Ss��;؋z�*��vyܲ��f�M�qY]n�*� ̺�L�
:t�G�����([�"�A�gVgX��2�V BəԻ���,M�
[���ї�A��cTD}�P˔뎽�p]0�1���g�u��:�Ŷm"�I�L�]���b1X�m�f��,���F]Ó*,�a�m$%��S����B�LAJ��5��s���]#�U�����g	�l��Q�K�e��5�5j���V�N@K83{k��wv���v.\a�C]nj�̼�R�l�G*[�T�zg���k3>����t�9�!�W��!��J�U����G������^Q��
�cg\��R����,Y�1��u�Ë"�L�� Kr`Mܕ�������ue�5y�>L�pn�����\6���qWj9N�³�nRJ��ڱ՛o��r��-z������ay�:}6T턛5+u)rwF���]B�y��<�JW���b6at��/�5ڍD�����ly�w��@�I H��
����������Οr?$%I$��,Ec�X���d��F��8I�u�i���5�9-�'��[�����r@q�=���՛#l�R�k��/�+�-��q�m�Ju���ۼJ�ܖ������!��\���;\9�m�go���)��c��L���hx�B�V�q�xb��㫙8�zHđ�-��s묳���or����w8�u'6�PV4��Mٙ���J]���L�n�i���6��cNp�-7��V� Z�44(,Z����)RX����q�d�黷s��Ҷ�**�e^`r�bYؗ����d"��5�}X�!���q����l�����c��t�Ξ�٨,ۍ�h�{5K�bk����a9֨e���FݤPk�T�������l�u�-Յe�d����}�$��d�
�l;�zȵ���Vn�KP}�W.�;9I�#��tC\x#�r����QRL��L%���̷��X�%���g5�U�P�KՅf�+�a������09n T����t9��xn��>�.�ZڟbS{�si\H�T.�<�.Q�>�O�*p�#��9Y$6>�9b�kLM
�n���еف���=�J�h�)�FM{J�<�ï���6X˻��+�J�����f�o��<<Pm�겺�#���9 %�hU��,��W��+M9��8,�k\U���w�:�x- -�;y��cՇ�B��->���'�UU{�U��}>����:	�x[kq�Ce���Ǖ��� otY�c{���q� �nm�Lo,փź+6Kx�<a#��̺1��-��FA�q��!��W����n$�V�Ŭ�zQ���ƜU�$��TE[��
�m{H�d�WvtyZ
m��{�n$m\"��-�V��Nq����f-
EW�<�*
�bY)cY6���ō҄�֥h�P˵0Ü��b����f�X���>TX:0	�e|n�V�Ĳ9D��%���VK�1b��ke�
�A����U��z�k/H�ɋ��n1�#�q	��˯XDx�
�)�dĂ �\���_Un� �`�2�Tڴ,���i�2��9<=̨�I՛����,_5�+��O#'p��aE���(X=%o%raOz��qޑNq�^e\Þ�C"T��W�+�XmWh��w3�s�nArP���i���^^[B�p�"�*�>˿Snv��Ww�Y��ģ �$AɦH	Q@FiIFAJ�T���Y�s�u������]6u��zoJJӁY����m5/V�����l6�@�4�@�M�xp��[�<}�`*�:�{���8�̐U��p�@ؠ١UK���	�
znQ':�{�5N��U���p����%wG�<0CgZ-p����K&�j���@��LD�K�HG�4q�n�N�HB/u^���q>�F:�7*�G�/��d�r�K#-ua0Ŋ�9G��oUP!�g*�Dc4j�-|c32�7=�����9��#� oV���6�C�W< `9TP���u)72���.�G
wIzCCݯ-]]�>�d�\IT��E��}r�K��( �T�U�t%��GUK2��8���
zĞ�K�~�!j"��,T{B퍁���k���G����z���I��������whwdLE��wS��B�-G��v\��e��O1A4�U^ZH��������y)��'�:�{D;�@q���F
�2H4���%J$XaU�#p�i4�5����A^�s���V��4 ����O��M�4J4�E�R��YA�컍֎��SWAn(�d.�nk�q����t0��u�l�}�亐BHXk8�0�Z ��!Հ�s���ٕ)��K��]{��ު�Q�<F�DNHߴ�C��4��i�ͭ�S^���ͬ�Т�8��+n4�ozJ|�Bh`�j����钢27� |>3�=�ha��y�O\����)v%�;F��t�A@uv�b'@oeԼ�M������`�>�O����@���̾����kr�En-��Ј��Ӏ��m%Ӓd"�={��-���m�"���S�˺c�V���ꯋu,�H{�ՃKOG�of쮈��5t��x3j���5j?:��� #r�Bѯ@v|H�t %�UC������˚[��ɦ.�d�N����9�VZ�Y�J�KR��K����G�����W�W�9�����(B��g`s�������"R�2�
�e���^�y�k��ǫ�����jgB�72<w0m�]L"f�<�i�5��W�U~���X��V��>�f�(�jQ����"s{e�Bp�
��`�d�	k��p�������~�~�G��~��G{<�߀���W^.��j
:�0�Nn:5��@��]4�E'�끉M ;;��$.�D��i}��}_� U�Y)�>�}�ޭ��>���[~�dB����D��t��+��&���<��M�e|mI=YHn'q�$| �C{�A���Flw��z�X0n{�KJ��i��i�5�c�DF��Ɏ_'�t�W����s��9�	Х�|A
H�0g������i���,�Oi���[ŧ�=�wm��K1UH���rx.��^���ˁ:�p��yny�����\^k_����� �;�"a#�7�n��r]��"U�Zb�%}x�Χr�̲-(�S�rU0
��!a�@ԑ�/B��a͘0
yÆͻrڦ� k��
��8�[0*N�Y$���'��n���'�X���G;�W U`���@��(>cH�������4W���,�����ޣ��ί,\<4�Ό =r��x��,�jYr,e��J��}��wQ���>�9���ي{@A�߈@ٓ��P�����,��q�����	���p���x�J����(�I�G��~����&�au�h`�z�2փ���}�S?y��L<Lm^&	��y"].h�,-T�R�q*PCp+uh~�[b�q΃��6�DǷ�z��g�Nw�-�e�������K����N���:v�Z[��d8 ��
qs�x	��g7"��6G > �>��>~��p�s����@]Ʋ��YB[9����Ɋ�~naX
�1$Mڽ�2�XJc���+�[S5�|>���>��k��sٖ��2ȑA�)���ITel��V%"��P�
���idDd��2��6�II`�p�9*��L�}�����6*�4���۫+%� k�����'-����h���s����e�"����uj
���9�8�S��R�4��GR�F��`��k:��i�e�j�m���2_`Z�d�NO�#�l�b52"�q VF�~����"4��^|t!E���z��b��1���*�TO@����
��/��q�06�݆e�hҾ�i�zL��۶f��*�����>�N�Z�N\q/EO1QQ�b�ۓMq�0�Z��7�� C�h�`n%Q��Mw/,ُ%�%�NE�\{'G��}��M��$i.�Δ�=��Vl�b����u��iVt꾣[���`�Pp�m���+ޠ�0�P����{����}�V����|[_G�ږ���M�KLj�<�]�VVdi���a�r�8�ʵt���y-�GS�<��P >w���b�n���mc���A�{���!bIF�'c�o��9�~�#���W�}Ԏ	���UF�����P7J�[ď]k"��!�ȹ���%X��]
u˛���2ś��
�v��7&/�x���8K��˜��M���l����<�Rb�����}��oc}����v"*ōz*,���͗��Y4:C
���h���:��z b͠ �;P��^L���}��G�}*��F��h@�Al޵]�p*����mƮ�-亖fM��@%��%�ّx���W��|  d,}�%͡�谿`�!/
�4�`�C�uL�;��p]7�z̞Z݆��{��e+&c�pmŻ��9�-X���ꪽ��W�}Un�Cp��!]�~�K�[[�f³L�V'D�yj�BΘl���+�.W�MR�LLa�t-D��{���/W���y/�Gp�j�Pp�*�ݢ�e^k���]�80E�Y2�
�	m ����8��`���{�-;�SR�F:�Y'6��{�^���T�n缪q�h��q�D�CH�>�j�
ʔd�&dQJʈ�($\�kh<̚��<��0���ȱ�oʮ���co����7.�\�;�k�t�Y��r���+�tB��.�ܳ*�I���y�R[D�2�D��A����l�Z �G��5b�UW�I�	���_z����+�!=�]xo�K���w���n��B��ǳd[�6-�B�
�D���U��~����}�}��
�cdnw
��I<ЬwŖ1Ww%M]M�G7��;.]+� }�)u�inP���K=��>"�WҘ�^���G�Q�52bF���]��F�])Y����P=�3��8�q�W8 �}�6��z�����c���^B3�}_WՎ ,V��6��<v�� �k��svK��ʃ厂]sOR���y��|ywWt�����ꪤ����#�.YU{��Ο|����!�s[9�v��ʆ!��5*fun�;�0Mh�"���0��+�9��u#�e�+'������	�<�3!I+"���VB�"�s��[�g/�=`)��"�t��K��"���s6ޙ_L�� /UdW�+������x^W�������-��<�F��5�ҍ?[Qh�ǌ#�I���d�]u۴��ې�[`�!}bN-�驊�0-f���x9�����B��%�B�����8����bY-�,S>�G��3�{�s�i�<i�]{�'�ʜ�����λ��jk�w�I$j���;����)��;+��H��rLsR�
P�Zw*�~"%1e��f^;��#ٖS�P��e@�p�z��}��3D[����]�]?����<̨�+�39������=�����!_\�Im�H��~XV�)��i�V�(�K��%�����a�t`C ��&a}��K��L��W�eK��ksLs��v�&t�fo���#De7�h�{�����m71�
�m��ˉ��Oa��F�K��3��i�Ԭ��d@	CG�@$���̮�6�V�*�"E&D��+��U�)�m�N��������9��q^��)�`+�Bf��4��В���h��/sLE��L� B���!�;���~ż� #��	�壼C�}U��|�ĲJ���h���t������y3�L�pÜ�8)�t�
���L�t.́�8x #�� _�O2�;���(dʭ,���ioV�>�gh�;����o�XI���(����j
�Bj;�Q���p�����ZL�����_���Q'�-��y��^Mz+1�&J̼
�UŕOs���Э0#����[c'cB�lJ����������_T�&k�z�@ْ��X3Y���.���C�
5�]!��3�us-MNRx��@�]ճe�� �v�'���l��ު��;���!���,�#�y�~�}�{��g<�w�.�n�!)���\=����&/<��⨆�j�%�$�h��a�VXc��G�k���J��8Y~����#����.�l��َ�SB���R�y:s�:��MʖF�b�f
E�t{��wt(���RU��b��@��}� ����$U�Nb���3h�O���)�/n}�uY��(P��� (9��6��)�]Ab�c�v�F�7���U���9�<�/�۽)�:�<�#�֬Nx�N�8k��wA��TS�f�̘��2�\8��2��U�#����#U
�Ɗ�g9�q�,�fXH�q�s���٢a�G2�%6����v���b���M��]��x0���$�ϑi�K���A�j����}�k5ۏ���&}�ѷ-y�LM��f�
�2���. �kM��Z2���f��D_�UA#��U浚�t�Z�(������ý�����A�.�s�̣�듉[E4rU�_+o.�����Q��u=���]挿a��! 8	 ��:>̌f�(0���KJ^���J�F�n�DY�L�7�U�����Y�)%�z�����Z��AD��B4�����o��ɉ���W)�4���\��:7-�v라���UPRt֍@X����޺##2�
t��NV��� �U
4% �8]��DcuJ������m�c�X5�"��@TDK�?wY��Ɯ����}
��u	�(�@����$��m�p�dܷ>y՚4�v��,��4o
�ݸ2�e����{�iʫ�|��~y@7����Ȑ%�[]1�G\UoKUV�f�$��#^}�	w��#�4�z��iͷ0�⻓��$LQ����`��=׈������.v��C_5\�at�J��1�r�Ҿ-O\�F,v��[m�c=�����̀��NP�!�py��Q�!Ye�*)WX�32�&fM����2Ξ��doG�c9�4n֛�MdIR���NG�_��W(��g��6iv�M�v8�麝.D���>�{���%>v�o:�i�V>�S���t�EqK��k��w��V�2��k�[�\Ⳑ⿸w���Q��1��*�Aɱi��]��(��!�9�����B$��wL�U�t��e����V�Yg� w��e��8����8�vXY�By�dx����;7�����:���ػA��u�a����/f���rQ��m�R'�j��T���L�q���b�+�0w�[��\���5�T���W6W`1�r��=�
��'N���ubX��
���F��2h��]�ke@�#�5rŨ	�yx�X�+��f7�&'T;�|&⦃F�N�κyyM76M��]�{���:�t&�w+a&���f��݋ZSn�I�#z�jzNXYXh�aе�faw��eDc�=�1tk�H�ve2�ů^T]�N�3r�э	G{��N�F������b�x���īb��߰;�Nk��M�]��7��7�Cg��o��$����A2q�.R׼��6�p�C�E����hPw�f4s��x��_��-�����L,,
�(�=�A�u�/b,�W,�q�vzFg�)���饖V�ir̽�^�+��_���ɴ��|����Ne��� T��13i�c
��d�J��W�-��»�4���Y����M&��~�� �?q���%VWr���gL�{�������ڬ�!�d�`bm?�B:!S�����a�kVBc���C�+�]���>a��ٶ1�����a����i�q�{�~�}��}���?3N����~�i�Au��I�h}���O̕'�F�(����z��PY?5��L�`bO%0��tϘW��q8�M?Io������~�����BM���?���11�3�8��*k�hO����څN$�5��g�/(�Y
�E�S���!���g�L�zʟڼB�`]����׾;�������C�1��&}f0��ߩ��+��e`�^�Ę�Y��i�4���!���a�N�����V~IS��T�F2��"��
�,AY$E�d�H�Q# Q�jm?���
�O$���<vUN�����c;�a��~���,�Ő?+6��`���1�(T�ϓ�t�_�([���m�I���Θ?4�T�L��a�+��	��� U����a۝�8Q����G�|�`��H��Y6�`[~CL����a\a���;lĬ�?� 	/���%�&&3���O�?�v��C��m���6��;��^}��{3���,���	�,>`(]Өu��!ܪ�O2W���aR�d�9�1Ę�񟘸��T��3��f�T3��P��v������~��{w���=f1I��V@��f}a\d�Y���?`T�W�@J��i���J��i��z�m+��L@�eOe�<�@į\LI�|ì��e~�`D����k�R��������c'�HT�v邟���+���?&�P���b��3�h����J|���1�/_!+1�z�?'y@Z������Lj��<���� ��b\i���������ٚ��[*���v�W@�f�5�+Y���Ś�M�*z�u]��b��6�V�x�R-+;���5*��)� ����O~�������r��a�*i&�k?��4��6�}�;�|�g�T�M�2/��{��4�����u?8�'�c1*e�ֿg���ￓH@�y�	Y��c6Ɍ>x�V|�P6�l�I�i'9d:�I��`q&�<��!Xc4�3�kn���}u��ߍ3��J�XVc
����V~@�LO�+*�v�}�a�*O%z�Y��~a�l3>Èm?2T���`)��'�i�����}�ݿw�gw��6���Y+�?&$��&�~��'\a�*m���|�g䕟��i5�:��p�C�����ٽc%a��wO�8�(��0�,�g���
R��s��BO�Vu�yh�&�}����jk2i��T߮$�+<����L?�+��~���2��+���t������Ry1/���i��r]���럷��]~>E��]��i�?̛Aj����PR��aR@�&�|�Èi
�2Wڠc?[�i�v�u�f;@�1&���u3���w_9,� �!���-/��F4�:LIP3�a�}q��1�
ԟ�t����f�T���!�?$�?��~IuO�Ri���1������vBM����ۻ��|i<�ix�0�+4o�_�H��Oɴ��d���A�]!�~Ld�k��m��1�f3��c4����J�l�}�Z�?3
s�#���p�6�ｽg��O��i�?&��̘��U�z��yY����a��3���/�N&8�[����lϩ�4Ͱ�3�?:AAO�0��� Q	w~��s]��?��! Χ|�fz��I�i�g��
��u��+H�����Y*q&}KG��9�E������{�>
��Hf2P0�����$�bK@*�0��Ɗ��· �HBDH�멈e�{��]��ֲ.�7�1�3��pTU͛���ʁtrY���s�/���a[}�U�=n�,�BR���b׵h�c���s���ɥ}��R��}}o��!��*z�+�G)_K�"���[2��U|�`P�o�l��$��&�f_���U�N��??>  >8F8v�_��Ɛ�}U{Y�^IW�n$����[\<v)�~1-I�]�V+���dN�����/��݇�f(6�Y�����PZ��zЯkÙO{]f��]Vfm���mM�kX��9�'�:����C?`b�҇#y�GΨt�F`HU���� 5_q�ܝd�����i��^H@9*�1�n�F��=P��&�!�j��!�UNY�VBv��j��UW����Y �NX�������8�pH���W6�`�*	s�hئ��;y.��9f��AтemFDD�j��!����F��/0�����98��&+$�,*2�D�_!_M��F�#�b1}IX�O�p�b�)�J%D9j��Pr��5Mt�D��kFJ���ܜ�	��Me]=����h�i�y��������5����"tsQ��XJ��R�>r���g�%�[�h,�}u�Y;��}����� �T���L9K8�H���E);5�e\5�\껹3`V�WP|�bv����G�j�Rr!%��~�"=tQ�N}��U���=�r��Co��k�Q���j��/7f;��N���</���^f
��^Kz5�U��kb#����{�ۖ���S��<|X�.͔*����U�`���Cà�K��I�x6[7%���h >��j=��u��L���c�Ѐ�	��)�c�v�����#ulKT6^�!H��ZS���bRoV�2ok�F+�����4H(e��[�+�`-%��j�� }�:�g
�#����B�U{�y0���2��h}~�ֲ��;�g$��Q)�t�O�чnJτV��AB7)�=�~��}���s�w��j�]V������-]�ﮮYz")YMj�u{�H�m��u|0,�{D�<�k��/��^Aܝ��	[�ai�G,S�U~����~g�
���C�R�4'��g������ͺ2��o{�������y޵�Oa�ڪ>¯���'�	�,��_}^���� 4j��x	���%��!�jv������|}���e��)#�mՆ,Tf�Y���N�<Of^�~��I	��	�qWR��Up���\6̸�]�T<WphK�z�т�A�edU��I{�'v��]�������Һ��p�"�˞��|>�׾N �ȋ���t3����D�"�p�v�Ѓ2&/�P)�L\��hkG3���O1wAC�Da%_TМ{P�,ɜ }l�g��s�u/�=��J�d}��2bWJ��s�1� ���LWų�n��8p�w�}KZ��������qN�w5��,��U`�,T*�0dAc���$Q��_Y����^��"��*�gY��q.��:�P�XE�1�JF1���HŐF�(�Y�PF(fS!*RF��a��$PW׵��}���x�7Uk貉�����P_k�C.��d�Vn�C17�7�孇d����K}����{b���m)��^tڳz<N�-�Txx`	�pC@âw��1#{������o+��OQ�Cg.��o%��Ž��A�`�v6���Z={�.y�^_����Y��������%Լ�|�`���W��AL
Vr�{��(����+�@�6 ��9q<�e�ڕ��#I^y����nIG,��p�PiJk��z�O���ޣ��u���X��l5}*��wa�������4��i�]����,Od[��r�uUz����)>�߬�^e�G���I���=x��6_޳�������g�`�Jγ�S�5E3y�S�
���L\#0^�� ��	�z����W����|+đf9woQ�w��S��TT�7�;1C�K��F�Yw�.���uKXbk!�Z�#��z��|���w��(J�ڊ���PE������p�~ɻ�"�w��Lޭ5wʬ%h�؍).�����xūe1lv�ɴZ�v�~4�.ƍ�A�0˷Q��ʵK��e&l��k��G�AÁD��}�Vj��7�v�pxjm�#�9M�BO�5�����U�(¡�����'m/������:����A�ɋĂy�_�ܦ<���_�����*u����yy��>�����/��0"��f�@o�����I*NC�����Ff�QG��s^CB�Y��i
c��:����mk/٬��x_|�1�8x9@ݚ��o�I���Yd�*2%ɧ=��̅!�5�H���>��~��4!�u�da�&o��^9��8}��S��ϧ�|4
eD�<	����=�]�Y���-b��MT���gX��eۤs����&����"�4 [���>�6��m��>��鳽�3낯L�+�� pD����i`S(\:7Wi�w:���!HAK�r�EP{[�
�w���Bx�.�6����(����:<���B E�\\���0�o[��7��tb)�=��b s�aE;��TkV�omE���y�{��M����_�q��������u�ڂ)h�g42:l�S�2�{��&�J�V��`��V�c�޶{3��^�O�����| |shx�̊��;O��9�i�8 D���L]Ӷw=g��q�gҦ�<��`�S0��o<��۾5ֳ��pr�U��πZsi�u(S��,�8��c��d�P�dn���&��1�xA��yI/��5HXP���R?d7U������7�t�mz���}V���Y��-��K<����!n-`�>Ǽ%+]B}'I���Y6�pʂ)I���XP�neC�w�����G�+���Ky���]����P"P�R�[��	e�6���w�AJ�W��9v)l���ʢ�λG�$�RE��)|~�ڨ7� �޽�Ä8����I �Q�@U* ��t�R������m�yr��D��3�����[w�S4c����p�v4���@�aڛ�����t�\�ЈgWP��/rRL�b�w�C��u��D�6���j�F�A�P`���t�6�U{ս�Rkd]�nk�O����������!�(t�!�q����`w��0ǘ6�{/�ú��U��=ˑZxpa��/}��|�UUn%+�*/)��9Z5�q�;N\_=x�5�F�&H�����e�Q�x�f�ÝޢF=�35b��y��^kLS�Dz| �}U���]F�ܙ�Kh���)���,5�mVQŀ��,}�ǽ`fb���%.Յn��+_Ը	���h�K�=��z���uU�z�uar��3a���&Ǹ.l��)���(T;��~>���HuM���Wu���� ���+7w�YV N�"�������!w��Y�jǃ�ʙei
��"��P+:��3L�Cg�#�d#�v%�������}3�u�(ҕ�K�K�IE
J2	R,X*��f$[`��d1�&�ꐰ�@dPajf��P0��T`�X�F����5i��&e)m&���GR33Bs��O��q�̌}Z�IX�4�9	�/r��VrY�-25� �Û1�Ke�{5,4&���ْ��Oev;�\ũ�Dv��z����S }�®��K�.4G�d*��Y�\�C��Wi0m:�or�o��)Gn/�	P�L�s\��_O��_}� r�$l�����)Grx�>�%�	<:��N��p�e%���n+��ȥx�*D1�����1	Q��d>�p���'��ǩ;���m{���|-mCzzV�{����Z&y.�2[�"A��uW���%��F;,\Zt�镇�i|��zl�R/�q#y%��I��bU�3v!�dg7ݾ���E���%�!�Ko�Y�Ԩ�J:>����]z�UT��'�r}�	�Idn���C	&Jckso:���L���=�x���V`�ޜ��,hQsp2;����nԄH��u{{�>��HEh�b����셹k�j1N�u�Ω��T����+R��i����8A�	[㎇�Gc�������U�b���2!��fS1C���̶4���y�Z/��=$������3�+HPb)��6}�pܴ.T,���ڸ9T��=�kMLߩ�+��ɯ6���B�^cJAf!�Ȓ��D�V���{{���sL�o*m]�Z���,X.�7Yql���GsP�w{�٭��§���kWH<��Z :���|2Ľʵ�(Iv�a��Q�1_�1���I�414�ֆ/,�j�i�{o����}�w�o�M���Dd��)�)m��Db��{��\��6P�:�:�������$+'�7Jö�r���d�vo��{ɭ��q7�ֳU�OS�3�o�IP��m%Q�b��H� \����7U�x�8�Aѫ��3�w{�'T�=����Ԙ�K}����mYH1�}�a���K��2h�w�Z֋ۻ�$��?��kR�iSU�:5���9ܩ��[��.��݁�v
^�뷣3Qcְ7N����(�
滴�N<��7�q�se����k���|�F�����^��0k���l�1�C�a1�@��بx�pG�6%v��w��љ�u�2�Ou�G�>q]I����Zͬ��(P�lX}�F��7�d^��D+���������9so���3���ä�R��n%����(�8�W��:or��C�}xM��j�l��*�6D��˪̼��=-+l������㳻��i��:�*ý�T���*V7c.��4v��ǳ/ �<^�h�uAG[x����nmm����;�)z`��t �>o(�)˻g%��[�M�L��m��WU7��7z�ݺ�5Z:�S˸2�s:,6T�u���oN%:��(��\�
eZ��Y���Q[ǽϜ�ݚ�0��(n�Ec��C�i��Oz#�jE���%�y:���S�T��}+�����x�.�7��c�[vA.��ԉ8�f|��,��U���0������퇵�d�*m���M���D�3P���[��i+n��*μW�r(m�'�q�* ��;9e�����U;���6�@z�:�u�r��XYɝڴ����sNvn���d�����t�Ӛ���ɰ�ǀ�$S���`���n٩l$it�s��fQ��Sc�nn�z�c���Z�Χ猼�U��;-����8ׄT�3[��q�F���-�"�r0��Ч�@9�=!�	@k]{4�y|��W�=h��t$p^��vpe���˚tB�cK>g<,űI��`
�wkA�S�ri�mBͺ��*������ן>�zL�%����`�s�	E^������݃��S ��*�4:���aʈ�2k �ܓfT<�H��q��|�7�]a���ݘZr��%�ޖՃ�6K6���p��L�<u���&2q�}C5\F�������m���X�����xq����UW��ڼ��_z��\��t��ӭY�S��J}�>���9�>uU�qW=��{�vJ[���z�վ�z�i�}j\~���N\x�y�-�F�ٺ�R>��o��V�3oi	\ �ex�`�(�-}�3Χ��A&�y�r
��c
�Yz�^���tx���Mu�O�wɶ�f*���z���N���7�F��߱�mr��Y.7��t��_9�I�l��.S;^�US�ު����ާ_	(��z��s�h�o�2_d��#��*G��jt�YX���Pv�jM�8����C�ҕ�o!)+kL:|f��#eb�!QF&��#PX�",r�*�0k"�:�GE��6�b�`���(�EX")5�a�EU�V�EVH����Eu5��i����a�E�[��f�
�#d��o�;�x����P�M��3�)��ua��x�רF�#�D��8��\�wYR��Uz����* ����o�����ZE5Z	��!�s�K#�Y�xi]��^�/��F�t�k�n������gf���rc��I�u���2]N�"8j�x��X�Dt/�������W��sh����s�F�m���(�����9R�r@�9�#(�R��������.����b����rN'�'��t���Δy�k�0"�'��U��X�0eAs<ս
fY���	 �"a �AV(]z��{L	�퍠4rj�$�{1l�����%��^H̬�e�TnG��rqe��8�<^��ު�\���:����Ԫl2LFuY�3e+� �tM��y�Ja�lX��E�~󽻻�����$##^�xp%bQ<Ȱ�T[*h�2V�o�ţ%ĝ9.�����]OK�{Fp���ܴj�]��KYaM�:�OvK��e��U�o~�{�g�ݒ>�����]_�&�a�1�������M�m͔��ג
�Uz�9�k���u�Uz���쪮�(��Z,`N�t�KP��l���'9��[�������#L���v~�> ot��7�t#{~�SX�=mk�u.ʽyIڹ�f"�w�VK�d
9_	9��=��>���UUU�W����T��[�{5�r���!���IgZ����S5���y襵6E�b[�0�_W�U�H�H����������$���{�sw������� z.l�Lv�L��z���H���������8炊{�f��瀭ջ�v,��cٓ�Q��e�Đ �)���\�
���hK�2�Ff��*�,4«���+XH��{jf�UN�կ�%���&����4f�n����Y}-Sᜎ���D9q�g�a4�L
j����PrI�.S�vkw�Ҏ�}�q�ѣ�ݷ�t��<߿��!A�ʸﮦ�w��PĦU�\��2�T.[����v����O~��o��� ܕ��a^���b>�m��߅��pRZ�����R�V\�.RL2�㽸�7�D*�>��};|�;}HGGxB��^�����|nJ�ى��jr1k��&��S!~]� �y�z��Ι<+NC{W������� w�}��,�5>ҵ���Qe#�T�1^�N̲5'v-3~�ߋ1�<n�����d�z�T�漼�M�b|A�bܱ\7�Cnw{�U��ғ��i0��YV{�{޳����_�s)�=���r�)l�j%�E�i)F,�I�"ԠT�j�ʉk)j��R%#,EU@eH�V
��і(%�,�����c,"֍��#F�-_!N��rK=CBY����ۈb���p�n+U���Ħ���0ه"��5䬥(����DG�^t'3{5��Ma[�kﾷX�[C[��f�]�E1�aǀ���2H��[��������z���|����c:�TՃ���N��H{� Y��j��"{�L�6q��G\7�&���w]+�U�_W�TD�3���]�7w̐�̝Ĩ׀�r��S�����_gr�$U����2����ޅ���e}L��u�P��z���kaq�S�=\���I.f$���UO}]��Ψ�����p=��t�mAh�Ur�5r�K�����+sa�K�ٌ�|z�̾�ԅ��������W���Z~\�V��$r�Q���m^vĻ*�1	(1{*�c�p�Y��+
��fd�^����oK�skqp�Mo����T�E}�;�ԗ�Z/0x^е�Uя�dղ+c��Ft�r�,j��v��7M�3��8�d��m3k���Ez���UyE|����=�=U�J���N��$�\�P�`4�$�ɼ45��̪��梳�N�;�#�n�'D'�ެ��ۮ�IN����33�oj��2�m�D�Pｯ��Os]��O���b�"+��r�}�3�N{����e�e*"�;��a8�Kk6��v��/�
d�����זQ�]>�W���V�>���UU{���q��e�p�	Wi*⶚فϞ�_:y�����=sN��Kؤ�*�z��W�|w��>]f<���x��<y�%ظ� �ZC��܆=�`���l�<�q`3�����Ի�uG>�}��\%߻���K�'�>��K��~���zƌ� ɐa�
���q	�%2�Sn�LYSY��˞��Ę˻�����kr�A�W1�TV.R�W2��|m���mZnطl�{�Z���ѵ'WR���^\W	5kn��A�>�}ݺ����ɭf�|(��d ��Y`,"�,@T?��'�e�h�_ :a�J�'5]{�Jo��o�hM�ơ��,W+���z��{��]�ot|�\p�{7�k�r�T���t�����a=O���n�*��}YW���/{�r+|���O���^�wU����|�TMo}5J#���\�
<�St�>C0��Ӧ�cj����U�^���W��T�Z�B{���.���CD3d�%�q�����(]��&���b]�W�:�e�'�0�CW����խ��0�ྈT�LZi���ʔ��L�j�g7q��nm3%�t�7��?@7��[N�c�V�ԿG�S�����\��fB �M�v6<u9ӰU�<�r�OM��u]U��;S���Wǥe�r�f�j��q-l����u�P��%��(=�w�0Č]i2�<�S`���=�V%�{ڡ�&���BK������T1()O���W�ޫ,�9sR�Z5m�劃���Vao_�o/�!�24e�_^%3�F�ܼۂQ�{�[��z�o��Ϻ���k��;��ql�����KgL�^o2i�U��*o���Z�A�x8��.�k�1�N#�q��:�S�Sqpc�ޙk��)����R����N��L�.ݗ�uܱ�Y�qmOt�p{ﾃL�<O9�uX�>��3�}��£Z�d�wed������Ffc��>���=�UW��o���J��B�nGٺ�Au)(<o�{Y�����9l+P���>��Nvn�L��L5�e��kz�+�Ftzl�<�H��������u�.���q�$�鱷��)�V+9e�M�2W^ݔr �cpλ���&�Z�Lkړ����_}C��Mvלnx����Vɭ��+��n�_�!;�JE2C&�6���� K�z�����WG�6ʽ�e����R��o!b�6�T��$�*���Sѫi@3#�����"I�&s���~~��EL�W#RG&��bQ��\W�q jɶ� sr���s�����UO{���|>R�~�.����J�5J��yBIq1EY���}r�5�̇n��y��TG�����yBG����6
dS��Lq��]ˀ1�d!��r�e�T\G"�I���b�s��/������C�����ZF��hX1���-l��)U�V��������ZR"1-��B�%�F5�`Y����4���Ϳϙ��4����=���rXG �
�9�[�k�EwX�"]��m��d��k!7�][Iڥ�f9��@-�-�n��T��"ժ.[��RQb$�"���Z�ZR�=w�`,U�b+X�_��^�tC��j+T���8����攧��k8�;�;�9Hc�4h4Lb���F�v���^�&�� ~�H;ռ�����P�.;(/y@�]�>s_<�.w8�r1o=�+`T�^�˞^���ŭ����
��y��ddy����h���༭��l��Z7h���^������}�� 	|f��<�hl{���Cn�ڈV[�X�n
rk�,쌹��x�5�t�ڄ�ݾ� ۻz�Đ~$�O���9��kѽ�Ϳo�R�L�zţngp*y��Y���p��+�kܾ	�Q��Uf�k�,�c,D���
�V �\ϫI
�W~�M9"�+
�Jҽ1�˝\Jo������"�4�?V^�[B�uQ�A?
K,��$�iŵ ¥}��6�����,���Uu+*���|*�[m����2E��w��m~VtT/2h]p�*(��G@XKJѩpE�����vj
lB��HǴ�5���շC��DUN� 
�]���խ����`]b��ѵxТA�����yxk'Z��{��$�I��D�딂Φ��>�}�vk��:Ƈ(Q`��W�sn��t�ʒ��w@�t0�R�-S��4���I ��֛T��ؘ��� �H&���3oa n�뫚����B�%F�{�9�Ag-  7)ߍ�v҇~g�q�Y9��mD;�9�!�`�f�n���c�ݚ�n���杔�m_��*�  �AQ_�x�n�J=�D�B�op�[ lٚ�_ٗ�ch�����s"�)և2�Gġ�UT��-���<N$뛫(����Y���Z82�ue�a=m��5n��swpQUW�	��Gz�QE��Қ�{�»�˾�Zy��8���B�wr/����Lα�(.�������:�2��9�kOj��^X��-hxq�;�_(�wOɐ����N���c�n3ʑ��V�wץ��[}\A�@����O.0�t�j�zq-��Q��ۭɪ[!z& ��\��@Q��gGf��j�e��+�\���hѹpϧj��,b��V㗊j�t�e�i���^��A��h��o�, �^�3-rS��k�q6c-��9Xּ�@a�6k�����Gq�X:t�(iʆv�:�4%SF���8�Bڽg�3Ͱ
���yc�x���`{(�*Ѱ�{ch;�}6z](���$�љ��]�0\��U��)W��Ts���U��a��>��Җ��J.]����,�yejW"�TaՎ��X���'ܨ.�ł�1D�]�x�LY*YɈm<n�d7�3,q�����(����얣+M:�n��Yʝ]p��w�Q�Q���,�	�$x��|h���@c��|g&����k�k�o1J�MIγ��op�m�ri�к=/�Q}�c�|۾��z��` �,t���Y��6��pf8y�b����n�?[�\������r��7��=�%���q^L�"$_\yGt���!��x�[���G͜2�tG��\Ǘ�����J�XΆ��q�T6���v�u��*��)�R<j�w����pե�1}34b�*��P�|V���q����d
Puh�y�w|��ӳ�H�J�����һ�Gt<k�d��r���D��L��R�Z͑��8�)s��5�z���}���߿N�� ���ޯUZ�;D�P���ƻ��X�Qh�T{����NAם-���0q��.�P�9[�G�t\G�bx���v�͗*p�J��U�p��o���w~��M}[�&�*J�){���4�Ͳ�t�^���T�u>}�[���SP`�'FR/�I|!`w9�W�*ǒO��ݩK�ҲT��1����������q��������r��PJ��TC�#�e�2�Mśe�����)^�W�����6���o�}9�X�m���?}����w��j�T���T#[���Ă��(^�J(e9�ق[�a�v�eud�x��p�;���_b}()���;lh;�޺y앗bۇjXegIplS�8���G&m�kq!����jV��%�T����[��'��1��z���.��nQ�ܶ��q��n�$�ܧ:9�K'9��vs��\�j��O��X>��z��y��c4m�Rh�|̀��;:����0�ܮ�;��{�>�uJȦPs`��7��G�G�}����'�Q�o�yf��1��Nj�ԏB��w�E{m8��5njr@�a��W�~�����݀��?J�Ӝ�V4c�=G�ث.���Ͳw)@��Gۮ>�����r�/n��^ur�va��f���;+��M��dIZ���Q)��{�[~�}�{�5��� ~@A�@F��o��o��c�}ki"����������oշ����כ��@�I�IB���|�B�f�¹��k4eEY�|l3��
�MBT����9W.�����*YG]&��6GEr������g%ݩ��^��U��-J�iK#�Gm������վ�,��|-���'lNl�Ʌ/&�9�XQv�Lb��9�9%��@%�Q�^N��Uz���$'��er���䡓�sq�s;�:�R]��+%
�sy��r�.#�v������Ŕ�i�j�>���I�����lum1I��ȸ�.dJ�NG��^�z����lύϝW��.�l�Y�Ⱥm1M75N6R�͹�e���/��=5�K��"t�;/VF0 "��1�~�>{�9�F�Ғg#��S�� 5ٱ�.nh�Ζ��;��*��~WWB�I"�"�GT�K!Ykd*��`i5¹������_\���\�fTX{)-�p㬮���,ހ��W3����u2����F�%�ru���8)oE�i<�����}�::Ky��S�^z_�;t���A��K;%����9����p�s��m΋{bUŪ/T����O7�����¾��7�E9ݾ�k��H��b�U�Os�w-�RVd7�&]mf�6�Sn3@
��^�P����2���FZ�M�H�9U�l�+�)�$�3���Klδd��Υ����b�z{�G�>��9�j���=$���Z ���vk��v^_c��y���b'Y��C�Ԅ͐�G�	 
�0c�{�3��Q�N��k��h�B�1�Q�/��A%�s<��4� U�͒s+RG���,q">ǚz%���k�{������G͕10�.8�P�
Z2S
�U�b�̥�`
70�Bc(�F����d)s�-�@�FM?�**�L�S{�6�׫sH�6���}���-�q�N�z��l���/�m��4�A�H�y��O���s���gg\��>�<�u�AV�W��Y��9;P�dԝ�3;=�{��^u�{V	+۵=� uy�Țx���gS��lҝS�����V�ˉ��1
g��ޜ�#*K0����z��v�;B}.��L��|��<b��V����Rt��!�6[�v5�&G$�=b�C���}�v@�J^�t,8V�F��	�PB��)�]s��ɃꪗY��%]!,\�fP=`ƾ�x+��E���,O텊`�Α`J2���nvh�lJH뒷S.l�}��@&�`[������=�UO���5��ǭ|��s�/y��L�r�¹�8(0�c�ol�y��5�R:������IJ���c����B1�
" �ŀ��z4.�u���9���y�S���wbĽz�q�Z׷@�i>�T<l�se������[kg_1���w}���d=��5o"NtI:&tI�u�f�h����y0�9
��/F12��*�O�ՠ"�3%d��̽r^�L�o�z�����Q���C���!�j<#2�ٍݥw�L9&9�Ɇ�w�^�Uo�N��v�r���ު�>בgۦJ�m�ѳ!�rb��8���`�=�.���Et��#KU}���|��h߹|v#��_��W�{�l��,���_tǞ�������>�A����2[9m\�:�Q�M�qu.�WNa[=�;��������v��{���eǸ7nP�w�u$�p�޷	»Rp���W�UR�J/��z��t��4��£n��F�l�{I�>�k(@4hB�V�,�z3XѬ�1�xd:��pcCLiv��M'��HDF�N��6�,{ы2A�3�vE\�n�mы�^�4�a}���u���}]�r�1������}�=�N���¯����eV�C$��Q1*�i�:���k�ӆ��[^����0�2�/3T�9���}UU����P�ያ۾˿(��HJ��5��/�`G&4���ݻ{�D�^�u9j�1eDD�z#藉3͇~��t���4�i���DT}���r�=Y30HJm-�P����e�<��}M��=s՚��7��;��APs���P�̡Rs1���59��a�_�U��ꪧ7�뙳��^�QSD*Q׶8=%!�T�^'�#��=-=�u�q��J�)S���^�>�RN���k��y���5 ��A��*w�ېXxDb�y$u`f��|�	�|����6���ss�[�Pz�+f�;�4T�T�V-�m�����L�0)�7Y�}��H��T�MVb��4���[`�j�r�@�I����U)�eA>Ve�7��%�lTRw<�gWb�Үl��94G��D=&z~(H�,�ax���_��{�Y�v�y�8^aw��{9�q��q8�f��s��P��q`�A}�R��U�z�u��Uq|�&�5,<����5�����r����L�\b��VNepY�,ڭI��1�H�bڳ���ޯW��g*hd|&n	["ɻ���S�wT�md�@���J��;�;������t4�T�U���% "b�V��'1�����n!̮��e1|�EBW�7ώ�X���)r��ZUTE�f\��\�I1,RE�ILQV�Z0�-PUKL���~����Yf��IJI��:�8��c9b��{X�j�;��g�P/�ri��^�Pevn�4V<��Z����JԗK�M��D]��������`y�*�����L:lcٴ����-56�P�)oJMUp�]u�)�+K��DA�|; �cݛ��ED�A�O;7T}o[9��lX;�J�W�`�h��i����*,�OI3:�s8�z	�H�m;�Dh��G&^������{]��w������D,���.�U�q�O��ކ0�}7L.XW.���EĻ� �+���T�}Tb�)��=ޯp�!K�97O^}{-��κ!{������B���B� t��k�֡������i���8VV�3���}] �4c҈��~�3�i�C�Tro��SR��w'8��ۡcc>�z!0���\\J? 7�}���T:c������G�i�p�t�i�ݖ�Iɱp��x�{%�w(񯐮VE�l�F$�L��W��w��%�� �"�j�=��T�!%���$J�kkl��
C6$��I^7-Q��A�90,�}�U�jb:{E��ĂU�̘����~M���W����h�~;�����s^~�f�	�2� ���|>S߭8�j~-�}��P�)c1v���M1|��Qä�p>��v�LeV�ɝn�e_>{]jj�SڊV�lkc'g ����}�!~�&_�� ����I\�!S���L�����%��Ø�3wn�r���iE�@x���$�N�ᝄv��R̌�x�茟�����׾���u�����A�&��sy���r��p��P����5�2[G��0�hĚ݆��jk3���t��}8���"u���_:�{,��W-���]�5�4y���h|\ɞڇ�4E^q�e�,ף�v""��@��s��v���N@gj�4z�:vhBROaTz_��=*�o�'.�徙�St�X��62cX�4���W[LO�)Q�L�_��}���5�C6�+�"ç��er<1��u�}�Q"��xaF���k��C��d4|lP!�{x+#`� �	����wX��*�;*�I]5���׹�|d�̚�(��@��K�~M:�3�e��E�[�p-.	D��^�ת�K��uN�U�¡r�e��,Q�bDC�Zs��h�R�yܚn���V�᫗�κ��4�J������d^�/�R퟈7Z�Y�)P�Ǐ3	(~�3���}�]�*�^�B�1�}��iUR/>���h�k,�(�Ac�U��k{�P̀��k�c�\
�5��l]�	0�0K����n*H+"�a�F�bg�vR�-
��wF�r��"�G]�pi��v�������5�1R��Ɏ���wg��0�k�6�]K��j��1�9�?co�t��B��{�`��/(2���j����z��Q#�̙��������m7�53��o�}�{�듷{[�XdTC5AB�:���̼.�3�9}������L!�T.���gQۮ�1K��};�P�� f��jv�B�;��i��O��mu�Y�GZUZhZ��"���D���:�wv7A��W'���[����+���}6(�K��ĪK��v��kB�V}8m@y�]*ɗF+�[[@�+�8j\wxu.�ݮ��m��n����p�Q�u�p�F��m&Oue�1wӅ�+0(m��j ��YOo�����h0h/�;��7��xZ��k�qf�\�v:F��k
ȍq�V��&�{�PB�[�0��U�0�3��7.������)�.4S0��!N��!g��'թlL7����Esj[ �wX3 �^./A��j�ڗ��TZqel�n��=�iWI`�
�b+�6��m��oKaݤ^�#5u�VhH�,�yх���N`���!u޲]��"ȣ�oh�ux�F����K�g6&e�K5�I5޻��l��G���(.Zn�i�wOtH.�p���cF�K�j�L㶝()K�k��{a١�_e͜�Y�[���jS���@#�GR��q��c5����I"m_��+�<Ǌ�m�e� ���,�ڙ���rlv�Ӓ��eT�+������&�YV9�N�&�I)Wzo�k�w E9ƎS���e�u�	��kbhy$��mӣyveT��t��,=5�^�η/4�;�W�i�H�X	יrcsEgg>��"����|��_t�Hœ>�i��l�۩i�&5gz�{�Τ{ZtZ�ǠׁW�XX�|
47���:5ˉ���e铟MR���*�������vt�f��|�	���c&�M����v�9�����sHTH���g�\U�X��c�Uj��5�\�!�X���f�B?t��G���tcנG�x��p����9%�Ħ���"��6x��G����}c�^��3�dȵ�S-�l���{4��1�̄�.��h�pk���Μ�}A�3`Ff����}�~��u�3=� ��|�|s+���G�����A-v{i��������N��$t6*���e��ќ^��vV���p�ː�������F6�\ߟK:���Y�8jta�NXD8ђEm쀝n����.v�ʔ��e��w�H�8�ꦾ�g�G��cL��G��gi��7��nܗdh��]BzCО]B=�R������.K�Q9px���;����|߯���́���3}3LLLL|`��||��g+���1v{�ا�P,ԡ�T�9Z�Sz�=�=D���|���W_ﾤ���?�/���w����S���[#��@�z�Q�j�7K�̵Ĺ˱;���T%],C��b����`65��+.�Zں�eƓ�5Ǔ#�j��y��u
|*��m�����LE�ĉ��YĲTd�s<���7{3t�D�+�h���#����pT%0� �#��'5���C�G�}6'跆|}'��>N�L��1�4vxM��@�	c΂9���H 0��X�F��%<�3�^�c�}�(�� �^�U3�|4��1'���"a�≺���l��kN��13P��۸�%&',<�(k�<��%v��������2���ut������-�Q]�,A���	���[��,�9o�1.m3�\t���aL�tNa`(\Tꫩ����1�`G�?�;�]��9:^�=�������,�y�UA���Bgy�����!S�Q\]d�}���w[y�����G1��0y��[���̈́z}�D�WU?�Z��]� )LIRV�+h`���aLY�>�����s��6�]u��m��xR	ER�
�P�H�S����5��	P(0��*vL���ȸ$�*d���ܳ��)b�]�]/ph�Ԣc�P�����q����F�[xj���%���FUG�}G7���z�Х;�:����9<gH)�)��Jcr���K�A�����T�Z��p��km����fwU�`]�ҤM��n�����Kَ�L�ߩO�#:��Y��(�N�Σ�9����[6��X5����(��&x�-FzӒ����9�:-�Uԧ�kI��J�}��/F�K#�":�Lϻ���.�������n1UM�Ж�ae�κ�_H��j�`BAߢ>��ڤ��A77d��Zhv�z~�g虑�(A`1��������z9�����"���Z.�z&�R��+N�RS�sJ m뙞E�
.��e�L��x2ZOhpڱ�iN\��������Ͼ��Dσ����bg���˳�����vBmڊ9е�y)��ZN���s�ĵ<��O�ɍ�O��5ֹ����wJ'츂���E �D �$�1VAP��f��_��U��gtvj_Y�i�Cp1Y�wEIÔ��z�V�1���O�|��o�cj�TĬ^��D�5ᐗq6��t���q<�=���r�y�l�)z8��GR�ޣy��q�d�ʗ|wMF��3��s_HlZ �^����L���1�}���x�l��!����zwx�͑�zꔤ����f%Stj>���lf��y���p��Q����DC������k�;�m7���� �ؖ����!Iw.pYTxte�\f���w��G�=�����9��f6sU���w��g����:m��o$	�`�o��}2��W,��/'p��v�����ɞ���/N����]�b.0M	�����U?�E�g�#��Z�{G5=7kqܩn�.���7��Y8�2Jǳ��z�����]��\J�fbm�L�V[������G���ofR��,\G�R�=O�~�M�	�,�J��Q��j4�39]K��[���{
�����5�)|���c	�
 �˳	S X�	�%�ݎ\=@�=�n�b��f:ɽr�u��/��-����r�,�;��Z�q���B�d�yt{���n�U�:�'T��S��T���ݿ}�?[p�~~�־�H+E���|�M�N6D�C��WKb�V.q���Fn@��e�F���Ѥ�4Ŭ,�wsbc�͘�{!\�q%��{���DzL=�Lz(� t꩙R��O3hj��v��������l��oR���qy��/N��w�	?�d�:��?se߿A`, P��Y�j� j��z�:ؖ�`l�:5j@P�ulϛ�'yL(0�X�Гب��>}]3�itD|����;D��>���?��Y����E�4����Z��dA��1s�A0���4�y�G ޺��]FmO��~���A����0V3s��׾έe��U��#�;��M>&v�uM�\z�_2�,��*�C�N�eY78�ڮL�}��hΰ'ɞ׳}����k�ٟz�1�m��(J��B�P�������������i��lA(퀓�٪���^���gG3�*B��˚-%x�-�_h{��@_IG�\����K�ԙI�zc�QP�OsrP�}ݎwr�%�2��R�ZX��7�n�!�}�f>�n���H7)%~��G�U/]�K᝾��y��Q%�L6���V9oڔ���%xpu!w�	����Bg��&/�b�+2�������������s>Ƨv*�F���vN`KL�a�T���1-��I�:��v���ƥ���:q#z/�K�e�44�w�*����w���?�j ������fZ8�lq�ҶE�����'b�'_Տ�OՓ3��Wj�]���P�Ͼ��G���/�,l����s=/����H󩘑M�N�횡��+�9�#���=51�q�����Q����ѧ��}#�����*7�&��ڄ�B��vF����O+�=J�rt 䙙֠sȔ�@�1ܜ��;^s_k^�k�Ts��ijX�����������Dƌ�l@A�כ#�*˲|9��CR�����nUݬ�%�"���""�DJ��Va7
�gF[;�/B��WE��,�pU�]P�&����}�Y���Þ�72�ҤD��;EK�f��-��t�
�'7�K���ӌ�(�(���q�X30�[��묧�~'�"�"�Po����rS}�V��ؒ���n�ν��n�jW7@�+5S���L��S�f�s��V�kM3b��OMn�;��̤���������4
�+�u��d��G֪q�村у���[$�]��Y�
��;-��R!�5�ۨ��W��4~�CG��.�v^P���0�}�⾀�����a��xև3�l�B��9|��b��ݘ~ۭ#�^��^65a��5��]J-u31���E;i̧�gzf�9�
^�.O�A?v^���P2��T�/:�J<r��<�|픲����36��I��
�Q�|�๊����꪿�U�k��A_zP��B4O���4�3s�뜋Z㘨�(��χ�����~�,�@�w
1�c�ڼEr\k{	UƵ֡Ο��,�6����]�<�uČ�R�S��13�A�R�c3z ��0�u���y�'k�g�R�A�]+B�1�Q�1���p�>9�{�
��k�[V�z*F�< b�����T��t�� �6M.�:���}����^��.N+���֏��4r��ϣ�T�/�0��qY�	��־��v�c"����Z͌�[�Hb@��d;,�bfg>�=e���u�P�RZ鈈�櫽�,gyb��؏1L�r3;D�r�Ɛ�|�P�Y�nk&wAsb˭�>�|!�g�XyK"����Q��>��u���z2(/�G�G��z���6�T,]Jq.�+��	�QżH�4�ݻ�����#ǩ��f�9ḩ���`�5Sk�T(��V!�����o��oy���j���,��WmV�Tzya�e=�*m�
��
�f����|��P�v66�:�>���+�S3^C���<wF�L���'�&~��E!�#�dXB $ �� ��� �"0PD �b1@PdD$d�Q$a ��-�����:�0;�Ә�r��HCqJ�Z�=��3���v���1�ᏻ��:p;�4}�{�*���hA7�mm�sGS�;r������R�Bq٧a���M�L�b}�W:mC���|�>�ŭ���<�d�-2��磟�4K��_x��}b��7��c�N��F�p�3_���7) 6�  }��Y���3���7=���e&�]37�������>�!�S��*%��yr"r�8���T%�����w��)KF�M�t�!�cK�ꠄ���LK"ۺ�}��^�菣�Y�o�_���[I�x��Nl
�D F��iq1j0Ӣ�+G��	�u
�c,9\5�Q&a�~��q��������|}URLy�\'7�h*n�Hn��*�����=[�
�P;n��O;�z����3�P�-��~�[��V�]�c`p�8�۵+V�d ��4TR���>�ǖ��X��\�m�=�g߻���s�'���Lʬ�h"KA^�<4}�V��h}ư+`rI��>ILg,Յ��0M��} 4��o#bӎ���QSo%T�#�+i<��'p�(���m�)Uz�!1*}�:n8�
B-���3���z�jӤlR�[<٧����g�q'D�5wp�*��5t��֢�W�}���zZ���߾��^h���&���hk�3����}G��Ry@fM���̙��^�!�ΫE�(�B����"=����%��e���\�7�S6 �W��zM�r*T��h�L��f�=5:��g�)u6�
:b�bU�H@-6��Ŀ���Z!�0�oﾏ��q}�n��|�ۆ1H��?����`�_������ِ�5n#�!fR��mFXW��˴}�HE	Qz�i^x����^_������KG3Y��s���J�8��Xl,B���uc��Mc�j8�.(��t���\���9�}�����
�屗J�i���y�*� l�r�G�O�X�I�g����F2�4	|�����$�
@�@�U�>�i!1_����9�����w�.5�q�y�����K޼���!��  *%����
��1+�ǘx:\� ���kt%��Q\ma��u@��o��]VdU��i招ͺ18|qB"w�{���h��|m��R��U�M%����Dr�,����J[[a+* �>�򚨆�eı���h^�cv�ǥK�h�~ݙ���� ���9Np�g�0k���Ì�+�$��UsѕF�aTD"�ņg.}�k�$炙�q"p"%����ԫ��``8�l�F i�S�5Mr�<�.g5s5��ц�5�Ȋ��a�j�1^o��T�W]�Q�P^�^腙h�\��ˣC�s(�;�֦(����iʛ����m��&6RE�Y������iʜ����u�+�iϳ9t�3�����{32�����ʀ0k2ϺX�1�2��uV�*6�Si�d{f���!U`$3o�`[��]hq�w0߮���mRT򻆟T��}�{}ޡ��7J������m��B�����w�rn��®a�K$��� ��;J�F�����;I>�=�b�#yv��f�X�k]��ꠏ�S���n-Ü�(R[�rn��� �o��M��t��<5���̴���YÔ���;.dkTi�N�jZ���]���_�eG�ł�N!���l졽q�P��v���l�LHql'_>�gH��i��i%W^s�;k�����v���n��ic���[r�b-�{(9���i���3@����-��m����:a&�q!�s(N�ޝՀVæ��s�ݐ����͹a�;�<	Զ5e"�q��E�Y���}\�V+��fj<b�}Q�����ڳS4�E�l.= ܬ�AM�|M��sP!�P��N^8�	i��v(��zf8KN��"�y���4���"�t����t��*�$Z�MNs]+-�m%T�U�RΖs^!�E���9�K���c��6�؜�\֚kD���fы�t���!F�����W(Eeg+/Zw�sďr
������P�/:��0�ݠ��hJ�ޘ:9;oT��Z`�ɎQ�u�4`�ТN]��X��YB���^y=;M1/�:l�w�mh�Y��Y�8�f��AG%5�a�4���ʕx���#X�!:ٳH0Vimv����>������&DsFٲɴEv�r5�s��IM�]�t�0��;@+�PdC'|{�1mm*d'��M\��chk=}7�XC�;>�`8Y7�6��(w�,��ɲWr���S��+
9"�haۭ�Y;x���r�L�4"_��@����0;�J���!���.J���j���T1��������Y@d�ˎQ�� ��A<y�H�����.�!�}��=Ͼȩ��YB�b��ˮ*Ȗ6e�3-�C<ΥW��f��*+��3z�ȸh��a�q����ܓ1:�Tİ˚�%��w^�|E?+������U��Ke��­�|o��Im�N��k���v]�w��W�.8v?��n`�]��s`r03菸���R���p�c]�NʮCfA��1��Z!�Y�M�:0C<�<3Ó�Ԑ:Gyk�o=�9��H)[7''y]���\{��v5Pޓ�ˌ�܈���N�&M�[��+�:��x"�/FPX�5;;�US����U,��S�؊����>��g�s�9;22��*|���uEӺ�}��E�H>��[yw7����	�y���[Y��`C�+s>#��o�U�%��~���l}�(��`\j��� H ��P~'�.�Y�%��(�V��wҳS��/q�Һ���v3W�:}�\Jq���2���Fe5�r,�-� ͞y(��d�����؝�$o(�e��uY���Hn��K�o$Gɚ�]�e�S�S�YAVC�L��~&�xz:,�19}���Wn���ɚ���.���Ty[)��
YB�gR�W37�Yb�W4��*sxލŔtV�,�=ϳTc��p�g�J�T��^���8^��~��g��oA���H�Ő��s��-�� ��	���<f4�>�������~>غ]=oS���q���W߇�}_�Uw�����f��LL��3�t��{�h���r�h��:���v=�*� ���cV�b�z=������wk����;ԭL��3+��8�S��-�D�D���	��ۣ/��3�1'-�.qZ��o�t�����0�t�j�ܟ}����W����u9D��Ϣ>��}�O�%��B�3R��jB�mR��kfK"z��7�3������TV8��`Ɍ(� �e2�*�Ž��߷����/)�Py,��Ɏ>l�;N� 		f*��|��|2����M5[\ėzt�#]>�tNC\n9o\�q�-�5�d������S��CT�iu9�ʠ�ζ�T'�Y�K�
�(��Ѡ�H���#1�c��\#Ǚck5P}��rZ�>���k*����\Twm�kw,Й���>������Ne�~��L�9Egg�����2�.N&զ�w\.J���!�DN:&nZ&�B,��s�x�1ﾊ�}�α�YM�x����;7�N82^��S
m����88QKj�u���X%�.�@�eܥc��\�9)2j����}�}��|��d�ʛ�7��%��P�w��Բ���)��;@F��T�r�F�h=H�M�m�Jٵ`�2%�2�q��ﾈ��z.��L��"� Mi�H�<��ܝ��e��X41��dg�F��\�@Kc7/ᐹ_Q�x*ܸv�uW����8Z�G�9�^/�k��fs���y"0H,�T-al�P�)Z#�bc�)b�0�A�A�0L��B�4���ʖ��VH���ꕰ���ϵ�7VV���L�쭻����r�5��3BÖ譧a9�x��x����3u����V;��2��@���[�e��N�.Kq*U\6ݐWI��5��eC{6���| wjV߫ޅ��Q2���>�:��g���I�NKX�s3a���q����Ë��1+��|ݻ�.���=��=������W�B��dA0��������Daᅊ'J��=Uռ�1�b�R}P�:�j�]����1n�"x �7=X�D�}�xex�u�K��`��B[ԫ��]�Tw��62g���6I<D���E�릘ll�}�'��j*)��YS�7$���&'z�;9D�>3xatx�e@\�A�:�t[�����lRQ�!{��G+���ʣ���M���uE@Q��F��7���1�~�c�u�13.�-:��ԍ9ٸ�|؛�E���ڀSBL�;j����S<K�I������4J@kA�b�Y�A�Y,�$SU��3-BS�)j�,��~
�Fq{�I}�"��%ֱS�#�:Hr,wrf�H$���u�m��YKC�q���@9��lBpk�/��7�[46
��,���Ŋ]�@�����ّ��-�ŹG��h���jÓ��0#������O֏��]M�>�q����Z��1���a�4[ѵ�oEʲr�ђk+��%Bzܾ|��U@	��!l�s��S�TsP׾���4S�7����g苕��'KR�f�Q�&oIE#NK���yop�:���K1���|8��]����%e��3�G�����3J������[ףW���D�pv,�.]�Eџp#I�Ѹ���Ps<}e&��o�O��vm�i��^������A���F"\�	O&�e2�:2T�<�Z���y5��E��������-�7`k��8�&fwt���؈-_���/Q�k�Y�J;�.�dO0�9|����/�;%������>�h�@~II$ ~%H'�3ַ}|�����d˅���X/|jn��\$���m5����n�זv{t.�#�`��Pѽ��Ք�:,�He��i�6��;�77H��|���Fi-��rۿ��1�G�o<��ħ�;L�~���NvN"�
7��tTͥ[�POMn�+�ݹ��e��L�u�3��x��\��ʼ&Ob�9/��ﾏ�31���\릕;��Za��}���Ռ�|�3���p�6���v��d�gyƅ�4f���%i�'���s:B�^�ٙ��
�����Ҽ��P��ע%��*�����S+�_	#�=��0'&�AN1���U�!fIT2}���l��eQ��b1�(˙�e��ŧ5�T��'��
o��Ө��r�w�u�lx�cp5H�Y0�) �Q�}j?}K�˟Mv��}�=�.��޶5��eK�.��4�2xYUM�����&4�n�>�j{_kB�ɡǊ�������+P�_J�?7�/�~Q2L��_O� 
GT��HJ�$d�"�,��
�(��XLњX=��d��b��5�q>Pg��ݽwZ��V��vr>�5B�,J�*��|"��m��^o�G��xt��p���Vz�5�kˉ��#������r|�BPz���T@��`�U�J+T���\+wa�*�N���]=�N�x��8zg�����wr���q��_����������9=��2wh�Ȧj�Հ�e{ǈ������r�+�=U���Ƞ�74�/k�s�Z�=(�X�V&�g �x'e�'N�3I�bgd9Q�r�\�]Ԝ���)��3���O��?D}%z�z��Zfhu	�杒���*^��:8�
��ni�Y���o\���I����.B��y��b*�O$f~��ġ�u�]9�ՠ�k{W!^�-�U�&LK�n�����NJ�º	��O/iG=�8�t.�۫�-s�~�D���}11�|��`���/�W��9�H\%W�\(5iّʩL�f�����I]i�mR�S�*nr�830�.Z!&	+��J̌de`�9��+I-�b#*��(W��'V0}�m��K/�����
�QK�a��W�.�����S=�%�Gv $����to3����5�IpI$h^jq��_�<�W���"�0<s�Z ��3/<�L)�OM���v���j���)���&�x��=���ɮ��ZdȓA��#�)9^���x�ŸP=:�(ǰ=�.�m�#+�f���]�HGRY�۴�E�7�O`���k0��죎��1���d��x���O����+����o��8�M�e��v!܄��PX_E>�ƻ����g龣lU%]��>��c��o����l��xlتCW>�+��thzz�C���z���&O�\ɏ�峻vђ�Pg��0�q?OT	i�-�^�q�y"/QWu�/1s�� R�092�LO#�0ܩNEp�V�ohs5�Rs��3Az"f�_��x"�Alh�r7i������;�����`1F�dbI)KK(QDR�"J%`Vm��6���g��W\����5ݜ�zF��g���[�2G����Ҫa>涳A�
\,]+k�ͪ�\#tg�����aa�G�6k&����~<6oz5�4�CL9L�u9��C���w�6�<��z��@��/K���7�oBtr{�U!��Dd�Nme
���*..���Cʬ� 7��_`���=n]Þ��]�r�ߴܝ��fɢ��Z�	��FmF@��� ���G�̤�e^�_G�|i����q�N���і2m�>�.<3Vg�L��Uޡ���#�(M�5+��=k���dm؈tas1yUJm��v��_�-�����{ު�s�v���p��N��J�>�>��?@�Ϗ�x�Ӻ/<rr²r^�����o8�=	13l�`0Pva��f�-I�\g�i�=�R���Z ����˝.�����l��G3@�\J,�e�n�O#(d�b�i�w^�M�y�o�:��U�1{�:$
v�uH�;��zO��d�	ѿED���B��H�k	{�e-��ރ�]=��(cZ��<����rܙme�VU���s�Y�f���])s��V��T��C�3k�t��F�v�6*����o���g��>��a�0FL7��a;�8C�MT�v��ծ�|���e�l9��Z'�ё���G� �	���؟t?S��%B����������ü��#ڠ��L�<_�Fr�.\����aWm`3t�9��=��>����g:�*|���B�K�3Pu�U���.�z�O=9TGy�aN㓱aI����9��	 ^Åo�5{��W2�ڻ�����k���=��x�}�x�����dX�	{3�sp�d��,���9#S���V:^��>sh.ۚ���#<?1A����w㼴\�V�T�g]7�3�W4΢��%��7��ٮ��Z�;3��Ӈ���7s�'�\D}Ō�R��T��js�K��{p�5*d���ډ/�Q�=0�^����~CԦ��}.��w��}=+wI4*sM�4V^�>���G�B��;F����0:�;��0��(i��'	�+E�ѭ��J���U�/�ZWz��3��[Cm2��AV�UU����=�&�[�7���t3�Q �v3�+0�(!��sB:m���vm>q24����ۀ��Ba%����WiL�ֵ��Vk:p��s��ӍqA-��	e�*�PF��ڎ���?\�뿲�J��T;��;���� �u�[PN��L�k-�VR�׽����5�%�iL�M絡Mw6�d�1abWyqv4r^��3BSF�+D�*j�.�V�؄��&*��}���A�ŲۈUf2��in�1�)�sy�h�м����.����B,���
ۓJ�g��z��m�g���nN�ʔ!�f�Y�7�J�d�f+t�m*}{���=ް�U-Ű�,�4���n7��s�����,�v2V�Z�����$��_}�^ ���(q��o6v�MP -%1S��x� M*Q�?I
A�Ӎ���fH��,��%��`�O2!]��20n	���
2�_<��l�}�UE������ݽ�Ep�����ކdrq$��'�������<3���O�݌�j�m����od�D��ܱ!;B�(G��X�z=���c���ųX 0b�yyke���)�^�b�c�x��k}�5V�}jC�$�;�9�.6���Su�Y]|8�Yo��g6t�a.j^�Oe��%�۫�']�������f��|��&.ww���]i���z�D�mqw:��h�!Y�I{3k6��R������F��Vu�+3�e��'D�;Y�,6�@���e\� �ν�K�c��S
�D!�l7R�X����B�L��uN4˕��01�;J��!�/R!���W 4#��9��odV
��+˸P�gX͚ƺ=!^�,H6���n*q�h��Pާ�%��1���.�o��Y̳�W(����WM,D��쭕�X֫:�fc�A>
G���y~���]4�t1��ـ�*���U�Yq��%�hdR
�%�ղ�P���9��l�Nx.�*)@������.g�7�>i����z��W\���vᄗt�M�&��l�����k1|+:�0mc%�B�]Zc��;/���h%�s
�Eȹ]�T��`(1Vg5�zdg:�W ��p	>�-��xR�2��yk��]�t(A�-�-��,^��7\7�R���©��k���D�No-�ݰ���odoW�D�][np�F�u~x;�U�b�kjA�$U�� jʽv�$nh)�9���wݵ}}M���A1��!\{��d���
���!#�5���պ����c� d˩��r�{�p���s�j,�8Y��T���w�O��Mk��ʜ�E�q1y��dڽ�uY\�,�f�h�hWH]uUU�t�Y���`ͨi޺-�1����u�p�Wŏ}J�(�݆eh�y
�gAe�@�-�Q��w�5l�椮�xx�e���l[6%X3Ƨ��P���Y��>��A���/Z}��;]q+���cԿ0{;m�Cinv�<��Q&zU�ǰ��y��MNh�5��*ݻ�`�
T�L�}��ʩĀ<-2��ZC0zևdS9"e�k�g���'���b�ҏ��z>�^�tֲ�_O: >F:w��?9'{R�=5�vg���'��.)�{](�17|L�`�
�R�Rr��<�b��mYc[WqQ�yc�`b�5��}Be�dT��F��>�~z�]v��*� >����q
Ƞ(~��o���sk��ꆹ�A�M_��Qk�qV���(�W%��q,`�۱����[9�l�'�O�+��9-y�GI�Z�7���6tw�j���3dz��QD�G�O4zz��>��,��tN��O}{�Y��-9�Αtj%�1#��d�Y�v�u�ͧ;����RבiCȃq���mec/�����ɉ�gdY6�$� ���f/��u�̖l�\�S5ʕ�3M�{�SX�`�������;�qz�:^�"�� x��?w�R�V��>���U6�ru��ͣ�0�b�\�yK�yQ�Bjud�"G�}��Į��Q�f���Qݥ�G��F�׷�F+� i���Pkҿ#ˌ��ry�T;d����j#�#��������W�$��=y���$�o ��F��LZu�1+R��cH�y8v�5�:(ڻz,��%��L��3�b��3�JH���L:��:�g��ےU��T�#	R#B�1��c�`b�����UeB�Hb�#s(LE#R ��J)h,*3�3�?vf�=eR�B���;|pZ�b���v�r�q���� '6���c�� �n2�9e�:EK�ov����x�n5��՞="Z�VQ��ɭ��{��!F�J��ʕ�}r����n���uW���qƖ�}��>�D��e7"����,��}u��2��t�U���zp�Щ�E�Qq����ȴ��9���}V�Y�M��17��:�:�f��UH��.��5. M�������'K��3��oMM1�3S���Q׾L�H�mq$x�k3���/x�n�xm )7�������1���գ�z��&Y�D�f��۝Mc��Q{�	A=3�+$�X�V;ʳ.y�\Ɓ+��LD��Q���z�n���7V_�`Xg"�Oew�K�)�+�\[y�!>�o��L��`v.u�2�퍩����5��!�S2}�0c��s��_�U��4�'�L�eu#�:{˲�^�/Q�L�>V�����D@�J��,���)�D��N#K�d�t�����un;�뮵Ԑ}��{bV��3Fk�qf�vk���Wp9�(�zo!��9�|��i����̔�(Fx���-1
��s\�oiՖ�e�v�l��TND}E.�n��d>\9�������e��ꓐ��3;7����r/Da�o��Z���t�� "zP=�g�z��:>@�y&�ʽ�^*q��:��W���\�h�`�a��k�P�	pu�Z�+fI���LR�c�_.�Qz~�>���s*F0}*&gk�gcZ���]NL �_H���bN7�Z��pkk-�,gr`��Hz�㌓&�fo�����������>�Y�S��Je�����l�gtW�6re<<L���zWIv�^�<��1'Y�t���M�'6����4��3�}�}�^�NG������6��b�4�s�[#B�ZYv�S���Kl��fՔ���}:��z�f�NR��X/�
��  �o9�9w���??{߷�?���}�X�Q�M���}��l�v�Re��b�=݂L�5��%N��8+O`�0�6�[���r:r��.�b�;1H�](��gY)
�2�Bťhr'�����w�������m���l`�HN��c0�\^2�#v��n[�j2�,�B�>�}��'Հ��R�l�O�6;��9 E�\yS�	ĴuR������ܤ����N���fTRɼ�����9��}DwH�z<6�w]�W�ʩpZ�<4���\��Z�!�|9q�켮�`�wo�Ď��qqM��"���J<v�L�[�ff��rgJu�g.�rs��y�ᗢ��"�:,T��b�`)L��vL�Q�^k4��p�cJ	��Ƙ�wr6r����d�v[ ?��'����~���Ɲ���U5}Э�j�}8���-kI�2Eʊr�%�D�:�.�j��{�CӧZ��rC���,�Q���X2_�A�q4����*T>��SQ3��z;�[��;�˦D�y�{�(Ԍ/F�/�(� �	?b�����iZ�Q��-
�2[m����F
����fB�VE�R*,U���b �$��
l��H�PN�1WM��-�r��ٍh5JG�/ݙ�Ak�n
�m9��t*R�gnײa8b�F�U�<�;�f=�\TK>���S�� �[e�|/G?uk.����M�Bn������>����y�m����+�uH&1HS�S��4�z}�A�T;�����7�V��²%[&e	c�(���T�E�;(��]l���7�s�n�RRyp�)E�0������נkU�d?��E�6��m]��0ޒF��Z�����ccl��f[�!��_}b�kX�d�,���/p]B��<��}�b|V19�;$�O��_. �7]nh�q����FF�.��v��M0a��Diy����UV,�C�]�uW�1}���%J}$x�.g�� �,m�q�������V``��U���F
��oHQB:�X \���U_f����Rh�s��thl��YX����.�_�o����ﵘ?���N0�d$b@D�d�	~�f?n��q�5��=Ѷ�^ˀ;�7Qm��ď H�7nc�6��9�e��P�c|��t]�ʾ�G.����� ֺ��R(��5n]l4κ/@��c���tGF���L���WUt}�k�xN��k`�cY3��U��]��Kx��[zr�I.�����&w�h����wa�[05����ާ�|׆Jɪ������_s�!�R�\N������jW]yW�:�s�CuӒ�:\����
�q�v��l�p@Az���"#�L�3n����ٙC��!Eϗ߶j�_}������(�%���;��� :MpX=1�G4��A��cxΐc��ս�˗���Ϋ�4�0�C�O<ۿ����C�9���$c]N��l40��c�2z|���v�[����Au,��B�M�m굡�B�[j��KL�Q9��Gi�K��tʩ�X��X�эc0fs���� ���r��z�G~5{�B?�S2S �[" "1@���^a�C3%C�1�A�0�l1� D���E�DkXUh�@���eM�K�(xn��R���#%2��]��C��y�7z���t�'��������	B�Z��31;�s|��e����#DAV�b��\�1s����'T���4;�KY\YxOl�9�Us��9G��
�ͦ�6�ؾf��]�4>�N�dlla^wj �>�B���偘i+c��͵2�%b��K�Nh{��5r'����r���7�f�9�i�J�_p�?���UGɗD���;�a�uw���:�J�
9�@�{eіC�lK�u��hL,
��c�7E`�lW�}Gѓ�|����_W���>�A����*���J�f1�tS2�_2���5ָj�XY�ٍ	���!&WZ����(�TQ�4�"�+�������W�UQ���y�����+�Z�eY:3������J́���%��;�
��_v��4�k4���gp@!��Lz#,��O�@�����xBp{w�Wgq ��!s�EV�,c�fHH	�OI`\v>�>�~�<ɟR#A�H`�J�+ ����Ʀ����#�]��p�b�q��Z�!cu�o�8�'%G�tz������w.Ez�l���(+2�9��jJ�
�l0��y�b`V��3���d4��b�`�3���r�R��{���*r��$q<F�5���.>�QJ���d[:���J���+��z[F[����S1�D������?E�G�#��&��s�3�p5��z��Ғ�<�=�{�\+1NK��vI~�-/-��h���Ic)�'���DDs�G�I����;��>C$@�������r���-��%m<
ƅ��g'�ye�q�VUj����r��}uS[e�!�
�U�fb3��L�}*gKZ
�Ka]m9�OZn�3��o�bOJ���{uoTt4b�t��g�Jt� G�tߢw�'��>AU��O�{Le\7�%^s�MY�Z4靀��c�;*f��
1��)�H�+)HTRޘ�"�3���v0�S��+�����T�d"gҊ��	�}�To�r��!�%��I(3j���̗�&\%��k$U��{,ҕ1\�kJɖV�Ei(������c&�[0� Y���5r��I9��W3o/�h��&��tc�W�����;DB��%#�/X��bHs;!���C��>�#��|���)��R�q��K	��{���BHG�gs�>��$���
3�1�uT�T�<���ea�&{&��ﾏ���<1Cx�%��:�����$\I��*z㲤7�CT�k'�}6v�a\o��÷{��px��Ȣ|3[)�V�1��g�>�������z�f�M׍�
dRl��ɇ �'b���[ϤV��/��-���^�Tf���_L�0�� ؠ��C��@@H겇A����?�1e�ݓ���/��O\��(�`ۍ���b�[�z�9S����}6���L.�?dy�UB�X�7�HxY�z���PxV��ݳSV;8�Ք��5��Q�dE�}��~%�U_�ʒ���PqXfo3_�����׻~l���&��1}��8q�v�kR*�SU��Q��Vm^.�w�z��k(
��W(f]�Y4m�:���7;�^J���|1�UJ�X�U������������ƫ�8e�7)ʚ{w�x���[ε��
�NfO��mm��&Xժ���#��fw~�-��-�h�����I�j�Xk(#v+�2���5�j�
�=�o��m�:�;.��=`��挺�4c�f�;y�W���6�;�7�q㈢��vf�{5���BeS�ޱ4�EG^n(�(ӹ)�a��heG|�֚c�id(FZQ`Zf�Y2��M
ZHۭ���%w�j�no.X��7��pEE��nz�4�|�z�w0b�zւGbF�Z�h��5�3���u�n���1¢���r�s�g��s�82�o>J�¸��a#Af�k�M����M�o6|�s����lۢ�Oo��ۭQM2:v�b4�y��d��2ֈQ�rod�b�liš�)���í�M����81�}��w�v~������U�{����z��9PQB�v���I��ٽ�e��k�ݝ9խ�[������4�ێ<Z�8����-}W�*�[�q�;fpۚ!4jN�7M�1w�-T�D�]r2����p�Fq�)��N�\m�瘝�lr��;VV��c.AHE�0n��F�9���mW[�*�Z�T�-m��{����c�%>	�ة{���-��% =ӟm.�w��������qXW�^�I��wN�3'tP���j;̭>l�(��YY %A4��O^��Wq,:�Qӆ��z*���ӡ&����ٛt�Tր��H��4��Rve���y|��B�-�Y�����.r����p�V7	k4;��ESD��4[�W��(�_��}&����ҝ���խ"�2�l�L��q���/5���ՉLv�x�2�>�ぼܜ��*�(�Iw_mc��r����ع�.�!�5�.���]@�Um��h�BP�2�� �Ы\��j����n�F���M�N<�xօ��QΠ�,���]CZ��� i�,�����eX�[ڜՋ[��n��T�� q�;Ct�y�8���J�#W��^��h�V��B -l9�$\u<�е_u�Ϣ�z�Z�M9�^�����\�LD_^�BK�0�VgtZ����X��K��kٽT5�9�`�ʏ].{ɞ8;2�a��=k���^���n�
�T��r�]ʮ�Ok2��\��6�R��9.��$Bt1�V2>��tp��FzI
D�b�Zs]�9J�E��;9�ZQI��Ɲd���^�Mӡ�8d=B�R������^���ޮ\g0@�s[�S����[LØ�ǝî��M[��bX`8�	�ml�+���?w�_��r�]�2�t羏��6xJ��Qv�#7v�r�\�q9�F��qŁ��N�,��ͤw��ӂ
�t��c������G�n�Q���(�l�#e��i���s��*;��D�s��|�dι �
�U����v,�+���uMkq1(��zk�G���}�1^#�*o�<٪�t�]C�b���tOJ������"
T�4ĔK�\-ae��:�F-#�c�r�_�5^����ɯJg{f��0�=C�;��V�d.E,���P:��WKn�om��Û�Q���)�S�~�h��zD�~������=u�Hl󬊽M� 㗄1�\��0��&�y�p zs�\���>��U|Q? O�ڹŴا����y�r�(ɇH�ի�q�&cn�R��U\�T�����Iwn�D30�cn�Ԉe���6�2���;.�l�cm�l�؋����#�&&6��L�`T� ^����-Xދx�����r��<w���R��Nt`/Q����9[ˑ%Ԩ�Ƅvq.�}����4w��_b}�g!��(����~���N��VI���5f;`���iWV��[�0�d��˹�e�>��Q��b|��B}�R����,�E�R�S��{��j^Mv�S@T�x�%����q\]��Z|�������\1a��X���
��*�������R�Mo�^ꌷ`.��A�طJ����t.kX�X����+��k��z�ԩi�'��i�J �%��9��F�`-�^�P���ǒ�ߺk���	�D���T҉hhfbM�4���`��i����>��Y}�]����&浝�[nqʪ��E�}��7$y)�.��矒�[�@P��"�RK!d��"ȶ�
�ƭ	�H��"0`�1X���%d�AH  �B����VId��%hVP����%\��l,L�����K���w��_gdaʂ���c�Aչ��ҭV��/pq����5�Q�'����o����ز�n
�r8HWG;$��g,���嘻R���z�z��2���.�nrW���*B�g�F@}8s�={�r��E�*�.fg�1`t�va��O8�|y.��sU䧄�y��rp��*TP(-���G����]χ�}�Dv��?WtO'Ց&���:e�7ڴWa�p� x�hB�/"�$�ڄ�%�RcG0���9-]:/+��A��#���$��it��馭�3.xb7�9�j���k��gy�GL��"�+EoB�t�[�T���)�iM
��NyVO����o���9kEpo��2Gr��ip69�aE�V~H.�qۮ�߰�����S,n��q��>�-wg�q!�z��~�{ޫ�1����q��:==B֙9��y����J�]�%�]�	U�弪�K��]�������E�i;���<~�Ȁ�������[�v����H�L�,R��j<wrU0�B���ޠ�b�n���̷v�S�rc�V�S�B{�!z�\tw�#�ֵ�i�R\;�W�x�6��<;�՗�� �e;-#�!���gѣ�`c�3��Ӑ��*c�!%Ļ��D���|=b���-��R�܏�����X6jF���v����ゝK���r9�/�H�%G[����{�������|��՜�?��'��~��o��{��[>x����E%Q�?n}�p�-K��e�$��L���q���8����fW�^���z�Ͼo~��y���a�����:z}�yEt7(''�L��A�a��s�N�vOYO	C�߬7x��������G���
�
i��;�1�M��X�ijo*]<�mĀ1%9���jeS�z�^�+���L�j�x,�3��X{�U 0D֒ɝ�7�q3��_'fZ���wgKgIw���)"??/�>�E�)P����������޺;��?_N��f��V��3�2���zc{ٛC�M\U$ޭUl�y.��ǆsf4�����ܞE��nT�^��1�ߠ��T�b	�a�5��^����j�I~�4e}&1�=�sn+7�X�{wS܏ �`��̪t�Rf�軇�x\�����W��΃ԛ��hwq��چ���5����L�Sf�� ��l-�)���RQ�򨱙V�Z���]�,3!Qj�U�m�\�"��bB�+��=�s�E�r�NN��Tv�U7/����=yX������\���9��ף�{]��(�� ��#ﾙ���c굡����_h]g�k���%ͻ*�����!Tt2���� ]<�fr�^P��ݺt�;;�����D\�i�=�#���Q��D}��{����+���lp���ŋ�;ݎǥJ�.�b��8�vqV܍�E�9����fӻ�C���������u���S�<�|�̤؂�����R"B(,��u��Z�������ߴ��c�p��-���&��u΍Hl���ä7�YlX���
u4O`�ͨ�I�;��LKhS����l��IL<�u�M�52�l'��-ad��t���ѬJ��V���i�����Q�,)�Q(?3��}�Y�v�\�n��K��<Փ|�����c8h�'�8���nqY�3˕�R�R3�b{���P�)�4b>�3�,s>�[9vG�H��^��Ș��f��j��	��%���.&�K���.g�dOL����&}�ML�|��<y/�5퉜�
ܗv����D�7����q67��̡H��Twe ݣ�̞�)��i�Sg!����y]7ω�)�;\LJ��9�m�=������R���zz�F��.K�]�Tz_2tP�ɩY�U�U��'�*L��>����E��W� U=����J�+rs�r����&���ꇷ��{n�v;4g%�ѡx3�W?{V�����KK`��d�!%AA��*��F��~������o}y�hw��oy(:��SS�r�]f.j�|���k�%��ڝ�G8�M�U�Aq]�zp9S�jwf�(�Of*��J��I|�I�J Dm���Ѭ�R�t�k�}�vq�3�̩�a��j�ۚ��l�;^�0���ʈ%p��ٌ�yua`�D}��춱��E��%G]H
V�$o�f$���[��1�������祪�@t�G�Uis��N�	���T�[.�~�?LDD}��~��>oʏJY�u�����l���V�1ݟ �-�%�<L^R�׃QQ9�.I���5�wG>8x��ĵ���>��7�b���	\�B@A�Ğw)�C{}z���kE	�Ƨr�@̋A*5	�nu���D%:�7�m��c���
���.�oԵ��B]�[L�%�8�-D����N���N���"sg�J\!�9�#9�MƤ� �͢�5���J̺��kM��=��}�jk�8j`߼�c|0v�K6?#�ɬ�>���� ��12��Q!��R4�)U҈��*J�HE!�*L`U��b6#T�"�Z[)���/��ϼ�����`�(�^i�.��1ɭMd�dڌ�ͷKZ]b�QJ��t�]c�EY� �ĝ���|��m�;�	y���c�:�S���@�3fe��כb䙷�̗2�W��ޤY˝E��9g=��U>�:�(�a��7��2d���Ŋ]ODJ���Of2�okw$�˜�.����m5\��c��"��A��"z���}�[����a��-����dS��so<�d�3e�tg[�X5a_|�9蔯:q
m�;	��iX�=���!eN�Rg�"wE��'k(�u�̹X��+^3��=<�UU��R7����)Pt��e����8��\�R������O�F��C��q�B����v�-F;��Nk��߾�w:OC[:t+��Z�M7�#lr��Puˣh�S��þ�-R��f2��}�C�6���IMc�ϝ]\��}%.�R��?iT)��6fWp�s�����~,Oá��$�XIFT�V�\�3~�bb�w����g����+Q��W�ɔn�@*�x����U�bJDl��0��<�^e)ղ]^���Y�^�S�w�K�wҀq`�\�v�YNE�ON������G�%OZ�[� 9b��S�s3�90�����}�}�t�ze��3�<��ͅ��MZV��EX�.����:�P�x�Ź���I���]j]n�β���<�=��O�șv�r蘗"hvm���x��}r��q3y��b�d\ռJ�X�$a�ƽXw���g����,��ʈ]
��˜��:B^ȩwt��a��s[������Mr�n�Βح8����UA7$#�����X|4G�;�^��$d�����x�)��7��\4�V�����;n7�1��g7���F�=/��) ������ѕ�}�xnS��+7�O�}�7���77;�g�lʼW�<GQ�a��}�-���e��_���O8ÂGUa}�&1f�j���S/7�|6�B܅���Wi+�3�[w�I��(� Ufl��d�eT`=Zp��,�:�����R]�W󞺘x�-�lU��Y��� dl�=Vm�3~+ ��>�x����7nl��J�c����x�tf�ф\��;�3/ ��N�n8	}O��/D{*�|�T�O�� ���|N�Ct���B��}��8s�n��rS5U'R��{,��rB�4�x����)y�����z7z̓G�ճƕ�K�XY�Kl�Y(���o���t=v���LH���\�����{�8>����=}:o���zr;�=�?m���c��j��bhewW�P�P<fbZ�u������R�vJYA��K����C]]2��Xg>�W�.-�5�G�"b_�ݭj�I[+�H��+P��j6W[�ng�i=l���\�D��,`<_)�`��OX�������k9�^��d1�K)Wk%;`����9�e�-���^��CNZU��e<�jF��}�h�� �`@���4��G>�[�A�A��F%V�y~(�+�i�,~���ˁ���	��)�ڂ�����$����_��AWA�ׂ�/W��p����㚺����Y�4���u�ru6�Qji���;�����1əi�ˉ��J%k�7�P�W+j	�M!R��G�>��'JbG���W�����mhp:b���>�k\Z�$�U�H5�&����Ba�e�E�N�����g��"���H�M
��T&0�Ɨ2����u*��{�ѸC���8�c;����u�90��{�)�9���7m���^��gK�)�\~td�T%�{�`�i����>�q�{�i������g���o{��G]���@�J��Z�ғ)�u�M3L�So�2�
l)��μ|zt�-�]�|1�L2FiX�s'J��P���RR�PNb�W��>H����惣�X�Ru����0�'�gV�z��7ur�Q$�w���1����0�3��m�67㨾���{	[�Pєܷ�$ڿ��Uw��_��H��GSg�)<�]?��#5���Qs�p�|{�U�T�����2�Fs2�2��rE�*�����A�|�4knsj���!l��c���3b1�!���i�<��|�RM��4�����y��h8Q�`5�^Z�>�Z`�N�%�.=qk��R���$�a{���8�ao��BA��b�Lj�4����6ؙ͋�o���9�F�ʎ�[<������t0�4J9��=�g)����ovlef#
*r����]�ú	��g��"�h�� ׋�R��%I|��W�ķ��qD���S�Dc<y�����dO},b&4X��l	9и%��M�<i͸�o�6���n�ٗK���Y1�(i���kF��;{k��I�mm:�J�M�Y;�����49��H���/Jys\ܾ�U�[z8O�3$ݎ�e'	���8�6�ݔ6]L�y6<�c��%6�@�4�S&��[@YB�ܾ�����$Ջ� �{�V�Qv7�2ɾ��s�W�u���rY���k�x�5P��� �o�9�u�+�7:]d�t�h��`J��P��l���A�u�'ܯ�Dy�r�w��JY� �3�{d\��㏍��u�� �X1��cɝ�rP�yӐ�x�#��fh(#\[!�p�k�K��2��ې��	N��۵��G$�z�.�[���Vf��1{ǰ�u�i`�k�����e�b��$w{{��XJ���ԙ}Ml��Gn��t�0��͈NN�ؚM�n*�u�[�r	�WP�����Qn�Z�6��:� �����z�V���WW1+jã��.@��o�����B&��9�դ�/���ղ1�鳅1����̓�T�)����r��=�W�<�?}�w"c��s��J9��m9�n����|퉛2Yٻ;�Kp[��
zm#��9\ݪ��]hz�P��O���q8Jf�sw�{"Z����dS[>U�ߺ���lX���s�W�={�p����{�Jk�
������ck$22#w}�����8�鍣?���Tv�
�c�1���4��TL��/72ԏ�-j��ݧ
�Yu�g&r�:d��=��нu,�D����&+���/g��aj�;�i��o�kį�4�0^�d�?H�T><��>��J�B�|�r�vGNv��O�o2U�����h�5�3Elqz[�}��r{}%� ���B�yh����ؠ4["U��s�:��9�"��0����*bQEF"�Eh��mKX�D2�1Z�Z�XR�Y(�"�Q�-r���ԍ���m��,�2��D��iQH�Y��GSZrR��_���p�7�s��7M�7N�Т��>�Y6K��U����ϫw�]�1���c1�6��HC�^�.�2�僽h��������n�rh��1����b;"�K�	j܌��+���G���\Es�@�	a��w�tQ�<ӷ�����	�^��x@�]����!.R�;��2��ʢ_��ھZ������؀�{޳�]%�z��V��2�Oq��Ԇ�G� ��_�W��l��ڍi;�goX�Xq��.��sH+��D�@􀃺1�w�a�I��c�n��nb��o[*e��:��S�/���.y0"UxCҢ��h0�9�H���Y���ܜ���fz��1*�Bg���d�Z�W9\��# �s��~����P�凃�������l��gY3,�۹.�N�.r�h��z�V,�уPCN�)�z��ât;�s(����������ڋJ}9N�a}��(s�`]�m��}.ϋ�k��?o�u�|߿_�8���PEP��\[ �H/1~��m�zv�n/_G�,EwSo������G���|lk�YK�p�v��\8�s6���+ݒ��p6޿h�c�h�����x)�2��7�=�FD��;*dx����ѻ���y5���r)u)7���q�8���(�SfF��H:���wh�SC��[�e���c�GEz����F���(�Cj��Y����jd����.�[�����%�m����0fS�%��DD}Y7����&l��'}&˜�z��V�k�D�%�ױ#��J�g�op�j*�8#k�?��<q��
[D%Nv6�\;����箺<�~
 ��f��@�1&w��F��t᭞�M�$�3�Ոs��rF2X����yN�C˞�5+G/���ag��Q����ktVƢ'����T�vg���)�e��=M.�����ٷ5��p�T'���}��z�3�В:�U]J}Z'�1���PP4	Q�)�/e�����z����N����,�&���nJ{�Z[X��&�����]k��)e���5ۈ�os�M�{{��^�a�j����u�y��إ�C۩�C��̱�� �39�L���T�4u9�������i�r;U����`�xl;���	a�<���O�{�e6ِ�2jr�#UJv7N��l���pXz���L�^��i��_��(�s��)�8'��66�6��ۼc���*��\��)��Q�&Y-ް]�k�No�8�����v�=:t��H���Z�����DZ�}�(z���|�p�U16��,S����9/l����671u.·\әT%0�*&Z�[`ĸL�b#}EB<��#�m_H��nyۗ�֡m����z0U.�����&���S�ي�R>�"#���Y��0C�����K�.#��m��°��'�_�VY-��֩�ԧϯ-�������O�XJx����opN�2�+����y�7� �q#J��V��PR-������g۟�[��xkV���zX�5����;�Q�t�+`�]"��c�O
����ݫ|cO:k*�R��­��!lx��¬ĸ�����v��>����ݩ9d�z&uA��U\���,�\䮷�r��׭�Ikfy��X��9QE.@Ќ}����Sˀ�
m�&�#��6ʠc�5�[�:!��|y�K�: �\k���\�s�����%�"�t�<�ު	���G��mٕ+%�t���Q~�����L��HU2Ъ(oV�H���l�E�Յp��b\tP���3�I5����(b�$jC:�F �<�j�Zu��+QɰmgCLb��jV������,��`P�%�3xv �sw��������7���Z�;8�>�>|�NN3�֓+���O*��Y��!Nƍ����� �r��;n'YL^��e4�g�-��e]қ,��%֛Ͼ��J���p�ؗ���]�t;�lT�Ǧy��h�6���S���IO�D  d�>`��nj���Ml�\�u�̾���)ڇU�[{��_���w�Ɖ�h��}�J�]g:Y�ؕქ6�kY�}6���K�Iv�D�9�����f5."3(��rDMo��u�8b#�\Ͻ�h׼�@=t���ZE��N7\�y^��1-|�A�����K�q�t�Y,��kJ+y�s]�"^��-)��'rF�jɨ���
��F��*�fd����#P���#x��]=*��ku�����ŧ#���X�.:��s����R�Ѷ�V��Ӷ�;0��{����Eg�fݗ>��x�dX�g�[裉5ڑsx�be��%<��"�8����_ tb"�RR3f��[��J)5&��A=z�a��^��.T��tI��=)��Q�m���>������`b, 6p��sˇ�/C�w���r}55�{,ﻀ�T:g���bФ�>��{΅��]�7�z-K�����T�J�G������[9�&S'�+~���<�:�[�>��y�1?��>�5�p��e�nD�±��
�D��X���mb1Qk
�(����@q���0ʸ��4P�.Ffbܥ_��P�&):�<[<0ͻ)�]H����������ie���׳�=��L�if�α�����Aj�E�Y����QӴ����H3y2�dJ�5zv��S�U۱ԓSv{�����[b��Poiʯuȕ�f���:�e[��ӿG�}^V��'}X*g�ڌ�A9�4�Et淖5���|gkd<=8IV��w]ir\�%���>�P^���ʉ6���~��i�2������7qYo���c���ݳJ���p��Uد�^�O	��dtec��}_}��	��M���i�n��>��#/f����g���N �崱2��Κުi*��d6jp��n\�Cpg�q��*n���k��>�s�V3Ѵ�oT�k�~���r�
9묞
��fG(I��e�L�#�ᆂ2#���m��(,�5>���ub�G��|�J�͏��ߴt#x%�3Ԇ;)ּ�϶����.�]�x�����NDQ�T&10Z~�]�c�'�T^�#����M��8{&�P�̺a���Ս�ox��&�:����{Brۢ�������m*�R��ys�)l��lN�Q��>�>�sBfbf�ԍ�):άSM�k|ʉ׌�h����Bb@O���ڰX��ʃy�:�����l7�E*�5�}�>������jw�!�e�K�KA��Q��4��-�����»����S��PzI�fwC���#�LCf�B�>������*vɞbwLJ�[���v�C���J���<��(6&w/��]�4^�M��b�!�d�rn�p��*�����>S��jf�k�[�h��|��@�6T���Zt��ݠ�6O<���9���R���3k�:d=
s��h�k�2M���{��Ϙ���v��e�#�^�v[:8j��*d⩜'��z�H-;֞�n��
�&�U�6�~]i �ceS.�c����ŕG�L7}�>���]��5��g�<4�KkX�@��$�����c�m�>�\�V���ʣ�ޖR�U����o0�NL�jdJ�d:t�y�0��/�f���oz�x����(و0�MNT�e�`�o�G�u&�˩j�-'U"'�Fq���87�~����DE�֕��wo��Ռܳ�Q"H��
�A_�L�ΨNJ�X	��Z�]]*�t��c2�N����t�3f�	s�}��� �l��oIx���J&���!��̫7;r����20q�$z>�ֳ�u�i9L,h�gd����P����U}g�*���SՄ8���n���¾�S�#���s����I����@BX�eQr>���rW7�R�f$�+@\L�^<��'P��vK}P��V�)���/�z�����X��p	�����|K��l>L|�\W�t'�� a7�D�h�D�m�U�(WwU��-��W��}�ﰵqtp�d�r�u��{7��X	�8�+�;��}\:��5 	��A ��/�\�IL�"��H���T
�0
0�.��	�������T^��Za���4��7��˨��hn�nS��z�U�N�V�9r�_�^�[�I^1��ԇ4�uzx/EAy���1�e?�fѭ�Bߍ���Pz*I��Y!wV�C�`��S:SrXX;y�j4�d����.�[7)�7� }y"���]wδ��@n��v���^T&�<��UN�jӆi�-�W��{���-���#��nn�r�O�\�N��Jn�~o?:���*Ŵ�";t�{3�[��l�	ӭ�\���$K,�K��3����ڛ��5,b���aS�>��ڲ�ϰ�9�.r<�UP,R&Y;ף�55���@s�̱�:�ir�E�l�(]N���I6�ӈ�*�j5���qm@������< ^�n����ķ$'��mZ]��:���t����:�&��ɂ��LK��c;#�`H��{�hx3���A�+��ҼX�/ ��V�A⫸Kȹ������T~�����B�;�'gsp�]W[�u�����k�E���3����k�x�L)L՛u��jg7��H��WBP�ԁ$A����`�C>{'3J����2�o[dX�@�֝|��t77��o3S����m֝�n�ĴD��h�l�^�.S&�\j)�3l1 �)����@Jʕ_3`b�+�G�bq��p�6�44Q5vT��o(��O�lM�^V��YE2�o���>:����Zv׾
]�Ϸ���4iRhte�z�3��s0�!�E~�Bdq�]��I�X�:�L4�:������-QK�@�Y$�V����O�eַ*r��殻��/�^]��Fw� (
Gt)lr���[$Qݕ���"�
�:�ba�"��P��cfQVs$��X�m(�s.�Նg�P�@�x.��~�Δ�s]��٬KM��Zb��c7��xǓf��ڣv�hp�[@�v�Y)�x���?0�4��U3ksc�͸�/5��w&�sZt�їi���m��h�L�x�*����{ �}z�{�CC��yw�$?3.@��*)>{+�m�Θ���r�bg�=�aP-P��8^�m
��ͤ�q�L}Z*�}�fw2\�ȗ(P�G^��T�C̷o��3��s�7�Ƭl+'�ٜn���f �t�ph�ɼGK-4CT�C������p*��F��[�`��o�7�ȱ��0
ŕݾi�\l�G�����k2wvEXk�e��,Ys�(�9�VG,!�N�r�"�y��>��gP6�h�]�E�����jf��t��w-�I����-�O�ᮗøZ�ѓ�!�ȡ�\�{nF��pD�R�s�jT�.��0	Դl���� �`�;�XP�5����9w���$Ȟ�ʼH��9�,�&��Y5�Zՠ3!eJ!g'˯O���#MZe����l��.E'.����ҚH�/�j.$�����,s,��6-�XyM秇xx?a�5�7���Uo{��9@�it����u��r�4q�a�|���RP���A6�ֺϺ���͡�m%�r����Y��eF�ҍ�_��RΦ��6����kzR�`u���nSV���s���B�Z�ՠ��S� �:�B�iFRQ�Z��u�+��i:��
�JYwPb��C\{w�uu6�SQ����[�|�ΛC�|��5<�5.��Z���&��XG�:��pY#g��ne�X��=Sy�����H��9�|�:�*V`�8�LSC�r�%h��.�6�o�}\^�@��aquP�g��:�^BQk�<y�I�h=9�����H��.�)���r�=�0��W-�C~���	|ٞ�ڵ���(��vA��9�J�nc��m1�Z�4�[�mh䕆�����,�j�1��$?���e��@��E����DM'��®|Z�����V�>��ޥ�����ʴf[NM�hd��vY:M�;=ǝ��wN��:��u��p��!o["9���z��̀U�°�ͤ�i���ldk�ү+h�6���e����S�����Xڳi�D����S�i����<���/�Vgʩ�.u8�&pk�S���u���9����g�1&��sA`k����ۧ-���|�K�����O�mX�U'�O�(P�AA�?���V9 &�f���g��܉��d��Jxpshfb@��8z�y@�C(�U_W�ׄ>Hu)����ޙ�����2�)t6w��켻�`�{2�F�%eIj�Hm�=�/M\bյBfښLT�5M���8��ow��Z針�3��A-�-�M�b
��Pb� K�hc#�@�����l�ő �V�2�TƩ-��2���W E(��4�
��Sl�3r�\��h���d��o.��ʒ���$�\j�TNv-]���f۱���b�v�+{e1���X���	��$�������p��덨&�4�PsN��!e\��6WC%���칥Iw
PD�l�@Q|
-0h{ލ���8$�o�	��<����!4�%B#�z�:�2d>*�q���)�=!�͈�Ĭ�O�UiA���HWs��d��U�"�^��u�Z=&�T�mK�x��-@�����I�;A�����������v��[8,�Z���G�t�\u[��u�X2���S�n�W<�I��u�ru�R洦�]���?C�96��s��yH�?����0G�\��5�<A�}o-T.Ԭ�g.�m���x �ˏ�un�Qv_V�rK2lJ*w�D}�)�ep���z����Oj;C|q6Qa��ٍ��P�}�;-2=����/k�c��!@X��G��W^�X��R
G֢�z=�6��������9IՎ��5� Od&E�;2��(*�p��9ZhNj�R��V�_d73�;��5D��1%�曔l�sz6D��÷�rT91i��{''`��,��(��'��S�'��{x�8A�y;��}���+#G��(i�"؀�U��D�;�=.}�w�q�S4]��@cg%n:��b����xZ�Nn]d۳��B023^k����@�f�0�:E�N�D�k,��O�DC�E���F�4�������N�T��	N���C?$�f%ĵꀾmٝ��aG�����en�^�z��V�ೕ����}�R�BYUօx�R&'�c7\���h��_kT�e��I�r����4�t���|z�k��4��%e;�&N�^7o��� ֪=��������(o��=�v5���B��6��z�%�%[i�m������tv-��bK�u!"г��#Dz�������T�{��=��2Ĉ�V�:��W����jz\�Rw�'̆�E���u=�M5*E��E�-�P@��h�c뻿h��{CJ�ђ��wyV��\ݮKR����U����LmmMŹ� S�Q��eNV���e�����\dWU�mb*�=
Gb�ݳ�D�<T�	�f�91�1����WN����2P���in�'*#�R��)�ș��Oo+�j��#�y����(��t�G��TĞ�T��ё�o�gy�r'�.����Y��q��*g9��9��@h�J�
��*�j�ү<;�8�m�K>�]`>��=��{>�g�\���8�<m��uUb�Ⱦڄ�\'��Y��H���^�����m�e�!�N��_s���g��wYщXt��d�ٱ�G�1�jG��#�m	VF^�rG��{�eK@��l��ռ�|�+&o�s�bk�J���a��2Yu3W!P-3_}/�����=/�5�x��۪�y;j�¤蝀�O@{n��T�d443Z�8�ko�T���z{M�� ��*�.�ܿTm�\lF�.���<H����(��d�$�_">�Q�ʫ���N�Z�S�4S��ך�����)�1�5խ�]!}G�֗���q����'J����kvUL|-�!�%�ʺ���}Ӂ9�RԲi�h��x�"�י�l�������¢�dQ �Ү����LD}��r��:���bxZ;�^z��3ݗ�M� ���+�Z�O�dZV�w���(M�.E��芪�[�CWB�':����_�����?m���~����LbyP���9�|�4�X}+��;	�I2���٪Ǻe=�*V��̽S]��c���֊�ÿ���1(��@Ǝ5&�@�.�{*�]�BwJ�eҪ�xq�b�,��l�g�[\}�}��m]B3��]�ݶ��F.-i�j�m��m���IĊl(�l��J�:�C{no��3�54[�K=�"���SDv}'��W����΃�o��b�tٗR�����P�HN��P����&���{�s,	`��̴��	*B�b�"�@����_���L��]^�)�HV�>�o����^��8 �l�wn}S���꬐	g�H��T�)��Y�Eݛǆm��<�;�ܮ⑧��G�?`tG�0�?�l#�t��E��+�\��Qz������.�d�`��G�@�UJ�����}%Fۆ�\Kȕ�ve [:��icl�1�0��iF�\��]��'�Vls�%R+>��P4�w���82G�}�R�9G�}:�m�/�BVH����V���"K�H����� 	`gk�`�8�Ƽ(NM��C��u��Ԫ�%��;���޾!��	a?l����H8�~���e�G�!�@=�<&�):���^��ﾈM6�©{ا�B�v�=>�}��S���fa�{2�9S�M�+�r9�����b���]J��+����/���)U2�9���>�Mb�+��*�kC�>�>��u�Ӵ�S/:���q��3<�c�(}�J!�(�A1�B,�� � c�K$��PU��D�(|�{F�!E����13Q�6��9p �^�hnr�B�eˊ�!)��_4Gt�.[n����W��\��2��tܽ���]:>@�Q���M�:�;2���)
R�Z&�@����Tˤ�W����m�c�EKS���N�C
n��Ggeq�q�څ;e�M�85/5���d�eT��&ZdpŭZ�-����
��yu/�UN�L�Ӊ�9FZ�r3������Hh��r�xS��c���~Ծ��y��;�^��rz9ͳ��E�������O/U��3�� �ӳ!R�����T���E��]�������>!7,,�UUW����Eܟ�ib�zʛ����7��:?Dk�8�~�DZ: �g����v\(4�ۅ2��� L�N')<�<�������F_nU��C�������3/5_�D�3��Ӯ�ն9{�f&&Ӗ)K�p���7p$�K�kI�����F�xq`H+d2�j������
R����ߎoon���g(��W�Ԅ%oD+N�t^- @�mǯGh�ލ����k���2�1�sF�)\�G&��9��f5N)�olL�B�K��jR ��syW.�S��fe����%�+�l�/�9�g=emܞ�]:��2��>Ͼ��n}x��g}S7�G�
�P�M�̪L�5�ː���j�%m��էu�PC���B�9�̝���b[DBq=�������Џ�נ3fY:wV0�u�t�5�M�É�o:�܎�����r�b`�k��!���w���ʼ�Py�H��|�4bIu�v%�<���e3�Gqi�}m]�����6�Ơ����޶ ���SHη���z�K���>���=7_UK�X�{՞����v1o
��d�2�T��Q�PU�=��	�Y=ږ7P*��R���A����������ZH7 ��]���R��� �,=�z�H�wp��9;]!�e�������c������߬���՟��4�V*�#&��B+Z����;j��f��G=�����i[;Mf��f.����%�A¬�5�$�|�e�ٽ;u�A;����(&2v����J��f��ÂJC8]���S�NY�q��h�;K����[��۝��a�d��7d	S����x'Z�ή@Ɲ��Ѽ��;B;u�������{!��8*G�D���%��$�"���o<A������1�9�]S��_�%��.�/�9���yH�ך:e��J
5��9�)N,*f�X�vdX��x����:K�mpt���Y��xby���P�z1P���A�U�W@��9�ƧW�{4���]u������4$V�;ڷ���%+�Ɩ�`����=����dH��jt�79����ݻ<�l1�F�,�=�.Z�H���x���tdv.<٧G9���s��wE���Sa�s���-/F��Vy"�boLY����mA|�J2� ",�B��O�%�}V���߮�"0;b>GoNc�B&�W1U徳g�y����r���0��^1��/ S�Z/+���9�l:�;��M�����y�$d�X���3�v\�ɘ���Q����=��|{&D��|�dhv)a�{HRH�*x����B�ey�0T�2o�y�Tg�9�0���)��Ų�&�h�Ja�܈���h7���;Z��f�=�����!,6�c�ÈΨGge4���0̳�7�q�`��v4.�;g��`�3y<�M����jt���)��=��L�nt��`04��C��n�Q�;������_Z�s�uhK|^M��l>�^��f��]#<=������;k�����V�QFh(�fe�;O
���:-�<{���T]aDE����Rj��������TBp�E��2�z���:5���p˜|�XgsHw����Ş^�f}t��y߶sx�[}�~�� �	$��@$���@$���	 �K �	$�x�I'�@$I?� �	$�x�I'�`$���H��@$���$I?@$I,@$��@$���H���I'� �	$�bBI	?�BHH��I'��$I= �	$��
�2��;]@	N�����9 ��>�_���zpA�X �a��+Z$�%"��$�*�����E��M��T�(DTQ@R��h�͍ �E)@��@�  p
�� ( R�   P   �  
 
         P   ��{� P     r��ב�u���)�{P="� =7���� ��#�WP� ��T��A�R���Wf���6�v�YE��^�ټ��J��� �t=��G^&��۞Y���o'QI<l{�:��ޠ�Z��k�f��s���/f�ov��.֢�b� � ��      ^� ��VJ��.��.t���������MM��;,�T�ݶԤM��� x�\���rz{=��lճ��j[ەN�坦��x�'��=Zm�� ����Y+��ޮ�v��o'r���)@T��T�&QC���6�ĭjS^x 9Ey���sn��f��W�.l�YR��Y�v�o1����{�P/Uųl�j����M��X�4�e�ǈ�Wl�{��㻆�h�m^�@P'�v        /{�%W�ܶ����y��^�zb{)JS�ހ��UL�w�·vy��^-)�g^�[[^�;�OM8� ���V��uy���5T� ��[��yS�t=��G�  ���w54�9���^&�����o ����3�l�+��\�N&���\���l� � ���@      Δ�X�����z����@�ؙ�`�����m=�t����V�{��ڱ����z��z��K�Z9=�^���2��ʢT �D�x�)��.f���
�M)��y��<M.��9����<v�F�� 3�B��+�vvx��V��nl���7=�E6T Uh�@�        ��3�TW���`�*q���Jx� 6�b�ͧ@.`n/s�纄��s��� �(�{��FUy���P ��cEW��[Fm7���o1�[=/;����]�u+�і�7v��]�e�
������x����(y�v�=�����헍��&K騥/p ��И�U  h )�IJ�2& ��#A5J���LAF 41��R�EH   ���Ԫ�   ��	�U   y߶zz��K-��NS�~<w�����M4�}�ii5��~\��B��m��UޒO�T0�Wւ������t��,c�1��O�����9u�vo?��둙�Y?��вM߅�W���v��X�^Y��*ZYE��֗T�3��a.�8����Y0���fLalW�BX�ŋ7�8kX\#F�R H��sM*����&1�����f]ɹk���X1�:�V8H
�3G�=�n��h����T]�$��k;o�T�X쫵N5�!M���顯k9b\,����5tGѸ�m̙�o�/���<a����["(7��4n�[&EN^bq^�N��K�fӕ"����sm��B�7�,�8p���"lff*�hSt��*g_!=x�Ʊ��r�i=�َ�cU�\�Z�K�7�s�H��RIP���Ѻю��1�̺�bH蜩F-ٕj��DE����W1fE=���xHy�xe��bI�i��Ҳ�L:��g&�_�ZT���z�Ք����c�wr!���B���_��B���sN5xugëh��`y�FZ:�6zK��3��Z��%f�ɔ�D���<ޜ�}��dY[KU Q8��"��Bk̅���/���Et�t7iV����&%�n]��w�u��n�TKF�Y2adXфĩ����0��ŀ���\0��0���-1i�L����\qs��ظ���.�0��&adX��C
\%�]u@�[gz9�3'=�ـС�f.Aaۄ��3n�
b���r�QY*f�O+��f�"�VK��v�x�)��k6��P�⏹Kݵ�,}>�֍�P-���>�a��Y�Է�;�kxݭ�zI��g���{��$��1��'����uR&���u_` nVZ�:��UN���,��^7:��+뫊�o`�䝕Ք�������.��Զ��!����c6�^(w_wc�*!�Z�횛�q=��o�)R�:b;{�X=rۭL%L4�T
#F+��D��ez�x�w81XH<�s����9��3mV�Z��R>���7�F*�3S�Y���v:Z_��#���$��[����q��u�e�Gb\�v��mp�q
6f%���v�YHU͉�(FӪѢ�^;Y��c$�VF,5��Z"�B�j�X`�%"�7�
^�5�M�Yi
�Qw��z��gF���k ���@�ɇf��+d�NLPQ��XeD=� ݃��/qT
һIő�n�$�Qk֞=���O{�ږ����g3���F7�poJ����� ��Y{`٢��4){�@�'��t()!a����!�3���C�Ȃ�&���ƣ�d%a��i�wZ4��P�a�SGB���4��t��z;[�D���@�j|�\��c�YIǬM~o5�(٥���4;�N��&��?�G�^S�m���ތV�Vn���PI��i8�
�x~N�c�E��a�YOQ��N��/Xr�V�IC�,�\�Ԧ��kvq �4aka�a;�`4[m�:V�j{��!Ĳ]��
�+��4ljØ�tܻ(�<SpaN�D��4�Фi�R�Q����f�&jM@7r,,�����L�T)0Ԫ�"Mim���̄���tA����0Fn�,ݗ�E�˭Q1��J�`��r���K�S�
�ʶXK".�6���c2Uج�Gij��n�K0�q�wG��C!����+�8 Ǡ�w�
Vnd۠\L#���Ne�fV�9�ń����$*6u��nn�1�>�^�F|(|m�YQ5N�b=0�E��	��n�]�Q��T�QI��H]��-�J��ܢ�0�����Ufp��P�16�2M!�ڪ�#�I�Y��(7cSj7�z�)n^bniuVcYU�iRn:P;����$��Lw�]ZV���hӻ$����]ay�p�FS,��!e��9V��(�Sxra��YH#�6�څU����#|�P��bG�]�U���3��}"��+�dF�4]�ec=k
�Kz�3�� �0��l��MSu�+���:N�S:���f�jc�R/k���Lޙ6���#6Z��Www�� �^v��m�;cZx�˵��:���n6�9�V^e^�Ӈs��	��m�,<ܖ	�墑�3\{��u�5v���)��%(H��~Q�R'[��b���, UEh�j�@ģwdnإm��m˦@Úf;2�e-�/0�ˤsi��C�@��B3�B�QX$mI,V�/M�VM�j�������T�AT�2���m�n"Fl-�ن -M��[;x2�[��'�r�ؗX�̘��H�q�rn<��H���JV#�.��If�:��5ko���ůq�~<�*�iF76��d��4������qe<�7I�[T!��H�&#�IL@i╈H��[�0�3")U+�{D����Ŋ�41�"���LI�fF�P͚D�7�V�L$;!��aĨ6 h�J�H�+�1�x�&�-GaQ:������)赚���eDC� \��$��r6��t��1'e�,�Q����D�hj��ȵ��]Ϸ%���¨���3�rʸ���'J)`o5Qv�J�b�#6�ݜ������V��n�T�[#�V�HTY��U��ݙk ��!g/F�l��f�%�$L(^^!�IF �Ȓ�
m�d�d�ʹ��L���u{q�ۖn������i�e*�޴��C�á���Ym�˩
���E�0��V)J(����֣:��.mn�ߦ���@�4�f���Іj-�M%[��E<��QaޝY�O�o,�|�2r-�i��5��dϐ����AEd�̒�Ϥ��Ռ�na�1:�1=�z�F.$��J�6�CE��`�J����ѴrQ��6�dP eAli�.�N����#�m]i�nm�;���f��ܚ[Z������aǑV)c,m[��ٙAYn�!	�.U�9��)��âUۖ�h��[Wx�H�-c���I�!��NH��7IjA��p�$譬sd�ɗ"Z��^�����,L�2�@�*H�3*��Q�+R��T\��&�IKv�h��6]-�NLZқ�e�4��n�n�+ܕC���]7��&��Xn��r�t�v��з��"4�F��@"%n�n�3#h9P!0P�F6�hvl��]]kې=ȶ�������ڌ����v��)]������bl�5�����A�Wu{�[�:[�VjxΌN �{�@��3nV��]LPa-�`�y3u���Ec�j|��TY�g�P�ka�"�|��r�g%`�:���� h�Օw��)F�VM�.�`R�h%r�*�cGJ�V�Ӷiʼ��^VR��t=y[%l�Mɒ8�/ٖY��.��6� L[4�ډ�oj�
�t�KFE�(�jܴ��#!����@
$��հo^l�_׎�Ӛm�wj��$l�����͊R+)ݯ ��Z����md3(f*(�HQ?N#�ݦ6�XJ�n�֒.��g>�F��l�P��N��^T�n�ߌ�y"���i�#���\����F����9u�N%mi�9�c۲46I����Ԕx�B(\)�Bw=b�����G�o���r���M:(�ks����v���;X��xK)�s%��]@�Ųn����u�Q.�l�!�,Z�Z5���%:�Y*.�㠓�]����
�,Q�[���s4�N�3�C���YǍ�*vh]�D|,� t�Vw�ipX]:`̋BɌlXTX]1�H�K���2k��#�����[ċJbV�iʚKvdLݛu6P�ݤ5�E5s\M���&�	7p�� bͥ��X�FXݫ���fV�]h����Z��錮�ȝJ������W�.��')X�%���Wb&_U�Ș���ah�m��a�\�}��	u���cm��o���ob�F��FVT��"�B��-���cFd#������XB�Qhfn�OK�R�]��X�Tץ�fVr�O�b���k�0�#�o,'���Ӽ+pM*�l��V�j��؆n-���֘X:S�zp�&lNȚ���#�l]��
û����:�z�:j��r-$E�!�K*�ڸ�a��h�-�x mn@�]�2���׆�PQѱ.��LX"�D݅T�Y+L�s&��� �G@	X�Ԙ)���$�R�L����ӰT;��z2�oK��2�n7CaБ�
:[�����5�E�Ǒ7�|N��f�-���6�-]^���Ee�Qͳ��ʫ�?�����	]�0�|x��]^ڊ�m�]�yY`�hʕ��V����3T��4*bP�6��1��u�5e�Y��&���hn�m��^ףl��V�=���v.8Sm�0Qǂ]����P�Y!0�:wY#S"AV�ŵ#ȷ\zV2��T�ώL
��M1�(c�Hp��Z��C�E(�W�I�BCe�I�yM�9�=o]Ϝ���>ρt5��jt3�����6�d�rY�V�~ys�L��U�
c�׊�Sv�r��kEՋ�rh!��Z%�M@`��X7l����az�P���`��n�Z�[�94���j%+�2�d C�/^����ױ"I�ZUd��uW�fD��0n9ϯXVk[�I1�M3w�,gue1;�bp%���~��p�
��ZkF����9�I�����)�C\�H�[r�WI�ӕ��Z�0�[J�*�g1`g��['+^ǋJ���,/%f*V�,�X�m�&�[G��ݺ'd�����)0��X�L6�#�䧪7r��(�SW��d�6���&�ݩyu�[�hc��C��{��*��7{H�86v�i�)��e��t�b��C(�� ��R��	V������m]�@j��Y"�I�l�D�p��ϊ�d�PL:��k,�i���Nۂ�M^�0��l�Q�ɵ�V�nѻj�v�0�WI
���f��ٌ1���� �'v�C�#.�ӖC��5�{z�ȩIS"x�MI�Y �nfA��n��Y)K�R=(�yvD܉��eܹ��%
�&e#4��@�Xj���8q5/cHk+^=Os��V��"�Z�R�R�q+�R����0^�j��f�6���Zv�m���޳v>a�WYkM�HXj(Ez��#{��vڼ��rX��	���:�e���Ֆ�2e�U��8����r��0�Wct��P�4��H�d���Qk+6C�*��ܗ��;z�oU��Ո3vjARk���Gp�..5��j�d]�n�� 8�pAP�*p[7�fU�(��5V�Qc���]�u1дi��u���e�w���U�L��Ȑ�y���\;��Xy�vd�z��ةn��Yx�V&f�F�溾=/ 6�z�����4�����,.�&,(, XPXTXA�w�*�:�:cRr,5��fE�Yx\1��N�U��K�pX\O��y�4,'Z�䦪�E�Mp�b�5�����9����;c�4,C	k6,-�+.՛Vx�߭π�Ҙ��ü��$���wz"���`.�x�)']kRڱfFwsu�Y�l�P'd�@[gY��VY!�
׬]��R���0�v]�]��
��]�6Me�0"�!�k���S�ʛ�)P��,�j�\�Y}Y�j�5�x�1MtڣS�7z��p�v�o�7�4���l�t��nU.��)��ڻ2:�O�1���g]
}`�G2]���]F�1�,��V�\�f�Kcy�̳��j���3j<
�7c*#�<[v�'��=�ɍM�W[ñ��Y���v1�i1��:ݝ�&��1�jȜ���x����3-^.U���_6�ܾP�Y�Vx�o�Wq�_Cud��K��F�6�tZ[�"o.���}wi��� D�R'5�1�s�Ϥ"�e�J�#+i2�YmD�Z�2��;7(&Ռ�)�
l���UL�XUU�zC���3?W�Cj�f]YT���CZrw�9^z��5�W,�u&0J��Ħ���!�@��9}#c_c�����P|A�5�>[���|җ6�ge��tpJZE�z�o}��Zj9[1z&�y0������C�E���au��0E<��)hͳ9!����J\5iG��*cS��n�<m�ٜ�:���x��Gθ�ޫ³w��a�K4��vm�:ؑ[9/VV�ۣ��]�1s1Q�xޘV�kZ�z�g�77N���R��;�Rqޗ��vL�����j��k��b��e��{v�[ċ
�M`���hY'[��0���w���D����r*�(�b�Y������G3�Y���C;�j�a�p����o1N�EvR]{0�㋥��v��!}��
�wV�^��L�A�v�-��'x�#�����`�Z�I��ҹ��i��V�5�u<Lw�#z��T[���lX�k�K3n%�alX뼻�f��>��U�
��C*����[4�r��.�_\6�vK�9�d��,��',�V���hES[w!�6�̲z�0w�+r�c��h7O4ws5զ�Ỳ��̢	`Zv&&�:���oR�c���S[�����a�(�>�rj�<���Yh��q�p�%���ɯ�����}�i�۩PU�V����+��}��}�����Z%,P+p%wk2�J/?���]�]0�'��7�ct�n��z�f1' \i�Φ�Hغ��[J��I&b�����|�Mn���w/1�Y��,@C��%R���(���;O�]�ʳ/i��~�\�<��	�ScQ{c�9]J-�%e6+3�G�7p=��#69�Q�ۇ/�la��-�9l�2����E:� ��S��܊�=N��F�2��Y�>sNYy��\�F�$?R��x��!Ƈ�+v��xcfL��F��qF��7n��{춹G	ճY/��\�-{����D��Z}q���ܣ�nU�����!z��̳�<�l��T��A�C}��:��Z�i��i_9ϥ�Ѥ3*3����S�}���˥�����2�y�SjkP�˼%�����ҽvE }^͋.���/�/�]�w�hv����ސ�.�V��M�v�̒�`�ۿ{*ƭ}eYJ����J]gs;r�JLւ,a�fWn���f$�d_��S�{A��~���\�UR��\SU]R�]*��UUUUUT�,ڥ햪�Z�ڥ61*�M]R�ڪ����5UUUUUUmUn�������9RF�$�����I;���F�II#}$o������K}$�����7�H�I�#}$o��>��H�I�#}$o����7�F_A�#}$�����7�F�II#�rF�I�<ߤ��]vf��������-UUWUUUUR���*�UU@N�����ڬ�5UUUUT�ԫ\���UUUUUm�JKUUUR��9��UmUUT�UUUUUUU*�UT�UUUUUUUUUU�U*��Z��%���������*�������ʵUUUUUUUUUUUUUUUUUV�UUKE��e�V�����������������ꪪ����������Z���j�����e���j�V�\µuU[UUUU@UUT璪���V����Bj���mQt\�UUW]�}���Q\V��ꪪ���ճUS���jڪ�SU�U�UUU*԰:*������m�;Ȝ%��'n��u��+���Oa0�b짍���{Y]��7,]d�X�{u�Z�ݧջ gc�(�7)n�ou�wf�ݷv�kc��.��1��r�8����s�k#�:�w�R3iT�*��s6*�c*��CH�GD��Z	{�*��&F�I$��A�+��3�4mYA�ꑶR��D�TE��}���r<��6�#I�0��G�^�&���5�*fPi��K'�G��d�-�h;7�g�/bņ��N�uW����*���⪝��2o,�Ęv��>��$�zh�[g㢮��k,c�v1w��h8*A�����	�wqmQ����O-U!�Y�3Z��H���y��XZdc�C�a�e1B�ޡ��y�F��z�V2��NS	KJ
�Z���[��Cp뤬ZA,b�S�G�-�'�<)]�6��d6B�xÔ6��f���s�r8k�,�h7w*�D0�*�ȃE/�bU_�R���e���mڈ�7�ۣ[�@U�-<:2�c��\Gn�x\�L[����FΝm��ﵾF��wb9�����7<�]�֙���l]����P§��tˠ���.�hݝț�e��Ҝ��]Kɶ���Ɔ:7sDQث�ػ��*�ۛ����nN�v�;�-����t/����v��)�]���\��n���@��jz���~}����g�G�<e�p�w�#OnۄM<�g�K�פ���q��ނ�#��\��q���ܴ�^�n�Mj�& ���IǛ]^_!��dᡲ�tl�|<��s5	�(�/82��V\F���pCdς�۴�-���c�<>����Ӹ"3wcb�1���]������n���q�.μ��c'\9{Ei�Ʒ/*=۷x�݇9b��|���ٔ9<�v��ָ0[ZsFi��+Dm7m�����,�V|��Ө� ����ֶ�)5�C�3*��q�	[X���w��/Y���j�z:蓗r�y �{u��9=˞U'vk�r�6�u��D���-c���76N�5�9�C��}�w'9���pɡ�?��-�kv3.x�Wi�pe5tr���e
L��!�[��߿��P>��NW�����Yv�vq�:�,P-B-Tj(V	�{qcԋB��~��kƩe1�F�n79��4�[�csn���|��Q�AIDP��UX�p���n3���t�n{&�lmn�n�Jt�[/�-���ϱ��t�Zφ�����q�uv�ݺCƞ��c���'��H��)s��wFz÷�\����6�Qȼu���
|p}�r���Hcm��W����ߗ?��~-�������ڨ.���3@݋Xa�6�6���D�rs5�(!�m������hP�\�J��x,�	�s��L��P�B�̳�d�K"��Uv�J�Q���ɕ���z���G&����%��6\֞.N/M����8���Fո�[s�x8���{n��0v^�8�L��S=���2^L\X��ʹP��J�'Н��R�.�I�'�)8��p#cgg�9:;8��	#��om����`��ۙ^����8�h鈗=��7�pF^�ڜ��b�e�;T$ݷ2v:9��}������	�k�<��m=p��H�ni�Y�z4�V㭫��e���j㢻)�����Xֱuh��V��Y�3����!�>2޳��m̺\�<��3Ă2^��8��p��I���'�&X<��m�;k�R��Ǟ{v��Y�ޯt��&�X��f�\N�f��m��x��=��u���r���<�6=s�k��]=�����rۮj�h���';}��ݻ |n%:�C�v:.,sf�z�v.�P�Oya�t��r�BX�v��m�8KS��c����{�˹�ɴ'\��ۛ���&�:u�i1�����C�t��nQΪ�yGq�����NEN	�9�J�Rv��*���ݗ��v�V����Ol���۶��\nfCGn�]���v8;�u�\Б����1�O\�s� .����K�u�@�n��n-�7��Z�����|��[��cMm(6�c����AΪ⋭F�la���۞�r�l��M'�P�bz�ltb���l^��n�G3Ő:GXגN��ۦ�N�.�m[��ru�x�O��wg��[�ש��k0��=/vɥ��R�v���uOlu:|v���n.��,�nw.�O^��r��g��j�&��컮��m�T����m�,~}��n4v�wԅzڃkڽ���	��o@��=6����%�m�0��\�/���h�滷�EmqK�Z��/1�������_,p��퍻m�:nt<�m;qݞ���yύr͝�n���/]\�Kq�1`���펺���GL�����׶���X��ۚ}M/g�"sǈ�I��Gb�Ӣ��D����PQ���j�&�:Q�\<��Ls�u��;���m!s��$v��oY�`�v|s<rՔ�W8�/��8�=�ub��}i3���*��WI��4�t9l\j97[9\�C�/b6�F��&��z���l7��h� �嗢��9_�.J�[���F���`wmM��[��M�z��#�񞶚�n��n��p\�p\Mz۵�32�=�mb���v���kWt�l݆/��U��\p���5i7nm��S4��=������o>��ɜ�]v�a��`:��k�f�+Ѻ�g��q�C؞� N�c��a�G�/�`x^ی�MU$��Ւ����Ӳ�w'u�@V�u�b{kv�%jF�Vxݻd�Rlu�B���'�#�tc��2]�on�\^�f�������9��G�U�9�Y�sN;Zۆ�1H��Wc����)13 �pls�5Ҳc�m��jz��Y۬l�uhC�(-γ�i�ƽ/k��v�k���%�y�NT���Gu�m�yvB��x�E�Gg���Xc���:<��ם���ݎ�[�]��eNuWOF�r�(Ӛ�<�+B�����{tGC//z��:S�����ރ��,��nۈ�2��k����^.��{���-c���X�#c�\ㆃ��ϵc�U���哒��+��;��5`�9���)Q�F�*�PvXCl�_Zk>�[m��Q&1v6NŸ�M��v�q����q�������(���{5�Ƚ�]�0[�����x�{�G7�ɽ������x�!A�,���q� �sˬ��ك���1vކOg�����
-�0z|mu�s˱�A�q�L�����4i8{:��v�봹�m;.7>Y=��}�52�-p���y,<�ۃ����j�wkaNd{l�Վ1=*{������Y�t1����kWf�ƕ,ٞ�:y�Z{8ɸ6��р��N|���}���ͽh�mS���gGf�<gs�J���m%�<:��l�/l����gNvrhw%b�v��a㶹�n��%�Ƹ8��d�n���ot]X8��,�7&A�:����;�4]�հ�m�f��v��u�!�K�ݲ�/F�����y����j��i�c��g� '=��բ��<��lvx���,�F]�ݗ�k���\2=�n�3�#Ɲ�[=����13���������vy�SA�F�ݕ��e����v�*���t'5�m��pl�(�8��p�R!�QZe���Y3�[��p1stqS]��-�,0���囐����3�ny㲝���:�n����:�����l/�ďI�V�lm�^ws�Rq�Ճg�.���l���l�K=b�v�m����Ken�9�9�ӌ��p6n�x���1�BCn˒��Ŏ{r�3v����O�qp'��kG�Ң�q5��۝��|<8��ض�L������qw%I�F]�޸r����ϺH��Wu��ŗ�3����^��nZú,��9í�[�O-��\׮�I����d=��j[^9���;x������c�ٷ%��>�����]���F�Xm�i95�>"ݚ��]Y.u��O\����\�3qa���6˧4g9�GZ:֤X{]��z�{�4ųŴ�t�Lu.���>�6�~۶��Md ����OBX`yw<��w8�ݣ�K�r�k[���r�m�y1.��=�;6�XC�گ��R������d��M����9�&x������wl+�WWn�m���9X��d�ۖ��r����l�2v u�7n�d:�f�SF�z�θ<��F�w���-;�A\䇇���n�bL�ټ��&a �;�]�����Ծ����qۃ���Mg�/`�[���oR�cAç�v.ݫ�RW�VZ{hG9�;o;�Z�]l�T�YU�*�cq89T�l�9�vlB9�ǵ�aո���s���g۱��\���{v��prp����A���Fs��8fnN���ظ��]�k۵�G�WrԎ:���9T<F�7��m[]�kأ=���m�^�mh��jQ�Bn���]��7�'u΍�vWsm����ۍ�%���\5����1�2��7[�&�xw;��6����Z7g���m������p��;q��7M]��6�t�5��qu���\�׋�Gc��C���e�.�	k��7c=��u�Fi��t���pFK��*8�J�⡵���n�m�3s�.������ċ[�����v�g�n��9�.{n����c�ZnF᠎4��֕�X��"3דn���ќ��wk���AX�ܛ����9�l�F��n�W�|��3Զ��V���ɴ��x�Q�ƕ���hVb�guv�Э�8v�n<t�j�'�ݷl�y��n��=�U�\4�Ms��;���������^؝�G����0�c�\W�u�ś��ӱ�\�/Xz�;���^��@vʪ�q˽�)��J琕U�B��Bp�w�����?�]���
�AskwwowF�,�����e��G�6�IJ� �)�.Q������꠲R�UU�AO �UU ���J���UUzUUU�Z�JHL�ͪerU$�Fx�g5��Ho�u��[I���������]����ޠ�fG�����ُB6�	����]�35n��V�jc���<�Y�;�-�W�1����>�ΙLZ�Ͷ놮#͘#��ǭ�x�Kղ���m��6Q��zQs�������x;��I�e�\���z4�J��MȨ���:�դ����n�bX6[d^.8zM��8�C��n��$�ض��q�U!��>�̫���S˅���k��I����O:q�۷���CmrS��Hv�[�r��;�n
��J 
�F7`
YX�[��Z�F�ѫ\<u��8�-q��t9�6��<C�\��a���6��EΡ��#Xj�bk;J��f��\;a��=N�}���;Y롭sF��.��!�p<�x�w]��v��˃&�!^�c� Y�۹m�"��� #�jN�B�t�݃0mx�1<�/Ni�s������ⵁ��W��^r�1a�ɥ���s�ϱb��������`F����w8��b�v�9΃=��{s�	�r�3�y����8���k�W�<�����bk��e�zͩ���f�����b)�m���c��tn�ރ��n%<�2���y��;��n��9Y�����\[e��[Y���e��۔;mݸ
�tE�-h��V��w<P�4V�\!�M=y�>��v��n$�R��Hu��29�zP&�Ӆ�=���\뗞{'�]���-��#��q×YI(=q3ǲ�p��.��'�=iɵZ;W��]��X�v���7
`*�͹8�4��5����2n�u���=�jz6���-�v����1[u���&}�F���v�v�6�6�=K�6�n��d��E
�KȧP��e��nw�Wi�n4�܃��vWb�I�ʃҞ,LK�nn��j�a�{Y���t���Ob������!���}uu�w��c	cX�ε5%mrS5@�I�m���Ѫ�^��q�[td5���_��^�.�ӻqX�Kvݏ7b��\j���9�ֺ+"g�k���E�/nݛmK��v��<kRuk�;<�ً���lF���N�\�]�[��n�[���m�)�g�w:z����	c�Е�֮w`9�x4#�넎c����m�{ncԥ�Q�q��X=��l�t�۰<��vpm��y���nS��n��=��ژj(0q��I2���|�~��0�nm�8g���[LNʻ�w
�V�Weؼ.�-�ptQ(�-����n���{��B�`@���D{���H���K^�oCP��U���g[vǹ��xhF���	HG#�\��eI����}f{�����Tݭ��b9uX�c��{�������}�I5ȃ
[p��5R�oN��=;GS��9��f�~u��]�������`�V|=2�f�y�V�z���h)F���8*��J�\��\{uPqɧ|�_�>&���W�t�T�D���ü�͏���:h�P�B��T�U#�K1ϯ7A8���O$kv|��8B1�n�I���C 2d��qwG�;�eq>�y,K��M_S=*�g��t���/o�v��)��H�R���]�+u��k[b�\:�^�Ҭ���V�M��v��ַ!z.,^����ۋ^��^�Xz��-�s6�Z"��tB-�;d?V���;���-�c]wC��5�����]j�qڌ���%i�s�v\D��o�\�{���g�UU��ntwXy�Gn/"d��59�;p�p7�!M��(� qF�)]A'Q���*r��Xj�yһ��u;��M,ee�3=l��驫/��߭�y�d0������n��O�.��[��,�k�϶]a��p�y��XX�n�����%ZX���!*t�[��A��Ӷ��������6�l/msF5ŭʒ�lY�Q&�ў����#{b��}���w�>�J}ǧb��"�9c��̱`��s��x*!N�M@\F�N~JCw
MVI��K.d�_���ܾd'����o{����jC�˙�F���p�scM�UNi�e���@�?8�`k'&�s�T�P\���ܧ������wj׾�"� 0V^*#~`��b����9��k;�߄� s՘��Zme�S�
�\q�io���+wu�6�%:�a�+�w��ҡ����q>N�Y���/1d�MD��rH�*O��%g�;&��pɕ��0qz!���0��W��.m��~�<�a,Op�\�
F���эHo,�S�VYR�-���iI��ɛ��4�f�V	��Sy�2<��go,Z���1�
M�D�l�l�����v���5���E���]r۳\��$P �H���;;g=��JXQ��_-���3k���t�ߣBW{�jC2�N�fU>F�S�A��N6��ֱ!��|qS�}}|;w��۴�ݒ0�i��h���\1K�Y�S�n�}�a��i��%�Lq۵���u���/S���{V�,;p�㎎�����=�}�;j�x�a��Ӽ�i!��*H�_=���(#����͛λ��C޿��k
�^�G	�����+���Vj�5_'�ЅY�5�Ae]��)�7B�;�.UY:J��ۡ���CH[b��Rw(�/.[-f��3��Q��\�O���%5-H���ԝ�ݗQ���imj��j����r��]�����v�UoK���+�R�8PbD��_i�]����8�;�T.�Z��I��E�.��[�c	U/u��u�����gb7��q�gyݐ�j�
M>��/���p�uZ�u���hR�`���Ra��ڽ��=����m#�^]��b��Y�|�d�9󰌖���f�V����L����R�������I3	K���[�'�;_^�1U����\�6�Ӳ���N��5$��~Y��D�~y���e��
�kO�"�&�-N��Z:�4�y�Z�XN󰧇�a�����<m�_�Bb������w,�)$��'�z��`�F�.��Vd�씬�3���dv(L��3�=׮F��sҏY��9�%0��Hi�\�[��	Ԁ�VQr3���Y[���JЙj���![vl)���܍��a�X��vT�e��fWں�Y� Ch"lV��5UUt���ݼL���q���l@�<{qM�năt\����rs���ۂְƻ6�c�ݹ���Y�+��"��	v[����lp���.�:qX(�_�/����Vݺ�G�]��ൣh���K*SR�,�RC�19'5psn.�j�j��f�.t�4���)�歰��c�o;}�p�Y��vg[qK�9�E��l��i�	��j麞ͳRb2"ۏ_ˣ]�X��ap���*�Ӛ=s�:�
P�Q�i�����=�6��c�'"�����r�b�O�vo�h���+|-��?O5:��r�w\����7SݾflJ�ѐ�����q[!?�7��{
��7��+���c�KG�{g���=ҡ`<����VC�C����9��[��N~���kp��o�Y���z_#3��賚��5���S�{�V��|V�9�f��e\���KJOY<28�#���>U]�ֆku���}3ˣV��2�����^�3��z|�cɤ����]�s釴c�8���y1u�EnsW�q�O���]@ge�w8�gkfv��e:�k�v�?g�9j4Ӄ˰K��[�i$�u�ˮ-پ�]s���������k��&�[��&�$��8 �H�7i�7zv��^�?�����S�z6�4�&�mf��m��f��Ţf)@w7}C��Y�p���i���P�}%z�%��o��6>L�~��{��.ǂ�}<������O��K�����5B�Я�BE%[
"#q���?:��T�-�ޝʻQ�̥u����{r��No�V_�6�{3z�M���,(H.��tyf߮�JUP��B�ؤ���%Tf��+�X�<�MR�^�Ħ��5�C�ʄ�r��ȷ��m߻nPXB~t8��]	�&��7�CCG�'/[���$���W��Z 3�W/>��Wc�ͺq��n�s� l�qD�筶q͹N3' ��\H�ш��ֹ������/u_^�ժ�ʻ⪯�צ��ߺp�Ww)��N�>%q�Ab�]��Ly�Мj����J�**�z|�
�{\�k堏���^n�匽7���\�����Bģ!���Ww:9���9;v�t`��,a����K�t׶ ��?W ���(<��%�6���M�|�MպU�G�oc��e�$Lu0{Q����2�;=���i��Ar�_f^#��<�z�%m�ӎ70��ř9ޣ�j�L|�¨�A�uKF��+"�U����n��6�_7�������(���d��nzy��\�m�99�z��	ݓ���_�^���E�oi�����$��
�"��>��']��o����ۭ��9xz,�Aݪ"]�{hN���6ūͯMp��c�ti�S���&�P4��x{��72T�Ŋ��篴Ko��Z<�vW�jY�xce�%Da�(Jn*�� �	�'G�u��&����S�B������0m�٫B�S֜�\�k*�{fb�r^SJσ�a�H��I��p�4��[���N��;�t��W{{����ѣ��@�8�}�,pÐ0��E!�yU�o#��{Kj�v�ntǰ=����x����h*��ut|�h��
v�q_h�L\ލ��wqo���{�y�Qg��"�[h{<��U݊w����c	Q:�_<q\��m�K����^�I7�m��BL-9�9\sy%����c��7�������UO{���͍�3��x�^"�~kc�"�Z�1h���}����[�ǣ����t�f���W+�>6n�e��5G��Z�/w�q��7��ǹD*����k(O�+|�7W�����.�q>��-pF8�MӃ1KG�qC�J�)m�î>{�U�?k�^�DU@�Z�����Y�TUa� yWKlӍ&#� �9/��R�	nuC�c�zs�v�.=V3+��זq�wU���KWBID\dG5-<3sI�|;r��,�V�6�����#�R	u7�����o�U���(��zύ"�.��$�!OA{���[���Y+%�-��#����W,c��x�x/L�9���_K�nG�VX��y�t���Wh�.];)�ca��7��vޥ@�w9ieY�s�(�M�����蛄�P��7��w�����m�.ZV��mU秃'�U�{���7 o�y��6�+�8�t����}�[q�-jh8�8
���z''c����a�]�<�V��;�=������ݱs�8�8�w:97g�n�f|\>�q���uq���\s�:�5�=�GW�n�6Ǎ���ogf��m�m�[�N�;��t'��z�j�<Ճ�sq�i��������W���\��ɠ���)�9Bz3���2�+��	��HӦκ�5�x����5�z9�e�\u�np/Sp=����]}��Vʬ���zp�`��T~�>y��\(������43�������f@����p�o��K�}��w�5��gK�R� ��_�M�<����9��+#�����jm���?~�������.�e}YU���f-���+���:K���0�{(r����k����'P��Q��U�Ε^ܻ�����}�"d}�-��L�:�<�܏�]��ށ��T����{����9�I2H����%�K��D��'.�>����"=��W���"Vm��|��'���ck��?c��[h���1c�	���uqM�����=H���T닖��H��d�[(H\���f{�;t<;+�Nv3ƈ����{#<Fv[�h�lgc��p�E�w��.J�b��M8��_2cy�H�L������0�(�QX���Z��-��(?�	[F<�$S��ۜ���A���[)�%vlX��h������4�1��n�>ߢ�4��������o��{Je�K��y.��RP�H�m���}Ӎ����ڶ�m�݃o	�8�:����c/D���E�_ԕ�7p�Tb
.D����v��}�w�}5o����)Awb���n���갂��nW�ԉV:L
m!Hs*��3�����.gx�3���]^ڙُ���Swoi��͋��NsY��&�^�ĸA|��]qnW�2۱�;������Il�����᠉��)@�Q�\"Bl��I�^=~}h�7�����Q�T��Zy3�b�ܐ��mx��!	�^
	��qȫ?~�Msg���SJk/:5u��J9'<��ux����)[I4m�r�����q����.Cg��o��ê�T�dPy��m�3k�҆�hʣ�4�QZ�ÛEQ/������(fԫ����G�4Ar������c�����Q�H~Z�f!�ř�
yL��u9[K��%K�#������ehZ:�a:�;�=�2:�Z�V��h�t���TVߛ5�^�k�U<�D+�i�q���؀��\�c�7�ʼb���P���`W�D�p�n
�9��7�V8ft��<���wpt%��`[��f���D����yP��d�.�m��ڻ���,�9*�nv��e#�_oe�_X*���γI�\��u�s���z���"t�Wu�[J�]uq#\Y�kS�mJ����*Ş�C���F�p��oo�,C�,躀��2�͗�H���`Q��#)�X5Ss8�b˫M�Gv��<�
�U�+.g������^ͤ��XJآ5��}s�(�o)��{m�9���U����ؕ����  �l	4ӆ9R޼��lq�Vh��z��]��VͶ�I+:D�Oۣ����	��qu9�4��yS-����1�Y��"XM��j�4�k��jk������V����/x�i锦�ʕ4NDi*'�7C�<�-R����Z���oS5^DB��s�]H�aW1z��L�8�,a���o��IMׅA�B��]�!Ź[��j���`>�j�F�?���%�p�ejvjpu�F����+��WQǤw;�V�Sq3bT0#�#@�vfl�}X{�t��$m���z/J�B�,�M�v�p�������!���^��tl�T��F�oD�C�0F�F0���v�_D\���G�4�ȉ����S����]W@Q��������ږ���|W�t�%{�s����q�
�v��n�>�/�8K4@��4т1�Z���K԰ɜ��CB�xY=o��| �}V���'����~��$��3�9���#8���9!�x�H��Pç�������kjy�B�qm�����<����8��ҭ��mЧ6�3�N������0��AT�ή�/�+Zb�~>�v+�:��P�b���	�!�$���TG����T�Ъ{�Q�#du��r���0�� ����F8[B�Rۉ���I��Ww����z#щ�k�����"{�d2�f�ů�� P�_UЀ���V���s��6lU��fӋhv�S��9j΄�l�Qd������sR�Hd#��*��je�������4����]dPӤ20��,Pȫ��~��4��XI�EUu�9t�����5����4�<�4�t�iC�Q���
����H��#:k��?Y��i(�*Ոp���|6Eee7i�)�)��O���e#:�l�zr�#�Nfmm]!���@��FU��ʡl!_�!g���O���Y<�橊zٔ N��nm�!�$m�ڼ4VA��vJ8s���B��̑�&U�WV��H�`���dA�_Q�)�L���GԨ��s�yw�̝�ƞ�Ԁ�n*���26�^� ujKqm�Z��pZ�kd��:�9f�c+�0��h&LC��d(��_-ھ5G����/��9�L"�|���9SɆ����v7�f�?"=U�a��N}����|��*���6�%�)sD@-�(�{����S-LT���(f_]�_�?)Sy@��w^��H�!�E����We.'���D��&k4x�\(B�fږ��Lq�q�C���Y[r5�;=$��3�ΓY��M{�8�''��eۑ�D���H[�#�i�/�6/�[��1��EZ��l�YC�QR��<���\���s1B~��]�Һ*h�k�g�2����1Lw��<�D�1�nGm�i̦0���f����u�Xk$�g�5��1�/�S�,�"5��q����'�i��~�����H'H'`��g� d���0ı3�me&c�1�pK��Ɍc���΋C��uP��w��f ���D�\�q�{f���э>�����-�i�����W�A�����n��v�+�?T�ߦ��\�5�j����٠�`]�}����v��|A���[e�"��؍ۦ;g��>u�ٽ�!�kgun{5�����B�9�\�a�%���Q3�F�B�ىV�ny˩P��䏉sI\ۨ��&�����J���zHV����t���n�an9nt+{Z���]&ڳQQ����@m����Y�tc�q��gf���s�`�o:ck۷c,�7U;�i��j���.����J��x�{X�o������9�[��ah����c
�� ���1�Qa]5���ԒБ�k
��t�ᅄŅ�>�ʢX��L_a$cTX�g~�2����W�}��s+�0��C���g{�.p��>0���bKB�ҿ��i�		p��^[�(�H��|>�8�u��H��?
���!�G�u�a|ac}xǌa3Yi�ƽ�eg�4$�JLcb��,pB\�>��apXY���bJ��;�j�m>�pH��.���w���|5�j��U(��vWe�H�r*BG]��Qu�}��&p��<�D�޻sgZ�
���2���#�A�u�~�3r��|t�J�>��ͽ?(�cB�Z[�O;brZVEc�ip}r��o��^ç���@t�!z�}>_����`����G�WL�WeI2�5K�7��P�FN�9��\Q�2��r{>��$�Ga��G%�j��4l�/�6G�L��E������l]�_u�Nr+��~�ޮ3����Wt���Tg܀%Ndt�P<,W�~����v��6��,�և��8k7��!Ю;��^:�cI������{W�a&�Ӿ�}��#GN�S�L�������2x��z$Y�d|<%T���}=n��u˲)�V�����$ɇ]��������g��4�v��̭%�� C!�y�<o�+��+f�d1]8�Dyj���pZ�כ>��Q���A����zf�k���M��:(���)�,0�ܽ�볩�5{�X���[24�<���\�K4�����Hx�hx��ڊ�6~NlIo"�h��=�"%�Ж7Kl�:o�	�ԫ�-�2���|~�>������n�H$k�Vjc�a����������#ƞ��C�@z�b�,�]w���r8$�4ۇ?����6��My�'���?x4���$Q�mxb���8��<p�F	�p��:*���׮����?IF��<���F�ʂ���;֕9�����)���c�L�A�XR�k�;g��3�(�8�|IFN�:z��T,@E�b��6F�\E��:Уͳ�?���sςq(h�.(�)%��m���V�'p��*��t�i뉌���<]���F��D�r>Qz0H7��������@��w�܍ {Ҿ?|"bOϪD���KўrE���x�VWD��* DI�h�uU)J:�H6x���k"�ϽfG�8��e%����Gg��G�Fr�4�(�j�B����#�w�Y`��i���S���:l�<6���)�"���Im���_@m�B���2�2p�(�$r���ӎ=F���R)�~n��g�w"ceL���,;��ۀ�i�-KWTY��-tM{5�v�n�_ݳ,SA��͋��b��f���S�H���qà:��4( xs�[�MoFV5SL@G�s�x��W!YB10ؠI��#ѷY�9�ς�;�x�?Q@�6^�O�k�ML�|����r) #�dP{�p+$�?3e����u�.������e3N��j�WI$�+�� ]y�d9���I��Y�n�$����	��2�̍?Y����/�5���� ��� r��D�܌O���m��v����c(��|���<X�r��F�u����l��m-�x��$�^���tn��ь��Tݤ���g@��>2����r��j���ƅ��o8�2�G�h��tP�0s�qI_̅K�J�}ՆQ<Y����~5�¢Z�DJ�e�\F0�(a�(�:�آM���FD,�7�">�@qꑪ��#肇D�č���0�bJ�]u��(*��h��"<3ɵ��~\c 7�rܥ�>��ϔ`�H�uQ"��[d�&Q^���R,��<��2���!�A���}����"%H�̾��1}�UE�T`��ᨲ#�#��D+�׭�M�=����ηäd�^�T���A�"�+��Y��j�"�`�u�_c��8Ck��#/��}�q)^�"���o;Q�AXruv�����<�7> uJ;> ����%.�c8bIf:!V,
ೡCOq��:�f�w����֥8`4)�ޞd��,�	���x�?�,���L�d;Pe/���\��ٌ��b<��V���$�wZ�����,���%�̐b��%�a/ۿ.�
��~��.l�M�ʉ\��'fsa\�B�WYޱW�P�8^G�,��f������K�d>·����V~x��QE�����`ɂ��!w{�#��|w9���0��x�=kۣ?H�7�EN�Y���']�H�2g9�tF���U���EX^�_x�eeM��
�>�3����ǅϳ �q����{��Zb�r�ΓzG�G �e�~�(���ٍҘ*㱲�,�k�]��"3�}��8��0����������7�aj���B'�w�aF�D7[�w����fd}%�ш��d�	m������k!>���� �|���q�$\/�V���?SGv��C�u=�"� ��v��ᇸ��4��4�G��4�Ȃ����l�KT*����>dYUx�T�쿬�}0O��!DGw��FpI�j��"���-Q
"{�N|G�F4/n>������B�}�OSNm�Z~�������6<A8��fA���9���SU�����q���t�t �9�.�U��vi$
]�U��N�-Ka�rF��Im$�n��m���N�aY���2'`5���g�	��y���f��Mc9i�)S"%B$"tTRE8�tn����ۧ��'g���v�v�WCpn�e�ްt97>�xNָ�y�Zq�m���p+W.|�g��Y\��F�j�g�n˶.8駗tu�+�۞����\/��׍��ϰ�p�T������e����ӓ�&QGk����v���g�gJ��x8�l��l�u���4p!-Q����Q�3�!�ɻ9V5k)�K��~MxLA������5iȈfR���ܤx��x��@��R;;��N7�p9�H~SK���h*Yd����A�1�pF�H�#L9�>"�0Qrs��}�(���um��#�y>#f�9�q����i����K�b���Q��θ����֍�ጏm{y�aT}�R�+t�٠]:~�I]Uʀ�(��_O����b�;�2��{�����;���e�g��ur�F�7��Aj<C��ս�UX���j�[w�/\A�U�s)�?G^
�7����{b�F@d�uS����1&"M����j��"0�!j��>#�7��G˾RR�z� �VDW[���㱨��m���R��'��1<���6I�X|F�ٰ�4��I����~ç�=yER���nEj�He�>���Hr�8L� f(`������߻�n9c�%���^S�umקY��0��H&�vػv�O�u6Ţ[��
���d��T@�BȻ�������$@ʀN���*E� ��������<����"n�g4DF�4�Q9�>$��v�����{��0� ۴r[t�p�x\��`���������q�/[�)����S�e�8QWCf��g���-�l2k��Ñ�Ż�g��_�m���Z<A���Od�|��xEg���ב"q}4�(ѳݷ�jF�^@�"L�,�^�H�Y�H�0(���W��<a�}�F5��Z@m��E�L��C�8os:�\��~�kk�C�"��FX_T�[�����p(�t�����A��Ŷ�.�4g������|D�$��$i���ҋ[w|dY���"9�Z���`�#+}ܯ�؎�w��9��Cc��/��"y�l0�D�T�ו�6���������M��aH�0<v!�@�%u0����9(qB��B3��p��{bI�G�#��lZ.^?��hx����Sb���y>�|[��n.@�n�,�sܹ��+���Y��=�sX����k�W77:3�U�ۿ{O�B�$���딏�S��'��Y�~aR�C"�!���"2_JW.���oS1'�[d[��$�Ab��
,������'<V�C�U�[����0Idt�p��xi v�kf^vq�6�d�s�"��e OĻ�3]�NB��a��!�w7ޙ[0�A�r�vN�;Шm�s>ύ�F�� �+��jɣ�u�pLǍIu�=��h^"�]u����p���Żxy;V�}����Y�����d!�.�\�W���l�5�r@9Eu�S3�Va/�*�/M����+��.ML���0�=���: ��� �A�l�|�x�?x�@5o�[i�rJ�b��Y�P�D���e�.�ԥt��Db���~���)kD����C��mT,,��@;���" �L����\�D���M�z���	�_��ZϚ�\RW)]q��5�q��
$�;��S-�Q�4o�:�y/?t��O������GOD��@�8�Lg /_����8��-.�4k�p���x���̄E$�����#u��uϷ5bbv���&!�۷ ��A����E+Mu�8�l�	���C-l[7�n�g#A��#�M��PE���Q���7�@�yJ�#H$2.6
^u����N4gR��?hהhq� ���%�Z(A�4j�"U��J���^^����4�V�`b���?-C���u=�2�{��G������$!����������bxS��c��V�-��,�+��H�F�6�'a�}�a��T$L�������2xViڽ�X��(v�����Y�_k�+f,X�������TȌ%�h|�����m�5L1^�����^���9i���h�����!��ѦM�C�>R6������c+�/n'xt�]�s�^�KX���J��=s���X��)�J�[�7U�*O�-�wOm��=�4���ٙs(�KA'�WU�Ȝ��؝�"\!ԇ��p�D=��v�X��;F�%�8WN�#xȻ��Pt���E�Ok�pU5�ӯ���YV���}ƾ�G��0�~�s�6x�e$�h]�=�����F�Iƛm-XM�y�=���K�۫չ!���MJ�Rb�´�N�;��̷5�
a�҂��y]�x�"��>����?3� �2���hz�j�Hbs;[� ��iW*��@�a��Bo�|J
�M05��Y��-������x��n��$����E�B?N�-����:I4r>=�Ğ�"�p��\n)��A�E��O���Ƈ�_y�Z"@Jl��K3�0���,�k�{�ц�@��
��v}a�".{xxY_�[�֔!���<�	�pQD�<����~7Ӈ ȜO�G��ZF{ө���""Ul�d4 O-�9�߻�O�,��
*�ݽ�1勝]�A/�-�9�#����I����x�F���uy�Vf.�攑���OȢ�j��#�\@\��4�AQ��$ۡfϒ[4�$A)�~&������>TM-������!	Y�W����I?�ҹQm�T�����N����X��a!}�EgH��M?�acPA(��]�����wV�&���K)C��������FZHH�l/�$6����g��M]g�w��'*�I��A�G71���=`T)��%}�w�n������V�w�yD7؝��Srj��-���'���˙���4p�9��R,kz�}Պ��m`ܗ7��y��)zwE����Z�0�_ �������Z5oG�»0k�L�w����׈�&mj(�c��s���`�+���v�L��З���v֟��w-a��uwc-�j�TlSBAJD))�P>a�d�V�{V�^�)#I�Dr��7��EV�刞�]����Q��֭6�Z��1ƪ6}��#E��7�l��-:$VM^��u�W֗r5���Sǹ�N7B�*L<|�e�-V���̆�1Z2�҂]��xn��X�PO8��-uɜ�Z�{��0�Qt���/����Ԭk[Gi��`��V^�U|T�͛��'N�Vj���79��Ъ�ǎ��e��ry�e�F1��0Z4��Zˎ�,���c]�]ս���6R\Z�BU�.�gQ����Yn�aS%3n�{��V�;z>�5��,� m�7�}��//X/�u�m�� +՗#F����jӴ��D�;�$��[�g^��X�D�R�N;s�Ef���fK���m��=>v/��
��"�޴�<�ګ2Mz���Ү�
$AT�=�PUt:;�ٙ���j���.j�S��:�ŕ�<)�߄^A&�m��m2���$&I$�l������}���{߿��������,�ZJ&V	�U�H��UUUOlT�uUUUU*�O2�*Ҽ�KU���T�Wʢ�mr�QE<�;0���n�λv�x�ێ8�-Ӛˁ?u@���i��,Pb�Aď���3�Ia��c�����w׸a�Yci�����r	%�,�Xy)��(3~v�1� <o���;�}��5�j���jS�v�'k\fNL\�u|��v��J�h�6����;t�y��2\�6͡b5���x��P������8��4�
�kd7k�g��s�v��g�[e������v��딸��7�p�p���eit5��y.ΓW<ܳ�;l:ݸ�p��������:纅�+�j�i�M�us�aؕ�{k[:{lk���	6�;s����s��z�����u�{cz��-��)�x���n�]�C�F���7a�6v�<v�9���+���IS��g�۝���Sۋ����#�ԗ\yL�t�A�!y�Gl�:��.b֝��x�j[a���u�,';��'��sPu۷��.��3��м��r�����m=����`��2{%30�����a�.x��3P��,I�X5�n�]��ۤe�{g�$�=��Z�һe�����eýUϱ�׷����p�ΛY��i����sO��u�&;'K���MC֫��Ì3u;,�=*�7=m^�Fynm<�.�p�v��c��j0鹩�N���hF������z�5݅��hS�v����jJ�����C�;��.LG��n��]��bN�u. x�\X:��;�����U�v*��X9$�ݡ���lԜcO8��g��&�˶�i��
�a�����Q����0�q&�-��h����[��E��6�f|��p	#��O[���c�qq�ה�*u�ظ�}׮�h��{u�6��Z�v���9��c���T�ٞ�gj� a�bXE{;a�U���q���$��f�n^3��GvM���r�\��um=)��Rv�7n��:�rpn"���3պ����Mn�����vB��H�?TqS	��jڦK��v�)2O�t���.��η9����Yc`hO.�DU\td��YV1c�(���wnv�{�w��5���ڝs��(���7X�cm��*VNc;ؼ;�v.�%�n]ƹ�k���(��QV�&�&�F!B��7f�N6�w���k�+��F�=Q)�gm�$v�ù�mWg:I�XM�����Uj�p��d;-ɒ^���y�l���=5��<������\�.�yw^�ح��I���ո{�ˬ9���8��v.e��o��{-Rڍ��t���{��6w���1�]�i�%RD�;r6���%�[�������ɬ����b����Z�BD���c�6)���`+j����%���Tv�ƃܐ�w�K^����|���f`�
^�W�2�M�Xa�O��U���XQe�h"9Vr�5�&� ��$�U z���Lޥ�{E�ߝ��������y��kr�P�Ue����8ך���E//�w�ykJ� �A{���5QB���(*���B���������}e�H�AhPb�54I�\�V6�U�T�"�	<9Sk���m�j�~N�e|{�󋜙� �*��G0�A��?Uo+7�P �}?Cih9���v7�#) ͵�*�C2���� ��H(�Ew)�Gp� �f�M=Α��O�F&�E��7�y�zQ�c��,�Z���m���6S-�����Ka��*3zԡ�Qoמ�7|��O�4>H�X�0����DR��g��(~$j�Z��lXW� �G�{[5��T%�'(�~���q�Vb19j����*�9;Es�CX�mA6�w/l�84���ul���h��O�M���e��j���C ���H�=�_��<[H�mb�D��fQ��7��� �zdf�AD ��ڞ��ᥰB7��*� �4G1>�׷�9Ymx��7v� c-�|g��$?D�t��2�^H�~C����3���F�;��jdK��Я3c���"N�g�jiw�CY�Ii���c]�d(nT� ��uyp�F[�4��e��'�A!K���j��� ��D*����tH��@ �����2�F;z��e�%Ua���?Z�UH��h,���), 9v�Ň� �R�
�������� �9Z���F��|f���bG�{�Z���7v<��V]�/[�M{���f�#a���U�M�2:��7���z�3�=i�h��m��^(�(R�Q�~/8�,�L9W{*�
"
8�2����rI��fG�$!kY���d{�'�&s��{��&��u�"�����1�2)}�>�����UBZik[�ە�c�E���Of�����y��ئ���},���n'X�I-)�Xj�8������P�L�)�1�C�߽��䛰i���>H�����	�E�j���Ғn!�.
�7\lj:ܮ-'Ѷ���=73'e�;P\���n�h�Ѯ���IW�o�{e?Q�������v�G��M����˨;��pp��Q�J[3�uƨ�l���|M�p�!����ލq�{n�"�ۙP�{���D����̵p6e�n��(�>{��T��V���	;H2�}��c��!����bЙ��{w&��ـ�\+�#n����zņ��(������,�)@$��H�a&��'%dXfqL+l3e�Nί��\�?�|�4W��
K�|,w�b�Vk���.��Ż���:�����ifq�С�M~��jw�͹	��<�c�Vj+�Mմ��e_�w��>Q�}ޫ�e��	\������{״���󑶄�m�s��~�U���9H���s� _��y��3���,�7^�c�J?�����d���w�X"��������'�}sAñ���Jb�
s^[T]��T���j������^o��"�����@��1����1�vc&t���g���B������o�Z��t�A�d�D�{ҿR��uY�LHi,�M&L�[��@�ZB�r�E�f�/s�s����Q��,��H�$�nV�pm�vu�޷&q�l]=��r�sV����[#5�-�����L+�����}u�,I���	j�>߷�VG�\Q��*�%��^��|�g*��A�^�d ���֟w0�1�7���.[����J䶸�U�׬��s�}�,�~�V\�A��z}e�Ϙ=��jh�HX�/���fA@���h������F�ϻ?X�m�![x�b$����q�˕�%Rr��^�?a�^���/�|���*;L�����m5ȜqGPz{�gC����V6��'}�?QӍ����R;�Ih!bF&yS6U��LB?A4��7{$ոȀ�������
s���O���P�,6�bť�މ٦ ��e�/w��G�Ӡ��t����L�@�\۾�(�z�J?-D�0�+/��n�ǡ!��*����y�%ߠ�<�퓢�
�Ѳm��4NJ�*P`�nl��(������3�o^��X��ɑB�ㇸc�o�.��v�����>��!t��	�E��Z8�d��GL��F>����x�^8Pm)1��p\�^û��TO�69,��E$amW�\����7џQԈ&n�P�fv d\2D�I'/�[|��# ;�.�|�xu��;���dƶ|oGe1=�\��m�-�0�u��va����z�{�:y�F20m}�<ioO�2< TW���;�B�F/�"�&��t,��bA��,��r�x�N�pe�D8@�N��z�mfu��xa�S�{�>C��4ؑ�_�PD�ҍ��n�g��H��gS��>jk�2Lw��h�F���a�N�ڹ����LƌL�}ʗG�À���̃���I�|�m �5�)l��ev7v��j=.�Pa#��۩p��cAG�uX�g�)�u���9��!�/<�{�>�fug��VL�>�}��� A���g����N�@���v�k �Gc��]s��=˸�O���9�"Z@�@2�f=�?[�c�d(���Z��$�(�H��ň{�L�H��c=�/�e�����xNks�ЮT"����k��@���N��=���m�A#�d�g6���򺧣���A���g�EA#wz���4i#�i�=;�	6��;'hU��`Z��z�|��/��ٯ��k0��BƳA҆��ٮ�^��E�5���M��[D�_+j�=z�e�\�mʒ�����Gp?<��Ě>s�Fۨ�i�$��e嶭�b��"�_��~�<q��o/5�����#�5l���̃;�Jۇ���ϋ���������^���V�;��
&�l�ܢ�*�e�q�Z:���L�j�Lm�J��K�7Q�hkZ��D�w92-�&��oen	�)
3���6;W��{C�nܸ�JW�g��4���]x3�/�5�Ϊ�wE�����(vhV{�r�|n�V��V]�je庮v��\k����%���텶�ޖ3)`��������b	��d8k����^zc�4��@2:���U�kn`�M�Z������Z.ί;�����i� 0YVQ&���U\����A#���}�k"��e�j���[�#$L�7;��
�>5�n�?�~�3�Yr��\4SO9�ݿy�A��HcB}H�)� ���ʭ��$:�oW���g�q�!8�9n�KZDTi�D��D�nqb1@�D�)n}睆6�n&�`"�;�D�����dgBFd>����CiD!U~�G�l�0����;�w(�F؍e��L��ϳ�k��[!!�����h�B��z���U1�AZ6�H(�F��쫢4� E���Hk�u��X���sOu?���ga�)������{����kl���� ��F���ݘ*��6�)$�kb�g�*|'�!�W\˱@a	�H@�&L���7ot�W�k��4�'�?2��B�E��}��6)��{�����1E�N"B��k�{z+��rE�eVF*��zr��9�S�ݺ�Ӌb�.���px��[q;�7<͢��7k�F���l���->�F�.�ܫh]9�a��9ߞtxz����7���[�i�ȴs���vW�;����ow��� �Ԡu�d]?@RN�Z�嵢ۤ�`|sL���l1ъ;�>�,����$���0������:΄]�]�OH�}ى\���wZ9v5EQ�:ٍw^�hVv��a7�߮����.��D��e��:�g5~{�BQ}3>We$Rd�
}R�~���i&��)�{e��+|pg����H:���ilMMM��e4�G���ޙиB�6��	���YkQ�3	G���WY��w"5ڿW�:���5��}Lp���R�i�S*��������7��� �D�l�4_`D�F<0�h�-%�T8��0�\l�H�>��L��(�oYٞ�Ve1�� 0w7P�]�y�b&�u�Vϛ[0��p'��ͷ<���F�0�0Ɓo�HW_�yZ��b�m�6����5�7���`��	&Pʝ�Fz0��#�~��� #GHY��b�(�wg[��,�8�;I~D�8���k�vu(VƠ얷���xH�����V��粲�I2��6�c_tL蔏1���*_Q��|I2V�����J�Ö��8D��˭��-���A2|3�J�#Ȥ�Ɓ���9#�aTP�ۓW��9WZ,�)e��i�	!E�뿾wdi��]{TsNx���н���$�r�KPS/ت��3hA^�y��n�cj��[�Dl�)"��)/��{�Dh�!Gq��c5��H���X�JYft���^&q�TA��n�-�n,֎�(i�އ�(�$���@r+�l_Ĩ����0\�>�@|��O��d��^;Y��t�x��<�^W8/bʰ�m%��ܯ(�]�C�ffN�@3=��A��frҀdh�_{�'Ή0;�ъ���~#��
K]dq���l<��%n�ȝ�9�H!��đ�E�Bm5�uߞWqf3 �;���Ø|�*����~��3~ ��k�6~#�bb�G�]�ע<HA��r]- �ܕe� k�g�:6&dh������g�},o�}3�bχ�d$H�@��]�"�'�C�� �A$���֪��:F��}�0g;z�^S�y�V!�Z�!@u��;1ד��i�z��'�F]�iͷS�#��씌k�2�r�ށ���3(������X�~'q@,��3������H�"a	�ޟ����D����$Y*���M }�t��ն1%h0�||���QY+)]�y6tx��FhB=u�hh������O|t��!�Yg�꟨�A��[������F(��6��%�a��RM䉋�uK�'P~��(�H�2��oC���8d���f�k��4��� ���$Y'
2~+С|� ���@ڳ�R[7|�����<�<���#N�B�4�$�/�U�� �}�I������vYPK\r6�B��Ӡ�H���ſ9�d"\�r�&��2RD(�w|�Y=�����!K���a;��ʳ�G������a����o�<{8��>W9Ŧ\��o�0ݔ����k$T�|eEh��}��B^���jj�ޥ�u��}��Wq������#�J�N-?A-+���G\����-���|{msƏ}��&�ê#� �ꭙ%�2������~��8�(�@��ĴI��?�.-2X�D�Is��z�M���@���졞p����VW�$�V�2'��>�Oc��R@��eݧ�NtW駴)=�ʔ�ztK���Z����u��5�o_oں��p�L9Z������ih]m�.	�A_�׮v���s�6���w)Q�9�4I�PG�Ȉ��H��}l'-ەWmyZZh�L�������q����[F�7��� �ܨo��KН� �@��oyU��2�Q>52:!g�{�Ih0sI{��"|�+����\>2z&#�sh#�k#��"���|X$4�׮9#o��V4��$1N������h�?���;��w���;uݽ-�H��znn4�ܫ/v��̓��ZV	�?&�%��[�ԋ ����]'�u�Ǉ�����EZ�E?<޺��~� �#)���s�g8.-'֬�3w�9Ϻ��n��#��l����V����M�!aG$��0�t��X���4ɔFw)�M�v�)# J�B��o�
%r�|i�3�*9Ɛ.�*�T�=5�� �*:����:����!�o�����*�&9c1�7m�'%]oⰬ��\`���	�-����Xņ�W"^�Ù�S�.�)b�e�Ԣ�$�p�+�I��6�֌� [��e'�v.�;/�I���S �����DcTl
:�ی���k����;�s�v��]E�h+��V{z�N-b׵��>��V�����:��v��:�������a6#u�p���R�+�v��vm��"6�vkVλ/�"9s�ۋ�2#�[��rv��y����0����s���dhj�S���t�;t0�F��=�ܧ^�����+���[j�۲R���#�խ�c�WF��ˁ۪飒��eՕMs��vۡ��(�7����P:R�n�(�*�H��"��@��ڂr:�(�u���DfG�P$	(�1��7ʰ�`���'���"�S�X+U3��)���(�ں����}
�	�3�=-m��<�d�Fk�Җ�I �x���Se���)ц#q���ޮ���"({
U��R8���E�د\���x:j4��|�����Jꐶ[�#��D2"�!m�tU�����T�?�T/W�M���9�ao�ϒD��
�pP$E�Ɋ&�M C�ܯ	?�<-�������pT�nZIk��3�ι�G5�)P&	ib�Ows]Q ���6Q�n	��˓>�~�d�����DQ>��k�E������o@�qE��>�9�����8�.z�4��ڎJ���a\��eh���3bf[	�Kv���O� ��|���㝃�C�.���hG�Vy}��$�% N����u�δ�7���_{���u����^!{2��*'9e5~	&�`Q�G_`��m:��ƺ.���2���jq�iݞŦ����
�(ԩ�ܿ&x:�E[B��*��{[��:�f84! �?k����s�	�HT��`�OtP�ɵ�{S$��b~� ���b�	�!�pF���馾򥑦ܖ�!m�h#d�H�
��U����p�S��Æ�&ܬ����FE�M"���}W�}������wMv(v����^��M�5�����͚$�z|���YR��M�>���fU�ϯL�V���Â��L?k�ZpeC\��$L�M9�/$����̦9苦�|0o��O
�I�e�[I����8����L��5>��6؀F�`p�&J�$A9�ؒO�\Z���dj��9z?��]�U�U����6�$GN����u�׋X��&���-b���H�
0�qW�h!^�iٟaƇ1Y�4(�㰨�0B%=\�{���_@"$���}��N����7�x��H���L�ш� (�]��vHZ�ڻ�6� 8��"J#,��g�B��UD�V&|� ��m.��pt2{36oʁ���� �Z옒jw��؏���I"qQ�N�_�/<Ǣ5�I���	չHous$��|U���A��e�He����#�3Y�y��ԍ��.���Nf��Q�Tv2`��r�rK|�/�y�4�,�c�|c��y5�.7# ��2�u���փz�TF
�D�cd�LI�و:,NIStx��|٤�ܿ+�m��c	�����I��h�Zr,�8�=hR�� 8H[�nh�;��.���6Q�[܃\_	�{]��Va�i�	ݞr�L�6I�� N��EQ�l�OT�Z���S�td���'!-�������ؚ�c�u�D�(L��ٞ��V	���|b�f�����5�̎�;�Ys��d��H-%{a��z��T��U�֛h5z�8\n	W��Z�[�Q��{��9�]���v�����7��.�%��<� җu[�,�s���UY�gS��y�m6�r��ao
�4��=�g8�꿠3���B�j�"��MJ9}�vvfr�������y�c�D,3
�7�c:�׺
��x����M�oj��H&�.��tJ۫Y�vґ�3��7�{�jފ�^JM𘌯C�ܴ�mk�mvr ������ͼ[����p��J͞�q��np;�F��3�10z����H�#���c{p�;M�Wh��HF���{n��[�9�Sn���mҾǆ����k��M;�':���Y5=Ĵn���v�5�6��#6lC��^.]N��v�a�M���U7V῜����w�p]�`�����*)lT>�zEvr��6,4gaC��Z4
\���2m��In��:j��i�t��j�y.��`+=�ݼ,�ן�$%ann[.�U�uVJ۫ͼ����Џ3/��e�>��B�;��^��M�U�-qΗ��/�9�Z��{�k[�MVwbZdb{:��t��1S8n�@��RZV���w
5�/x�z��n����]#|���:��U�׻x��0f;;�~�g�*�c�)��G�nB�1O��q�u��MN��K���=-�c�yZ�Gv_��a�+�/(f�wv�	4c��/���9�#�o��
7�W\Ӹ#�:�=)������_�I��]ڪ���#�Ek���k�4ظ3#H8�xOcFW�i�6���e$@�,�(�7��3���f��Ŀ)��sf�rd�À.����S<�x9H�q��B��o\�Α�A �I�! ����t�1��b縞�w��2lOVAl��O��ۻaU��[��hDD�e!k�}��|t��	
��Jn{gm�G�\�y��6}Ⱦ��r������|'�D^νt��6�4�j�y�^���6�
F1�Y�3���N����N��V��֡���Gk�����cD1���������M-!gi�F�� e�]�۸�GAx������UG�<F9~�*ǌ�@`�Ř6���(�JGG8��H�sx�T��۪�[�2�]�X^ �pY���}D�r�g�A�?_H�I �Cٝr(ZC������W�A~�����ďǲ ���D����6���1�w:}�X��k��<<���^�_�9`ӄX�����H�+�I�ː$L��*�O��S@I('���Q -��zOM�faj�#�9��ZI�PYF�(��]B��d#&�$�(��?�n��`��$�n��L�!Oc �׏G�/�����ɹ4�F��Ԙ��>��SD�$�0OŔ��HeYD��{k����� ~�T�㟚h� ��Vws�����PQ6��9��4�}G1���Q�|�7��m\���ޱ&Ӳ!s9l�_��p��j��� ��K�d�g�����%����du���>9^(��\QV��^�քcm�D���@dϏ��{���`�~����3h2�Kn\�yذ�q�R�|~v�g���Q�q|�.�ŤA�}�{k��I���v�q�^g7T�N|"�7#r)�㵫�ݴ�`��-q\V ^��\j���?��m�����1��6�4Ͼ�Y@m�-��nD�� y<��c��6Vʃ�%m�yؤ@��YC/��D�6����o~����q��_��ZW�k��i�*q�܈7�d"G���9�nh�#t�Ϥ�L߁I~&	ڇ������>+���Ġ�DuNtH�	&c���D��F>����6�9�7:�s��{�� $�~꒧-ErJ�k��m=a��в1r���^�,��	�2(���uH1�����<0��D{_x��#>�7B�V�"I5C"w�d�V��5F�O�x6�@W�>~�r�X��v�c�.������$7�4��*��"�e�)��~ի ���i��	�<�T�%���
	 ����>��]�j6Uϧ�Л���@�Q^���W�z��t�-V�m��-��N����ǽ�_E�:d��I���ȝ�)t�O����_Ȫ_
Wl���*�2��!�r@�;����������k����G���M]2�\/���7J�4�qy�kdY��K�S��\����ǃ��;�ԯ�.yp�w�3y � �||O��U[U*�t��f���?w�w����I��,N1=�^���:�k;m�s�b�S&��{]�ɬ�mr����d��&'N8��3�x�&�3���܆�>Wsx�N�mǞ��l������ �^�n�ڼ4�G�ջt�œ:RF������y���uN�u�8S��uG7G7��#�xzݎ�]'G-�Y�N>����8�3�vy2�Sx|�˹lژ	$�^,>� ��qWv�#�f9��F\�h�*�|fڿ �袭�}=����l�m��"7��o�<��\�`PQ�j;��@>�C�F�����"��H�ֆs����L�e�=j>P�a$EG%�K[m�$����>��|��}��0��p����\I���B�F��x0Yz�� �9�&�$�9���ð4�zP9�\�+v�ѹ+փ7�˄�`�P��r�x!2PFJ���̯����+��P���O{�Xd2IfKpa�G���K3k�u�ǥ��#-�ޞ�5����!b�1ҹe�b��iy{=���K1���HW�đ�Ĵ/�	>�б�m\��ĩ�r���)��$P�"�����5�������_�{��=,���j?(J����۬kƚ���Xa�u:nМBqV�HyEwةO_��d�W����BLy;·��a͐��m�fΐ��d�UE�DV�>w{���i�$R�eM�R��!��[t��a� ۨ�6�|��D�k��\�݁4v5f1�������@4P]���X,�9�B֧�r���\(��s{�E�{X���w�l�>��KH�H!����=�=H	V�	������e��Wez؎�#��}~���j������w5����̫�s�]�����^��:sr�a��?����+Qo=��ٹ�į*]]���f+n�
�Ç}J�U�����^���N~!�l�@D�>��vX�$g����(��}ʅ1
g��h
W{����f#�j�r&�(��#�(Dȵ���ip֛�B�6�H�ޯ:���6�֮�Ug�H1�!�|�U��

�Fh��WtMJ�_A�"�WHWê?���q�F
s�@��L�� �{��9��f�~$�Mf���-�!��}~��h8�CF@�U��J1h���ᅅ�;�;�\��4I��#
 YS�Q�%���9[e���8-��4�hd�����	
�A$��{"��Yי0p�Ճs�2(M�g�x�NR$߽v�����:3b_{���6 _6�M1����z�9xp��?/�	~�A�3x6���v⩣�{2i�7;�]T/X���C1�Fb-���_��0a����6D#�����`A���>���3J���w���$���r;��3��8}�_ O�tS:�x��ـ'�Ƀ�k���$�	#����d![b4�낈Թ�?�i=���)z@'�t/"�D�Gu�)�A��<B*.�@�k�狑@�iK�<U�<Mt�G��`,���=l#eDc�x�-��c�%�����_:i�	��2d���U@�q H%���K�N e�\vD�rX����Nl�E� �����0�o��q�:a��v8s�
��u�������f���({Ҳ�صF�g;�}3��g�N�����~�����jC���B��J�DV�5D�)0��p�lfV�i�%��Sd��gH[0hƾ��r����vr^<j�3ս"��#
$R��$�sշ�N�4{�>s�֐��J>[F�`���Utt�Y��щ3 dMg��߭Ղ4B��`�\:�q,O:g7��Z�C]B�OSމ��r1l��{6)w��{�!�<�3&@Qc�o�J��ᄪ6��T��?�J)��%�[9�n�!E۰�}t�Z3е�M�3��9�0��'#���$�nP#��,�[�}�Z�M����D�
�o����!H��0 � תz&�޿!���1y�>�(�9"���c�ʨ ��AMｺ�i%�ДjH�|,�!�?m#r�*����͍���8��PJ`#��B�����Z%��+_d�?�����
A$�'ޮ��#�ofv����p��x�4�Mk��$j҅Ê��n���q�c-�ƛ�w�=�\�?�%d�=��h�Iۿ��v�3�$����zN7oS�5�I4�s�8���/�ۢ���\p!0�6��j~�)���]�L�l�H�=W���O)�z��$�!�C��'v�@<kiV�pP��Ϯ�Ѱ2�&�oZYq� h"��	���ǝ�s.�(2��e�Ŭ�/y��ǧF��ר������Z�>�VR��n8����d�zv�b�;���0�����>W�S����鞛GF��^!�Go���%�+p�+���6�P�����}���HADg�<�J����uw0VT��X*��I>H��t�)��Mzk�d��L���9�
� ��&�p�@RG��;�RYu^tz4SbH�F8R�kC��R#�n��K�	�xI=��3Uɣd���l�[x4�irM}X����Ý�:o�YB�@d�Fm���D����e
>#�{�D�"��������PQ	?v�m	$�]<���H8�sP�$�FZ�:�uYSAh���W�+bA�述_�MEL���.v�UQL�tb�O��w�hࡎ %~��s�qHb2�?^�ϩ�� �s�s��?/�"-��-�8�[�b\��S�[^�U@�L�q|������!�b}A-�q��~�:�"l|���&O��_)���4@^KtdT�{-8\i�2I`a-0ﺮ?v��C7��uo}����NR<� �P�!]�F<C �z����! a�|P���Jo݃|8��s���a �4�d^����]�-#uf�[�#o��O��r�gccj9��EX�g�z�yP�}�}�d���܄@��6����������Fk�@�o^>�ο�A{K��2��A�73e�ms�r�J�ʱ�ws*��e��4��+���V�X4^L���/�7�1bM��g���a��.�
�BٵW~��TO2�IT�Q��&P]͡F6/�tz��.�j�s�;+�ը-u�\�/Sy�r^�9�fƝ/kr%ڷhnMn@[�$M�v�Yɷ6�'��R[>c:�7K���^;���uO;zJ����rs����D�:�DDӵ1��%�5;c��vu��nj�u�N�LV��\�hb��ç�p�<x�f��m�݋�p\vӛ1vz�q�][g�\�X*w\�5nkPu�Eͱ(Omy��NH��$���o����40m���׫$��Z�R��ާr�?z�Y=����:�^�M}�\_q�ݏs�������@��P�0K�eQ���npnT�E�IK,�����$���z\�U��	�,����I����d-���� ����Ȯ�6����jb�D��Ƣ��su���o'0��ggE.�"o-���H�b �DI�Qj!E��ހY��Ո
rw]Q��B����Z�_�$B�nZ�.���w��N����o�Q-��:�X׌z#u6�ݴ�',YY������+��)ã�$��t4�`� �OŔ�^��3�� ���&�$��5�B�^�	":s�r��i�߹VPmMo	�~���V9-f9bI���*����3��wگ�D�#
���:8���'U��u<�q�;�{KF����_Bd�5�N��60�5*	(|:Q��g�?��ӂ�B��Ui��m̅��jC���q�i�h��m��ä8s�u�AЖ��|������J�i�޵锪��p/LҨC��(�N�H"F �z���\�T�L\a�W�,F|��$�u;=ܦ���a�"Lim��k���K
Բ�u�/��������^�d����uB�e�y�t�}a�D���ӎ%)]�έ���[�"Nsj8�����M�To1�`� ѣ����mL�-�������et?x��${:��s��4E\A�.���_i�'pP@���LMG�Q�3�9�r�b8'���j�嶜n҄$ћn4y!�J�����DQ�F�wD�ǐb�6l�We����'g;Q��v�����
g�ޖ�]"(�q�f�>=�+]p.#(��h�Ǒ�M��w�&��������-dz]��� �)J��]cw]�%��̖��5����zc�%q$|+,�z���d���c-��+�7ֱ�`�.w}r���ASb"���5ܨ�K��{24�� ���F+z�՚���r��:=��\F�D59�$���Rs�<yB���Zծ��+-4�5�H�AF;WY�󵶯"At�#���7kr�g6c���u��M�^ϷVE��ʒN[�M���sf��n��)z]��B@�85	>����� a	0O�@�kg-���H�h����l�u��c-�[ ��IlGu�L��\��ܕd���,��现kH� �;�>5�� �����_�O�z$m/��Ў��'gi��x�ƫ#����� �X~������#+�:�#��-����NP&���WDa�C�4gw�ь���N��A�1���u��(��aęGq���MS���7��x�{5�Ү� �7!;��.qS���ࠥ-���mo�z�@���s�q�2��=�I"�_�I��deG�}-El��m���v�Z��ږL���]���F�7}��eh�e��4¼{v�w�RF���V�9's��TN�E�p�	�R5ox�*��^��F_��|�বQ��ei��x�U��,���L�ID#OR�&�W�,5�3�hF�QɎ|3�>��l��d�@3�gz�U��0��Dl��H�8���>#aH��x�h�Y\�ї�e�V3�U��0�5��ŉr[;d8e�
��K�3��z���1�.�����NTJ@���r٩�'�]��h�w]�b��qJH�_[������*8_�qy��),��P����Y����� �ߐHŴ�X1�&�4��@�$ �+r���>;���dA�߸M<G��T���,іص)(#�s5eG:� �����A���W�"�Ϟ�"�����0�TQ3ؼM���u7)�۬pK`��{*m�2U��#��2(���<�4�p��;rU�Ă3}�g��ކEHB��}�q�6�֠��nt�g�=a\v�`�n�^t��pkz�湇ߜ^�mn\�@�]�ɢ)kD�<An����cg���~��پ �W� ���~�����9@�#���N<��(�c�u�!����#Y�
<�r�:��\�\�sw��k��?j��WixH!�`����^\��Ʀ��΀�A��k:�����e��%c)C��:�����E�O<��O�P�fԛ4;��8D��P�����Y�b��)�$�U�`�"D�BH��[�� �,�X�����h����a��*A�vi:�z�����EX��9�&U�NK�,�%v���S��������1g-�}�k�� ��E0q_{��
�0J$�ۦ�${������9$+��]�gbD�D���`_�~�Mn�Fb�$}Iw�|�dA!�R;q#90	�Y3�T,������
���Uc_d�f���欄
D���Zr@�3}!O��ngb��έg��
hRF�!T���䀆�mN�-�� �8p�ȹ/��6�I*F�B?�R��"��O�Y��*��ܙ�[��T$�H�0�T��yN%`�NͶ0�*(����"���BQ� RH�_{���{��n�~���lH�AEZ�$���}�E��ԅ8k���dQ��D�s�cҫ�A�#=w��Δ}�N�_eH�9�m�ƥ�e��.��nx��"�$f������⫟�$|�)�C"�d����oZ���Q
�E�����7���hSqc���d��f蚆<ٴ+�}������N�X�:�N�����SU����k[� 1lĉ�:P{���)~8kՅZ��K�1�I����2p�(s��m�{`��G�x�}�%�8��2��&Ɩ�UH&7Qr�'-�w���y^�nɾ�s+f�<oz򣾏m�2�$�[ e��+��٬*�p�ɛ�Q3{�ѽЊ!��bJ͖�h'6j��֍�\-��Mn+KE@�]�s��|j:�.��KћZ�J1�\{�����`�@%gL��66e���[�:�^��QL'�M��r��Z{9�CE`wϻk�7/h�Q�]��2�T�.��>)>v%�7��,����'T���X�����S9��.v��F���gVRiV�黷;q�{w��"'/�M�G�n��j�4ۄ��I��F�3E̚X�z�9��jL%��pW{�����:I��x���7��=�\_9�&��vn΋ Y�,���'ACG`������B7/Z�������0��;a��3o*)Ov�n�ew�f�p�O[hʝ�K�ؤ�J�;��,W����s��w�󫧲�'���΢���2��K'o#����h+x�+�楠ԉ��j9ҤLfԸPR�{˝aߪY�{�����>�[��#Y����/l��ɚ���B��K(����V�t0���[�h�������4�YV1�spE�a��o6�жm>���ΛO��2�W����\��I#mĢ,�$�	$2G�{;;{;w33۸=�ї$�H�%�-�mUV���*�UUU�V�y���]�&U�v����eZ�UvZ��Y�dR�[SF�uY��I���%l�2�y�G�9�Rh5m~?�+wt�X�Q�������/�mR��lႍZ,5�)^S��(�f�����ɱ�M�8�>1�Ǵ�����ո�_2�1s˽��䲪緐N6]��U�ǵMş�>�}vϜΒ��ќb�g��ۮk�s���m��9�nyۮ�2S� �к��w����Y�{=���UB�k���de8����#Y�.x69봳�����E�Yz�k�5������&�����5��5n�3�:㎸<�=�gG:�����3j|�/\�ζ�N]=vΫ�����4q�_$uY�9�֘�hb�b��m������Gn�J	d�	{;�Y%nwm�#ɥ���X�=�Z+�[s]���m�ۓ��t�㜻�;��om��q�s݊�ng��:�op�EO
�Yq�[.�[�t�����;����l8"pn��#X��>غ��G�7X�<A8�mێ#�[�>}����u��)Vv�mN��ݯ*[�^�y��&�q���8g��c����`��pqn����0t�X�����Xݗ��-�����v���;9-8�ePgWm�����t[=�v�A�˜���3�öƼ]�=�/n{e�ݶ[���&8�m��p�s�E���e���=��a�qƳ�7G(u�.�p�޽��vr\-p�M�����]%�:�w��UK��\�`�1�=s�'k;�gN���ƕ۷c�P�8�����ö��r�؛s�\v�SN����n��݇x�{>o1v������3q���n;c�]��v㥵�ú�:M=��h4��sq�un{��{U��bLX�d�k�7����;��sˏ���/g������Y�Ǭv��.)��`�H�h��ŷ'=��4�v3���'`�Q�-�N���=8z!H�v��\�C�	ö�O:83^z�Qū����l҇��=;S���%�	���?>��>�-�f����&�/cun�\���k�Ů	G��<*CkY9�W8�砆 ���//n�f{T�6۷.��l/Ǌ#����z�&⽎B��Z�<;�ض�tV6�^p��\ק��]V��u��.�7�����<�͞7m��Y��y!ؔ�Ɯ��q݆����q�p����nM��5�$�q��nʗ�tKvF���W���/�#k����1�}��lGN��My)����g��^m�曣��Ib���_� �r�C1�{{�Z�F���(A��/��~��p�0A�d�FZ���>��~�Ñ:����i/3�b0��(䊴�z�^X���J��Y��N��Y~��ʏ
@��:�zm��	^�S���]u�p5]�R�!z��#pi4JbM��"r%��qdW���N{���#v6�r�=�D�b��������X#�O��6�OyE��7�;�/�M�������˫a�G!���|���?Q�^�cx��ϫ3w�\�����G��wzw�#��qjȹP��Te�$J	#�ٞ*_F�&��!��W��G\���o]��˷�2%b�s�|�}�\ws�a����XZ���L���jhv��X�Oc:�㮙68ژ�$c�qnD��v�k�F�ٰ�K:uΪ��N�jL�#w�p���]�]����qK��2yN�H�r<(ߔ�Ὢ͒7J��N�?�H]��|Z6�M*S�pz.��M��&��꼀M<��K��;#%t0d"���٩�b��|��'2M�Y�6 N��U4�b��ED�L�Ԍ�y�8���[��A��ř��&K�����T�!�?Vu�o����EY��*"�XI`�m����aSK�{�9���{��_x�v�����u�Vr�����m��Ul\�s��s_־��t�18����2G�!}�;l}�����f��+_����S�Sޯ��(�Z��uި�>��zH����>��[Tz!�a�	��m�ٻ큜8o�ܕ�F����p�Y�k�@�;�j���u�sQ�-}���ܸ�W��Muu3/�&8��=���Լ�R��xM��N����`U뫜���n�CE���8�h�b���6^�3���A��4ӈ��q9���9E��'��4�H�[T~н��wP~��Z��l�"�qD�,I#��C���#��tO���S�3�}�D��@�ʧ��h���=��!��OOUE���z�L��Yց�9�p!��p�C-7�32����+�q�C�)DW_S�۱"�Ngc�9E� ��C�U�ʛ�^sN�����;���'��L<��oCu'u֑X+K�6�f�c�U3�-�W0=���{��?T�_>�ވ��F�E<{�Bv`H�܄�$��^]n��b=<�|����;��.M���W�L�?e�~���>���O����}��<ByA�9��R��2�B����8���G�׽B�{_Dv��Oz"�<'F��܋���^5�_Nen���Q��ז��<�ڨlP��d�lv�d�S��n˦�z�]r�h�)������t�<@f�\�1�f���1���]������=�v���w:Wǵ�5�O�>�~���_�<|پkG�ݽ�>9�ࡂC	P�!M����ܺ��~��Ta�U&߫
o�J�z�ݗ�ߦ'{�Ϣv����w��]�\�|�.d..�G^��%*�re��tn���������P���TB~��N��^�«� j۝T0k���p�{����,���uJ䗺�W��Eɐ���#��q��`�L�5v�P�C�8C,��I�pᡋ(sQy�H��m������-�O�w�DEt�-�jm�{.\Y��7S�J)���%d��h�e�\�]:�;3$b�+D�'�5��^�n���+�}�Bd�j)�M��$ɻs�I�tNe��#��d7������rdf!G�=�����Ğ�f��=���R4�Gz��U�P��� ��6��x�AE]�9{�ɀ8���v�c�۳�$����	���D��H��9���>��� z�^ݷ���H�Q3;�?|��*�<s�!24�u=�w=�u	�W���D@˒^H0V��V�a�Ѿ�&�E`:��]����D��y�,�<p��u���sr8�,0A�ٶ� ��_�|�Eт�9/�D7��ף;yгO-����]�g��k^��/θ��Ժ��ϻWNZ�����̋#	J8JpF�qޔֱ/�_���ߵ�����k�W_y�*-"K��9���ũ�GT�m<���ϥJ;l=<f�r2�IC!p�c�C��v���L�'Y���Bx��V���#�[��ڔ�3�q.����]�Xk#�
���z6�܄��n����X2��!�^��2��f�U�L�zU����(�<^��#)_����/Hn�ˡ����fZ�ک��&��A�rI$�I$,��5Ք��6��/O�>ݧ8NH�(�C�T�`���$�Og·����z�8���A�ٜ�u�;s4B�nb��d#s��<ۚ�lt��ݞ:�A��h�Hn#<=8��Ź�e<��j5�y�������hm���L燵ƻ���rص�d���4�#�=�7�.]t%���s�Rl:��S�������;/��M�[]��ʹ-cƹ� 3�g����g�k��y��;�'�I��A��s���gm�Gb#�u�z.UyپȱH;�����=���Wa<qH�η� ?fT>��qM�Q�QI���믱U���|yz��N�����G����^GOd�W�\ O�gc�ۿ�!ycbB����q�d����x��
%���$��ڼ͟����;[S��r�\/��o��������y���5����U��=ZxgR(�0��
��z�;�Z�h�tV\���YbN���P���U\���M|����Z�G�#��Чla�J(!j�q6Æ�@S�%$�`��������-��m�����rs���[���<�9}��a�_k�V��M�W(���N@�v��v�_�A�AA����x{�GOn��ty��d�q��H�- �8ݱKh�
��m�{��D�}�@��7R{����*
/���i�xl�tw��ݭ,x��sX�5?&��&9"��C����cH�%����m-�Fd2a𝽖G֘#씳��&�L?�O]Âo��P�B��ԖԘ�|W���
W�V1ܱ2�,��98�^�̼��f��x����7��Vb�T��}e�T����S1����KM� ���ZI%�]!�.�Z�M�;z��s4�r�*6�=���V�_Q���y����S��H9=��&}�ŕ��]��0i��fE�6o�3�<�4=��:�~��]�cRP>kϷ�Ő=�x��� Jy߹k����Ew�Q4�eD��Ĥ�`iu�>���k�^�w�,��D���o{�JU���dt���9�>�h�a�SY���,�������8��C��wfk�d9-Y�q�	BW"1��W1�Z7-R���}~����~}�;�ti��=�߭���7��nz�{�#:A��{�1#\;��#�<�zH��i��AR?{�py.O��k�Y�z�����=>��'�^=��g�^��l+Oz$\�{�GW�,�4\��RN:��/�qo�K~@�2��fW����3�}u�[�Iح��g��댫��N|<� u��cf��H|3U�8��9��㥙��:D��}���n��fr\l<�k^eF%)�Lg+�ɤ^K\�>�����K3.V���@�U������?A�}��d�KF
����1���{lLǤ��T���p���b{7�9� ��;��}@��Bw\�wPp}��̾�!�{r�ϑ�1'�B�R/�9_\��qĢ��˝;.$����eǨ�Q��gS�h0o�nF�OG-�����"�C�w:�&�~q��D�W�]�EAkjv�ER�p/S���-�La5��=�wi�9�zա�mv�Ƌ��u��:R�^�9�9��fW�ۮN<bY�i��Ց��d�G�s�C`�DQ�0#!jG�F}����������<y���&�ˏ���;r����[2������M���Q�����)��^����l�
�w��3H�Uy�>Ÿ#�%�`��^�a���z�	Vs�{�Ǯ���Uϥ��WyfWl�,͕��E�ڈ$�՞������T/_ۏ�G��8�޷"��g�������Y�����b�ށ �gl��w&�̷1Û������7j�͓�m��f�� K�'L�ڔ�ʱ��en��B��ë3W?}b�xٔxo�e'Zm�z��������|���ꚭ/C�Sށ]��{c�w�fD���{�g//3���Ȇ�*x[L��@�;Q�]N�q� Mk`�b�xxz�X�L�e�-]�%h��{�S���A�;��r����y���8����g��>w\�Ʊ�HU�d���3��O%}����(Bx��V}7���+?y�	'�����g9�ۇq�+z���wT��`�����dg��{�X�����	&�$�!1ȯ�[R~r���3�D(�3�ߧ�>�^�>���p���N_�"k.wcG�Uv;ۨ���\\J�ܴ�J���};�״�;����a��~���޿��MN�R��#��q˹���{��}��WHr�,�9	�C�yN���vʗG��a��w+UK}��MO}�3=]�C��������U�v%UN�/��|�q�D_5������)�h��زd��1֫�'C��u�Zu¦�_1t]&�2�=ܘ���mi]I]�k#OL��f�dn9$	�m��n�ؑ{kkf����>~{d��؋sm��۬�:v&I��_�����%�Gl�ϞL���^�:�yF�B� ��us��{\t۶8�J���p �rT������SU�̊<֢���rq�ۛ{��bvVC\
2�H�Ͷ���[%Ԝku�v�Τ��s�g�ѫ����p�#m됓#�억ab��d��{1��V��!*���{voY�b۩5�b�N.:vr��4�����mc�)����+{.�TGzb|�>����"����+rW���9��3*�<�pT��?u�+I
��^���t��>m��*N�����~;D<��_J�}����ٕ]O���);��DD�C�y� U�<Co��m��Jd���K��Ҟ��!�n�e+���T���p癱ʛލQQ�^�wn�f_Fk��,]�DB�p�"��s�.��w��jD�]��x��O��sxqW��~�l���9?;�+"�s��髙�;�8Bj@�-%ERo��R�}+���o�!���*ˏ��J��5co::sݜ�y�}���g4dY�r֬Hq@:�Ů�]��1�{sΤݶ.�wQ���	��Z�����ZIl��;�o���}��Oke�5N:�c�n��M@��[�'^�EV�&�J����3��.���#��TE��3ǰ��o7����Z��>���ދ�$��T[+c���\'c�%`~�/v���ѡʞp�"��*�c�!��/TYOj)ί9;���vf����Qy^ڋ جq����Cw����}9��_�ّ27�pWƳË�V��f��[�ό�j$���/�.N��D�"N����eN�m��.܏b{]L��`UX=3��l�M(0T=�0�F�9QSٯ3l�4��*�tw)=[8m�O���˖��xbB�K�=��V��%D7������
	�$wgD������j�~�S���Ud(v�� t�uO���4�	
f�tՔ�ț�j���#:�a�v8�~SۙZye����E�u(-��/9�k��ű�t�r΅bR��j.t�qo}�}?a�R��34��3�rW�e�YS2�bs־����rI���j�d�aqQ��"�$�L8m�T-���>�?{�7f8�]�=�bj��J�}7���r/tz�����;��z����7~�}��7��)�F�5$�~�`�_D�)������ex�y�eQ�d�5Ҫ�O4lQg�ޢ���N���Kפ�j��J!��(R�n[m�n��`M��d��V]sW���o{:��V˻���5N���t�c4���a������{x%OXUz%K�V:ո�Y�B��o��J�"��T��+��eο�e�n^n��K+�e�Xz9�_����F��w,>��r����h� ѩ�s}Fձ���yĺ4�'�sgZ��O-�0�˻�!�v<��mn���%��2�V�q�u����6NJ4^�����v�%q��+FK:�2L�/4 E�X�֣J�6�{q��]K��Nk�%��2Pt5P��ʼ�neǣ�{�|�}Q�����ގ�Kn���g���ʳ�9G�q�{�ef�{���_r3*Z;@������Jp��^�v�ǕՉmZ�0.��ˆ�ը�;U��E��Y�N��{����м��wb<�z�Z�݂��4>?4���n��f[��G�2xɛ���I�b�(�^�1&nīn�dK{�+��l���fH.�XL�x��x�a#�Z�$����M$h7n���ڽU#r0oO�w[�m=t�R�����!Ѫ����å������~7R�"+K��5�ꕑ�|�*"�n%}�f���f͹�@�㑝��e���jY.lbٶ�5�L8:�u�ur���؅����&G���pW�3N~�;td�"����]a�L�#n�^�<��q�D'j���x������܎��y��2v�5�7U�Le\���e���rIo�}#�5��v�Y5KZu0;��~��(�^J�]��~����Kz}q�#v�dOU��l�S��7:��v2�{2����;\GxC���><~�'e_G[��g�dzw��lH�)u�����v�N4��Ȕ.4ԅ&���|�#�������f~�j���Es��2h���wQ@]�W5��=c��yI��x ϭ�*�YE2g&s�Q*�ũ:�	��O�̑okj��7e�uօ�D3���=g�������=��T�q��뵙��5���R�:}|��V"�im��g���A&����a��$�5�g~��s�Y�B�;q[��E�f޽�1�z�;��|��׬M7;:��q�gyx���Y�}�B�H($-�R��#��|��>�m�/�(Er�t��=w�d��:�랜�F���n�zXYN��,�_�M7�A$�.{�,�~��]��y��ݝyK��w�Z�̯N/Fژ�N���=��1����n�Y���Gl-�>���!鯬:�2|*v4��Ő��JW-��ۯv�z_��dV���Q�׈fή)���&�9U���0�
���CA!�i����+�����+��ͷ��ˢc�q@��[���(K��GW>���9L=��#��H���Q���̎����������qo<h������1�&��(�#�0��L�ĸ(2Z,K�oP�N�i5��*c꺉�팎R;V������v�.�
�P�wL�(�WY>��������P����0947c�\��R}�:�?H�%�D�Y�^\��:3sE��w\��Yn��}^��(xA�4����s;3��نa����:��Y��~x�Ś����vH��muIt�l�=�:���v>��C>�Œ�aU-$�m���~�'s��7̾�X�I�i��!T͗w�6#��G{�t��=ڬ��uu%h�>��?���p��l$�u�C}�5�J����>{����zGA�#�ͷ��ϯ��R6��o��7�^S��oa�����6�8;bx��{�K��2�YQ�R�%V��	upQ[�w�����Uv�Ꮋ����{_��o�3��{����˖�B���X�#,�IT��]��r�8֠��(���y�Ddrͩ�흴����ܺ�^�����9�x0��n0�]9���G�Cv�Q��'-�ۛN���7�'����=$\m��p��ݗ��y����OPL�]���i-�'3��s�.��8��u��v�oL��=�V������ϭ���c`ujܬ��J [�N�4�\�����O�z3[
	ܐ�����7h8�q����^��L�a6\7�Mί�/��hi�[�ۛ�`d��L������K�7��9�Q��O)]�����+��P�N-4�f�h��ޟ!~����q ��I����/�ǔ���%��sdKK�����屨�G��w#�8�V��L�8J*Pm��_��c�ِ3�ʺ��B2��ƆEDŭ��s�v��Щ�����1�=����E?F�N&�?�_��Ǟ�u0�f���yϺcqd��(��NWD��x>�	����s�z��H磝WAV�bJ�V�E�d�,�ۉ�\�R&���|��m�)�/V/�U�J�٘����~�`X~�=ז�׷s�>�H�,X��أ{<lv�E�=l]�,�i��;{m��B�M=��O\��EWn�U�4*��c��߯��쫧���b��&���,X�$�����:�=�9^>��z#/c۱����\g!t�P�,9�E�>�+�}soV��{}�*
6� �����=���@ڛ���Ъ��4g�U��l(�9��^
^�,�n}fVBʺ���f5��l��Ԟ#"<��](TPם�_��7ߠ]	�� ��S�v�4�\]>���������vR,�a0�����u�ʏ�߾�7����)��\9�egg��:��K��No�Y��F梘M��,0�Îj�r0sAnؾ�Z��q�����yv���῔[&;t�*�
�sU���w�Օu�;�8fm2�2�^�)B������!G�-�0��k~ͮ+�}����1v�O��Tf����k�7�`u�̧�-^ۦ�)��7m ukE���-m�sJ�nΑ�\e�^n�=�@ҫ	pBH�v��&���z�����M�����w&n���.��k��`�O+~�߸٢ZӰ�����3jDfp�-%�7��+���ޣ���KН�����G��Vת�����\�w^?`���b�B���u�L��ACp� �CU��tW~�aHb��#"���뤺ݛU~����9;�B���Y��=�롼(��oYlb���3ln�lgV�Rv�Z�&,������Gc�1j��"3?~0�>�f�6�߇q���^��o���bG
q����� �#�A�w �ٸ�#fgޢl�ᐊ��u|�C=�<��Y��y	���ݿ}�@�_��Tq L�[.G�ۄ5��������T�O3�9-�[�_Ϣ�|bR�VP����z���1�� ����6�=��cΙnP�U���b��uW�qú�Z�>
m!rmM]Mˍ-�ɽ��_[���׹+i�{پ�Y��&"{�F���^��s;�}�v�쇩�m�S�0���!�1$���}�/���״c����ˎ�~R-mӧM��-}�]yK���yXRvn�G{��B����jg���������!cg��3�B��/�	_L۷���T����z&���d����P9�7m��{����jE�����<cFϧ��ϔ��=ռ�=~?{«"<Ҏ�5��!�p�ڲ/*謔;{�zP\��X�7�՗{΍m"��f��|��˖�V-5�w*�vC�5q�W��HKjSy�k�	����k����5����!��L�}e��\!��T�;���UÛ�w�U�3Q��ڥ�r�����訙�zo�&�Dw���9��.lI+ˡ@(ח���m��c�(�¾@��]B�9�ѻ&j�]�q]H�DUi[�,�������k�9�/���d�q�3Q7B��9�N㲃�����#5,�<�6}J�]�m5�Wjx�]�DL��۰�ށ,��{}[�����u���{]�����6��X��)*&բ���m�,����]=n�*C���"�v�O_-�b��p���֬�F��i������s�u)	x��n�M'��ǥ�p'r�3�xiA��zX�s�]ݖ}�3`s�����~���������-�%����$F rI+"���Z��U�7�~�qB�l�t��ȁ�T�S�G�ψ��^��J�U1�QV��6�P
�AnJ���E~�v�e`�2���N���zx7����7��p����fr�lǶ'����4�x�v����m��UUVq4lulr��N��S~57]��̛&�V��ۥ&q���tm���M5�n*g�7^��;'���l��;��)�]�$��D�\K�)t��V�X,�s<���.ܺp�Jwg�Ӟ��5�
�+����1��b��yz�>�ļH��t���Yظ�ں^bu�u=�p�mҚ�G�c�q�"͎��oki��:1n�q���i�;'�z�~^!qA�������1v������:�f�^;P���z�o��oA�au�+���=达��G���*�S�b��3���^����!�q� �@�Lۻ����n������=��'4�w⟲{�{��	;��.�
�1�r�4�J�Sؙ0M#�.a��N=��7��pߢ-���u�do��~���ظ�׉n�ۖE�x���^�wS���a}�H�n#��ѵ�Ƃ�������9�^ډ����W�su���������܏U3|=�^M�tߪS�WPh��p�^�xu:��~����~�ъ�ɛ�vit�oL{�7��<}�+ۚUI��c).��;�7K�j͌w*�D;U0\+���7G��sc��u�(�Z�]Y���h$�NVY���S����Ƞ�U�۷������[s�6�=��
���?O������Ng�����N2�a�-���}�j�6����WƅЌ��(&uC}��9�b��WIo
�a��Z<��82�V��Ȼ>�Ƕ��b =��U��A��r���[���E%�^�ͦ+��D�?H�Vs,f�zo���K���8!8as��לC�H$�$������g��G|��>}Tx?\��+���9Ծ�9ޠ��֡�k�%[��iyl�}Z>R!pG�=�N�����k��ǫ�n���/b��@$�pq�|�/�{*D%�y��˃l{c�WI��f8�	܆�-��}�>�|t�I4w羑U�ޭ��W��豇3# �t�K��5�u���1�c;T)�M�8��ܸ��]�u�7[;n��s�+��zX�묠���aL�Ƥ�����&W��w��}��ޑ�v����Q�Z`���_v�o�=~�Y9Z�	���AFam��~jr�r�[z$�O4�ם^������uΜz4ߩ|��ԋ�M�O�UD�#�s1�/�0�.N"h�me�r�p�ճj��|�z�rê�u�؂ �4+�^�uN�p���g�Zo�l��CH�@	��&��b쌯x᷈9Y�4_���K�;���঳�.o�w2���ŕ�ߠ��-8+.WZ�a|�
�䉧!�(	r���u�lS�#Ʀ��K�26-��}�F���y�6gkyG!9~����4W�2wzn��!׬}|#P8"�(�J9��j�_gՏ|�׽�H[���R�7�Qw�;��<.�c<�k0���u4�`H�Sҥ,��B"]������Pph��:9��u:�'�[�����Z�{)\���컡���\����H}˼�ٝ��O\X��w����hB�I�u7=ORy1���X=p8�hs��p'�G�_������~��Q�Pg�Fi�0j+#ױ�\��?L��w��up�o-�����-r���5b��+�7
b!�fG�¹��s���{�كP�_z�ySl�G_^h!�t��=�M-�O���}X�̽������~l�Xe4`��K��=�|h3��n뿗`��Qޝ�9yy���:/�sє3;r��Ƽ��f���ϒ���t�qKeo`��:!\t�6�T].U�e�U��B��8�t3��WQk.�q���b�>~��g}ݵ�\�̷D���F[p(M����U���Rr�<��ܔ[d{���9G���þ����=�T��W�m�f����y�BD8���?���O'p�v�����16����6�ļ��ͱ:A�\�8�
��~h���и�LT+�����ɼ*��)��{�AAm���y^\a��������U>ߔ�T����B[+7�_�v�w7�c�ϟ�%���_}6�US�^�o(��z���F"l��5��u��w�ku�-Q��-&[����?���h�\y��k�����g�m^�����𺛽�~hH�>�݂���V9]���@�P��I0A�zc��s����j���ʌ����X�Ǆ�����{CV��
�zNCSٝUЮ���<'x�\�d� b7V4�w`�ud!����
U�o+`�$)�Z��:n#N>��#զ��G-ˑ�X:qb���s��I�;�#u����uhJ&t&�G~�/En�(ઙ��5D�ݒ�].��Sx��㻨��V9e���D��=ݮ\����;��ι�t�z鉛}8?��cWX��R��K��k��B@훬����}h��o7�/�T��>Û�`�Z욏EݻG�]yK'Z���]��s�X��w�����,�&�4�\�OV��N1����Pټ�-6�#��Ǻ�V�y�m+�Ti�8�_�mvF,JT���<+��v�F�V½���B��`5�=�ʩ$���5�g��nXm�Bs��Ug{�<��
u�;3q^WWqL�KΙ���3�%KQ+��-������S�0'����$^)�^�<���������,7C��#�ę������J��t�$u�ѕ�����+�tpѮ7�L �����}��k%�H�.��WS6n���-�ufd��#��:yݰ�,�����6�\�Wj�q��jfD2廛-Rr�=s�eh�m���xZ梆�W|_H���I�D�C�n�xu$N!��,9��c�\T�M�F�j�\X	j;�x]��u��Q��s��M�
�.���a�Ytz[���*���z�|��h�I�'}����V=}�5�Y|j�Pq��qh2ح<@cf��ф4�k��7r=B���Ww��ږov�C�Q���j�G�Nmק�z?�7"J%#.#%nh���������$�$��$���|�~�f�2ꕂeUT`*�Z��+TR�UUAD֤&U��j�F�
�����U�9Z*�A	�Wmbs�c;i6#���V��Z�deE� �x���k�*T��R����,�	�;��?@�dq��qxPK����[�y.X���Y��U�*K+#!�<���mظ�6���]�����C��r��x��:�sc����]kX�.�C�j��ɮ����:"1c�^��r����]mkֻR������Ii��2��:A1� �*b`�m�SF�����S��ky�:��ps�����e�6�\=F�0[�����?�v�n~��e�xRx�a������8\V��v�<:�τ�*E����s��r�=gq���E��6٥z���.mt�L��t�k���T��c���r�f���]����^��\�C� H,��㋂�-g�u�v�XҼ����Gm
�OO��.[�s�͡�Vr��答{J�c��N8#E,v]�f7.986��sBݣ�<�`k��.בY�.�۰�:��h��K��-��v�ڻy��d��v�t��ng���\p]���t��"��ɷ}W��zy;s�*��w��pn{�kU�JmF�m�ӱ�M�\���;�u�3�e.�[*6�<�v�p흻`��{;����۶��tN8As�u=nxn�v#��60��s�`�S�u�M;����v�����烵	��E���by�=2;
��ͱ������s��&��S�α-���	�s��-�y���t�-�[�3�;m��㚛�0�A�qꊅ3ЂA����۲X����l�4s�ۣ���0��&j�78��c��ƺ��.�88�X�8e�m�D�f�r���q�a�q��Ӭ+�B�=U�y�7lOh痦�=��j��ƻA[�8�6�pD�ò�����<�G�vˮ]�%�i∧��;\�j�@|��c����\T��-뵄�]���֘ù��t���s�˫=0���<�%�ٸ�0Ln��^��qnHv{`z�:-N������󪹂��e@�[k��mە���s���_�&�0䁢闲99�jqk��r"���tʼlʝ� �՝������X��5[bnh���h��<�uc7O���d�o`+���Ð���ù�շnq�ЛpwkqoK����H�9hUS Y�W������=yK����˛�n��7A����m��lR�WT[klu�!�[	o;\���w��>�z�k�[Zӧ�t;\m��;�Kz�d�A��9f�2���:��Ĵ�x��X��d�Ws���:���UҞ��)U�o��qE:�]Kڱ$s�=����M!Z�=��*��w�`ܙ��Va0'�w�wsLg�ڼxV)���zKȏ�s�{F#�0�Bo1���uw��P8ڀ��&���&3kyu����]j�g���e��~��s�*�Sɝg|	��Z�I5f9�R܊4�����|��Z������|{���*o�o�;��/����H'�^���O�R��>�/Rk\r5�NEYXXF
���,U�is,a�#�ìt�_<�3c�H����y��w�e�ׯZC�aͣ����Б�4B��l�n��6�gf�n_m�헛�PX�6ܭM��3Φ�B�9���������Q�=޷��Xh�q]=�1F#�:/�6*�u!	u��0Mo��s�>5Q':84ᑓ
��,;̻�]��0X����kE��p[��؄�l,�
��9×nTV2vY5AwW�}!�W�i(���'tKh�u�k�g,x�h�s<��˅��L�,~b�OOe�~3=�LM�=;1r��vxd�W2ӆa�7l-�������ug����������nc.�߳Oޗ��ߢ���f���__�&/�6�I�ĄƤ9i�'�x��q���;�?��!ฺ>��ڝ��'���"�k�vQۃe�2vy��P!&)�ա�w�%{�ϧG��{�\;��F-�z��y5�������]�<����tee���X�q r�0Ε��9k��j���㵭������y�b�eכ���QG�Z����� �����2�����ɗ����ݓ 렋���w��߅�DIP��N-իC�}�������OmY��O�χu��_�
k�M����_������7����ĸ.�&��[�E�r�k��d�����ǟLD>  ?=��r$	�u0c���n���sFK�\�w):���E9q����;gw)��ۥ��t�F-��U	u��S�i��ly`��O��h/}�_�x�mz����l((�)9ۗ(c�����qc񸹸��~5�>��ő�{��O�֢�g�
���w����]sA��f0XrE��샭�/���g�4�豝����^�
wz}�̕I�8����.��1�"I�ǖ�՟!��.�ڌ�I�^M�cn�\+�P;an�C�;��qv1L3�����>,��4s�\��~��n�Կl���^�����}#F�����,��_g��I
��)��	�^�Ⱦ�#z�*�s��{���z&���t��+:g�p�{A�Ι���P��nV��D?e�@JDe���%��{�}�uY~�3}�Y��5�矩D`WާAE���;{r�����^3������Y0	pYN!���Q��/�64]Y���s�Ļ\��"����/^��!h�����_͐:}��q�m�>2�^c�mN��4us{"(�_,R�4�e\[���f�㋵�ٺu&���5�쇯k�Y���z�em^�s_8�*B�qD�qV�:D���L�������^)&�SiL���wy�x�1{�N|\?LgGr���y���|�c���]�
U|�sWCL�N�n�0����fn�Hk���|���p���9p2���_�����\x�鐢sR�&,����ǌl-�_N�5�^fr}g�"}�+��L&!3�j"���m��v�#s��<�)�sƮ��򓑯x.�F�e��ٳ�t��������*=�S�hW���������0�6�{,L�Ur^~�����O�7�w�u�g�����n��7{���Ǫo"��M5�a�e6sw:��!�aT+ޥyҽG�Z�;��Ӈf/UjOr������Νh,��������N��u?lal��c��_��Z�~��Ob���^��4���uO����_og�9?vd�[�")#i��x��5�k`b87���8bf�}��"mx�!�/i*l�eK��ƣ��,([������y:�$�.e�VK��J�һ��j�U��6U���sK*���r�5b�;,hi�R�5jiuryڹ��k���m5u�W�wd��N݄F��q�c���vr'�:�G	�c���k��pg�F����=0<;�V�y�����i8�ዳ;s��/�m�5��n&QǕ�d}��s��������Co��ό��uZ����m�ru�-Xm�d��F䶆�=_�g��|�p�6�I�Ϯ9�F6�S���֮ʺ���M���9�Bw����H�5�k����huߕ�{��{}ܽ�b��ޣCOƯ��}5;��y�!T����#��0�fNF]���>�ł�ߟٽ��T��v���Nn@�M��}����"&����w�9�1�8�
��>O#/��Q�ʜV��8��ͨ�������d���W�R�:�/G_������
��_���&ۊ&�e�w�&���6z��'k���Ke���������r���l���$�s�f��j��uC�/�FRs�7&!��h-�3G��߰��lA5��5�����ջS\��T?Z&dǧ���c5�5����{烬t�õ��-U�T�l������a�����٧�!,�^�T�\�C
��l��I=��|�ӾT5뚬4/;�Ʒ^�v�y���Q���BW��:k2���҇�����@�1�!���H�Ҟ<���I>�<VL�Ԇ�!wg+F�l�bqSD�fv�wT��;)\�e�n<��Y��K�܆�x''ƸdnV�F�v�n�����!�����e�Fǧf�'��k�.u�����5�z}NNv��pG����̓	��l�5v&\Oo>�y�K������M\��@Em���f+��+��D����CU��P�2�f����h��][��BR㹅O+�0EC��w���1Y����s�|�O�rA'�1e+إ9��֏��^�y��f)�o;��&r����������Q����b>7:��-�k���3/��k@�v�߅�����am�>�j��9�Q�_N�p�k'6��A�=��f藵ְ�2먋L�Ų����/���uɺ��u2�u/Wm�/7�����}��u��fh�I=�w�T	�5�ˡ�_~�W���0َnf=��7U�o���/*y��"z�b���.�MͦFuw)��9"���]��og������=����d��E��`�<�f��S�*-��_-���P�������}B��D�x�T�C�{�{�)=��U�l�`o�:�[wu~��b���V������`��.���:�Ȑ8?7�������o���okN��)�H$�=V|���^��HA�V�{f�U����bj-�hvl��;�/�	�]��xE�����$K�����D�j6�rE�_������e`r=��H�H/7ޭ�r���UήEC�5�]��ۍ���f�RS�nR	e�K�+NpR�Xݬ�LU
M7Cݽxβ\�6#NF㱎��q��:::+&�73L��!�[u>�����RC�����r)�W�P��{j$���
��ˋ�;������Q�F�b
q�^c�#�܏���xM��s��7D����#+(Meꆬ�)��zc�Sf�i����y�(��-�ЎI�U3�������B��^]��[�������������_��g�1U_t���-���3��p"jEMC^�{'����Eώ��J
o��بg�1�A���ۉ�
�5R:>@?z7��s��鋜0�Г1�2s ?eU�[�+�)�;�m:�|n�X�s=�p�F�n]O��B��p�뭳��kv�S�v�F�z�~׵�G��pj��!�ؾ�d@d���r<ݳ���^�*�JƎM���@�^�赮�ɽ>�^���t�s���ǯ.Î牴�~���Be���}��
r�j�L����Y�7`����ܺYݴ��<^ѷA�9,�IhD[*cr�σ�=��5���D������da����&�#�͑��B��gE�"�$M��K�2��b�a�۟�mߖ�5Mw,�ѓUHC�y�ȸ"�\�[�ӗ[�W�,��ƑU=�mvl�p��g�\J;2}�)Y�di8�V�۞�~�>�>�^un�:��<�d8G
�U�Rʝ��i��r��s�D^���nP,V��y6/����	��ʅʾwؽ�8m�g���d>���r���)(�5�ζ�B������֗�S���L6�juI&�Y1-o:�^g\>���H�v�!{��;;�c4�CS�|���f�b���-�>�l~�Y���)�P�8��yo�Ǒ�� �J�d7N��Ѵ6��;3c:��m�+�iit�;q�)�}>��?���ܿ!�@V����JKYcM;c���>���F��7n��7�~ϓ[o�
َ�'.���E����]Ǝ�p�l��]i<E���\���z�N�:���|f�V3Q�q�`�m��oW'&�����!�n�D$���ۇ�Sw7nM�vuB��WPZR�B�D&l�q9�SǾSk|���η8�.��m�Y/�#b�T\�;�����#j���m�=b���̯`��F�M�e�/<�7<X��p	8!�M��'_�v/�Ѿ�[�3��quqFȇ��u����-u8��Q응Y��V^uן,�C���r	n-�axOu[4.���'�xP�����ɺ�����s�m'Q���ܧ��}��]�����Z֬nI�H.BԐ�ܸ4ZV�x�BB@����ߛ�m*�L�/7�u�n�>�&tC����>��B�+O�A0�P���z7/�W�����m(�ȍ�܃XV��v���uﳝ�E��޻lH����3�1��=Z;�2*�W�w՘xa��6�÷������Fn'�L�C�!K�[�3��w�u�9���̒^z���oD��S(A��N_3*�� �g籰�l8�ݻ=e�;X�"귲�u�@T�3�7	8m����N�f�{�Ձ}�o�6��y�����+���~��R�/���,�4��cUXZ�A��{������M{��<8����̮2U����h4�S���*�Q�K�0��ˠr�&|o`���4U뻍��l�S�!�n�nM�O�E��Lw��K}�з1����g]�G#1��S�ѝ����3����s͍��&Yi�(�%k�;.�{�w�c�/�#>���̬�Y>�R��_�(ӝʾ�k1����8��ڭ��!g�fdrf�A��}��/�����^+��wn92o,�:�"w6��,G�s4�'kg�3�,�my�Y��¡�6�N!<����ߒ��+?����"�����V��ȳ��C�R�[�����*����/�>W��+�¬5�ac�>Cc��'��ٹ�K�Wpd臢�p�;�Սv�(k�
0�l���Q�6�gP��W���NK�T��.�]č��XD�*S��9�����Y���㘱�{�cm�0H�D�;;�ܥ��M�٥��+ ���叧w"p��J/�z����y��J�az���<ƨq�L&�]��L�^Uo%�{�Ecz��m�����X�<o�����Sە��YPfb�/�ݬ�I��5Ł��*��䨵uJ�]�nKTߘ�
~��8�^#���%7u�y�],�eYZ�d�w��s͏��lպ����2�]ڱI:��Sc�+&X�z�_G���˷*��[f
<��2�7�}��A���W�u.�ۼ[�D""��c�En�y����베T�W�wOi{�Bx�Q��=���D0���I�K(�T��p������-�V�s0Z�z�ʈS�&�Րݹ
�s�� �љ�{�v��fӡ�[.w�j��Hʶ��3kl-�+�[Y.ƾ�^�
�{"5�# ��1���Xwwd0N�&�Iv��A���m�7(� �t��ݖ�J��������7��l1,��^e�оΊ���~�F���2j��^.�������Ri����֫I�woTn��a7:�y�xu�tͽ"�b�[��Z��yR��̽!VDs����s�V3n����g�:_�1��f�ƺhy�Ŀ�v�鳳VL̢J�^�i:�����l�G,jUհ-�X�e�xv�'�=�xm��l;ʂ�v����:*R����s�*��՜�Ε�N�����j��u@��!�J�SX�O.�M�|�M<���Gh�NV�:�H�RS�X���P͕�n���9V���^�%O��:.`��lD'�׎6-�\��ðu�[�cY���V�
�WWJ"��:��[@��m�ے�(@]����CQ�V']�I�]l��ߐ�]nz�..}���a�L&���;o�\��9�|U�1����t�~{ �.L=�F�%�<u�e:�D��S�/�j�E�|���p������Y�QEOt�e߇e��&���/��a\��^����.|o|������L�>����9s��W��-Djr�M`���l�!�8�g�[-;]��G�B4���[�sNnQᔵ���~��?��^E��~��_z:��Ұ�G�ﮪo�� }5Y�r,O���o��D�ݯoo	��r?�^�EF�1�cn=�����3����U}=�V_��z�bDVEEWn���Y��:o�'��yh]������V6{]��|N5#
�)�k�w+�}�>So|5l�e��qV�p��.���/*��n���Z��#m#�F2 ��nށ�'������Y�������Mh�)�o��^B�����U�������zw��,��WՋJ�cP�*�U�{	���U���k40/�I�=���y�-��^gvm��a<�¹|��Sٹ7*��8��r���$&F�.5�Uf}ճ}N}����T0p��O_Fz4���M�>���g�^ע�6�ϳ'��<�ߖ⟋F$������F�q%n�ٸ�1���և�k�Y3�a�,�..3��aC�o�^EOk�^���&��Y����n�{`S�6��_GuE��fǒ��f�Y�.Is�HÑĔ���x9�5f�$sIg��u~�~��t��K�8*�����)�,��fs ��h.�{����m��JJ�%
KN.g��u3o�c�Z��*\ŕ�A2s�mU�fb�8q�z�龔��+��q06l���
(�aLCo�}�^�m��vy��cӑ��J>�U���Q�>.Ѽ���������FD�쒨�2����r"�;]���g��Z9�{;9sz������u���a�S1�]���=�qh._|�����/Rdo��Ԍת��4�D���V�Y��!��m�rݑ�li�1�|	��� ��Y!�CsL����~�����YSG+*���Y˭�H5�^�Ae�f��"t4�����_N1q�j;vV�7bx�S^�&������7	Ć�/�=lm;c�l�p��3wh����n���\(���Va�J���&!��60pF����;��{v�=kMä��u����9�r���]|��8-Jۮ��t�Ɨ;J\\`�Κ��J!��f��a��Mg�{quMc׀�۷a<��W�֝�ZIvw+�o�z�����t�b�Z�a�"��O���I���j�R�
W�=�y?v�7�sr���R>��\9����n����سv��Ͷ	����S���p�ò��7��ev���t���y9~�m��V^���Aon˻��U�r�F�k�>s�����5�ӓ�%he��!�_v�I�I]�nlÕ{b�[�;�aؐ��B.z��5�kw����«����$N2[���Gz��^����;��jo"�;�"��̎��1�������7����Fb�tc��Gm�*�PHPQ�"�{���u�k+�(���T��?s�_��=J���Ǎ�k���4�n�O�F����<�9(r�N�4�נ��kf۩���L�n4���z�]YkJW*n�8��UT�Q�i��{��`�z6���M1�e[[�yrN$�n�ᘜ�a^��+�������P1/oݾ��04�%D'��4}&�*zu���Wټ���>ǌlJ�U���EU��6��N�����w>Cj�cU�W	��]�i�:���6��x(>��M�=�G���gfdM�� VP=Q^
ww�ۢ�u��!��6{�^�l����#0���7�>]�^Ϟ�:��E��u��!ݞ�u��;�����������#��`n�~>�����O�3����\����'�`5(��>C��8p��{��7]m���oir�"lE�D���)!�n�%;�}�^\�z{�c���5Dl�H�-ހo/�G�䊽q�
�uЦ��z��
<������~�F�vG�G8�ϋ'n�����[���ۭ�u�%h���z�tQ�؛�����������-zO����$�#2C�|�cxZ#��������[,ߜ��l�)hh��b�192�xa���~|tv�o�hϹ����nc+��{݁	��L�M;�����?<Vk�~�B�<��)��-@ܑ폟��
�g�[�
u�W҄�,b�j�X����ծ9\�t?sσ�4����ka���e��p*��]�o�̒^#U�.`�僼��)L����u�:�70�/7��޵��=t�lzaa(NC�{K�~��O�kئm_yx1^���S(?s��yﯦ�f�����bk����{�4��\�������Ų�i���K���Y���VZ�;�F[b:}�l�[�����>R+�5w�}�{���7�92q���T��%	��ll�m��՜�0=�m\� +�붝���J�e��v�`���V����Ϝy�o�y�=jn	��N��n�ș�5�}���8~���F�dw�_2�L(i���<��ToM_��7����t�w��h����s��ҟWZ��x��)���>�C>��4TIț h۝�O���u
�d���{vu&_��eO�Rǰ��lO%��lt����>U��B�3)'7hM�x��u�{m˚V��WF%=���wff���/g�m��}��~�U�sB��dwmh��!�Ku�W��m^��pnw%Nڋwm���������]�����m��z+�ww.З������s�v�u� 1D�r$�M���yw�ћ��AY2a��f
�,�:�	���؅{!}���u:%�K��c���MV���y��D�3k���ޚ�3�c�.�͸�v�X�W�d[�ў�͎'T~���ʽ��v̟�S�o�Q����y�ۧ�����Vb��#�j�7bk!cM�}k䛄F�i6T)�[����e���"l�ǥ�#��qk���0ͳz��=}y��?EWypʟ]q�z)WU#x����M�N2��:�o��k�y2������A�ܡ���/ߪ��;&Y��V�s���f���d[t��ʁ?�8,����=}�x6����w�	���nՖ��>��3��o�{�wT|��o�oӒ��.jk3��)�
*T�����7n����0�SX��Z������qL��ð���W{�"l�V/vĥ	��<�8e��.�L�A
G�Ǒ5Í������Y�k(��c[�@%�����T!�\X���؉ V��Y?��U[T�F�QKqs��������QXm�h7�k�_@s+з nv�|,��Q<�V5�g�&Z��nޏ7I�;n=:�K��t�{ ��s�+�u�<pi�p�>x�s]c{;�\�"+�9.���B��{<=��0J������lF���;�q�Z���upf�d�.z�tF��8P(c���Uv��⣯-�j;dn:��'����Sv,�#��Ay��^�C�ug��%�Z�=�0��5���Y�����K�����
����۝����<��Һ�^����/M�7����+�06�m��M̾�Ī/�c��n5e���w�����r�P���gc</V��t�uQ��`4�q��Ďs�(`����p��.�^�ʵ��_�xΞ�>�=�+�}��o=���Lq8�l�����.�F�G�и�n��H�W�/����o�]~��o�Y��xP:g%�F�j���2=N1�
iG:~~ʎ�>��d��ijL&���2bVoWgcG����c�v\Pۺo�N���fc����~���^K��gd��(��#E4��l�{Ia�Y��.{v�mս8xԠ�W6�W��2̤�4�FJ��{/z��[���k�����Í��I�55v��_}r|v;k޽>������
�H�N6�b2rmK[�c=��~9��$��N`fBc*D�ED���Ҥ�ʗ��et�lV���F���}r�0.{�(��B)�qN��qI۵瓘�ڶrg��zb?���h���7������"|�^��\�4�����g�������pTu�
pߏ�!>ފ6���^�WfIw�����Gڵ��^F�W��a�+߹?��K_�bs�G�-��|���0�$i䕕���Gۜ|#��/w=/]qq'���B��w;�fz{`�h�������vÈ���:���nI{�ξ��)}��AQ^�d���`(u^5s�z{��m̫ON�c���f\s{JA̹�I�z.W��rw]W^֯-$n^M�Z���F�b��˰uu��.k�r�c6�����2�����s�Ǎ�z��gT��O�7�=�߅��1�8��n��(T�8�R�TsL"ى�-���H��r\���.������N��z/W*��\i��\��R-V�;y'�$��)F�ݙ>F�Z� q� ���mHp�m��B�����1w?]|8|�5�ėQQK&��o)�[�n�O��8>J����X���Ȟ��d^�(J^��=�gL�^Np:Nun5
��}_��g���Ǿ���*}p��9N����G"A�4�o/3~gk���w���۸����>�k�Q��*����8��T�^Vza$
��N��(��co�������S���Q���Q2�v����U��o�gm�6N��5�J�Ϭ}w	i��}��v;c�:�n�vl��������1��L�Z�ۖe��[��P���������n�ms�lS
�nl�gl�W�����".5��.ҩ5�_	�Ȯ��ݹ��u%|
�MA��=JR�f��[@/�����i�PT+�Y��s��� x~j�L����{e6g�)��v�`n^�V`�_?t���$��S[��,�6�{$�����{���u�}��|h�R�#��0�P(ܒ���{�u5:�t߫�֯&�׫��6;f�'k���4��B�9��@#M70Ur*m͹�ySED����X�cqTyG�˫�}g�^�k �9��;;��38�l��V����wnr���q���q�vB��9A����U�5����eH����H�ׇ�~����h\�y	��v|@�x<�wo�^ϼ�[�`�J��>�������^��7,���[�-�fIT(��w���ېu���d
��Y��4�8���U�XNI�6gv��W��"����zz���k�ؼ���W��&�_�8��eѫ��Hn��]2����(ɂ��kһ����}���Ԇ_��s�
��~ֶ�eV_�����pL�9Gw�A=Z{]`��h�I�8�L�#.)ppyO�v,��	[�ƾ�U<�v�;�����	7�R߷7ٹ\��O��$�-�I�(�2��%�7��8v<�:������x���R�a[��7�+w�7dܙ�ok�T��h�b%�[2������闿�����f�aSB�G���z�.��~���vzcbxսS��\z��{����Q�t\X�fg�	�喰��h$:4Y��l�A�sA�g�(�[&�+2�h��o�b�n3h�7F��Be�3���{��:�|.�:�IOX�x��z��O�kJKDjʍ��O�Cu�Aq�� @��g6�Q�5�](δp����t����zE���ՔE����oG���v�=wי,�@6/����j2ir[�mu/�j��to	�|	g{g��Y��M�vf��1Q�cK�r=p�e���¬��'wb̎�����P��Wf�Y�Jտ�Q��jt�^v��}(��ܥhP�4���ջ�T��Gm6��!S
.�D2&+M3�����+_s��_]20J0^eeofQ̓��(�~!7�K�C3t[�;�/�\����u�ww�Ϟr���:�o�x^�0+����y*m���IM'nIю�|�o�M��P�թU��ଷ�R��aIL��5fۋ1���jtQ�y1�s�7(�ޖ^���,�c��S��R�Y�z���`��j��!�	{F����$l�V�]�xp�L���+6���t]f⡜��G|�y�׬�'if�60+�dޡI]?�S��9v��+�xY1p|��o;��b����Ӿ�U��:�j�8�[O��$vI:i�"��.2�����hv�bݙ�1�����6�z�T�� f@f�,dD^��/q��*ݼ�k�zA#憠��#�{�su��c��3*���o���R��A-�Un�G�\�F��d��%v�����FE�)Y��UUUOcMR�#UUUJ���&U��B��ԫD���C�ɢ0�J��@gb�3�;m*���ۮ�س'/"u�Ů��Vrۘ}w�c}mӡ�=�eV%;Gn�k�J@��Ss�T�G-�X���*�Р�?���N�����%[�;*t�,��q�����Ao5��������l���������'vϮM��j�R�&y��;h��a�7m�ZF�Ku�$���	����J�7c�㵘��N��ڟN����; N0]��-�����rq�Ճ�#WW�9�ixt�S��lm���{o\{s2q�ݷd�m�zq:��<��V��ʡ��ݷ���e�q��ІL��Q@n���m���:��{q.����c��Q s��d��������a��:�]g���v�=���}o��u��nw.ys��a3M�Gd�mb��zI�ur���P]�x]ve-�=��T�\�Y�{J<m��Cz����u�7*ov
��ט=Q�> �[���:���9xEM���S�6;k���9��;�v�[�M�� ��+x��7iz����1�˻�=�wfzg��۳�
d��6;�\i��:�lIۓ6��Ɲ���ok&��w�t?8�ӹɗ=��s�9��t��J��7k/k��/rcF7<e��n5���:�M���������ь�õW�h���yϏ7p� �6���N��hK���7[Q� /m�}����zA���r=��v��布!�]`ݞkz�ug���2������CƷ]�i����u����<�s@q�t�1�N20v��x�2Vl��3殜�nR9���S���;�z���k&�� ��ϲ�ts���5k0v=���l�����nاa�� (�n�����|g#��pKn���`G�#��ot)=vn�<f�/!��<���������ax�\�8�P��%۴�{\R��b��2co� ���(�/��gׇ;6�ۑ��F�ƹ`�!iݪn���򽵳�����#m�>��~F
%�
ym�
�C+�����v]�s���s��N�2��ݰ��yk���y��pvԽs���e��\c��w�Wj�ݙܽLH�h5#��
��Nq��7'<���ݷ+�6jn�v6�:�f�f�d��s���v�a��)�0�O-��l<�����.�8�=�E\�!_�����e��;��X�f����M��!���X��,|[;Omh��:'��V�m7b�nu�Z;$p�ks�\�R,�'M������ 6L���zU؍��Cw�j޺5�cD/��f��yUOy�Z�+���s��m�\1ɲ�B~ﾚ���}M麖j\y�T;΢��>���U����X�)�ޫf�3��h_6=�qQ���0��- ���{C�ӵ��9'�Y�s�ϋ� �X�qML�\ޥ~>����/�]��f��y���`ʉII%���o�s�&:�|fo�;#���Y���%8������ѳ�n^��Tq��d���=�1�	��P�!8gС�ou�I6U�v�ш�ץvE��(��T6`N-�:���
.���7��o+�H��b�cy��m��<���2�?X�Y����b#��,h�5���IŹջ/5=�Ēf����W�Rp�o��P_(��ޏ��{By&;��\`�ʚ���V���/�l�����t��|ldϚ�H��(�MEm�vs*^�zψ�,��A�A��8�v���aͱ`���@�ܓ��a���`�3���;�n�c9���}Yj��8ON #pT�����tw�\F�|����Q����'��՟�#���f:��=�j���i.sٞ�L@��؁�%�@�VPc.}�i;0k����A�V�]4�RZ~񶻟�j�2��}_|�,�1b�4;۟w�!l��%��e8{�)�>�:��^�{�ϩ��z�X��3�ٝ'MO8��3Q���C��zy�ʽ��C�W�d6Z����rnE�G}��~��Q����IR
�s���n�&��q�]�;��6��+��n�՜ʝ���'��rW���%P��E�ӻy���u݋mY����\��r�su��D�%��uY-y9}�#&����k��N�3����"��g���>X�+�g������_h��e����$�J����u�W��+����ZE������#��o.�{G��w�u�gU^G��.0Do(���p�%�I�nK�湶���r��S9��ߴ����W��y5X����~{A�
�8����y���Q�m���(��tgܵR��u.�C��&eI/w$@G��Vj���Sj��۪l����߿��C��ٓ���ʖvV}��6��d9$�)�3S�Ϻ�;���xg<΃A�[��}�<jzi�ܥ�m�����;ϻ"��φ{�:h�0�(� �m�O7.kݽ�:���y=�o\KX�m^�o��a��3�q�O6����_��2�DϽ§τ���2O.u��<Lg�������rm�G�.*D�������i���WS�T�_��������},I�ٸ��*C"���������%�9ZǶ��=�G��Yu����\3��MC	C�y�XE����{���Q��NBR�����љ��Wm�l�����<V.A�sӰ�;ׇ��3�=�����i�\�ɐ�U�O���{��s��Ѹ���U��:��z���&z�z���}��	0V$�"�rE�g��w<v��
��#�W�Rd���~�W9/]�	����A7�RY�\�[zw=r���v����ќX5݌�/�$�տ�gv�k͙IB����ru3����;hGۅ�8QZ���ߟ��k���URP�Ӛ���0N.]���Qk�;V�O]0Dxt��#z��P������=�ˉ�^G���g�T����mD�,V*)dj ��E�7C![7h�������qU�涶�n�h�3�Cy�ò����Q�Y�'�{�Tfd�Y�޳Y��Y��!k����[�d��p�=n��Ɉl�)2S�s9�ћNs��k�5���z=Sە�Ǖ5FEmt�z�c������l���<��;�ga�!�C ��E�6�贈#����]\�~�+�p=��z%���z�����W���썭C|�˵:�_5����*H�v�ZEoe^OM����M{�]+2�)�6=h�h��9>��#�u��q Úp��:���v�����c1&R���8,��g���2�d���DD*�q^��f���>�tUGm�]���U���|��ң���mȬ�c"�5ۺ���{�r*��|�p�r�.Z=���:79ۣ��/u4n�;�?����U��$�(�u*�s��,�]�`nk,����߇ߢ�����Sms�aVrλ�4��de�[���oL��Zw]��0�A��e�E<�T�Θv���M��n���v�]�Q<jÚgL���p�۶��ڡ.�	��['P��be�A���َ�i��|#�u�����Q^������]p������oQ&qX'��1s�x�.�`����+�ô`�����|�����b�ׇ]W3��9�/�n�W�elt�svVc$Ɉa�C��{�1~��e�<���S�X?s��	��5�}0o��2�����덫��E���d�¾,C�!0Sn;;{��T��!���I��e׵����d��2Yg�~֦�Ó�����Z`g��a�D�7馗� �I�%Q!�siN��e��[�X��&dEƋm}��O�1S}p��1�w���㗐�ҋ�6����'��%6�����/�)��>}-�tGv������X^�}�{�"aa��kధs#j&��k�2kl�/��9�1fH���w����G�ܝ
��"��y�ݬ��{=>���+�
��U�|�&�Z*|	�F�P1����?gߏ�f��Ȑ�֕8��>��Z�:���d�T�JL�	%Ɠp7����亳%��r}r�&��uN屑yS[]^�*g<�����f��&���2���N�h8�L��2��{�}=�7� �vb�9V����>ɳ��D�Ư�Y%�}ț�U,���n�YooEO-����M�'N+��j�9s��2i��奟�!�j�؟M�{�u7Qܪ�w�zm�ެ'{ϹD^��������а�D�����q��z����O������͙��}+�U������X���<8|/�*^�� �'���O�,]�	�O�J�P��3اE��d��tH�tY���/��R���k�I؟M<;�j�%)���0�ECa��d�"a>�f����v�c��Nd��t�Ek��y0��ٸT�]�5�����z�����m����n���5~��Ҋ���1cn`�@���=C�qt2��+l28[�Bl���n����/>��G&m��[����Qٞ�Q�BcR�Mf�r���p�&!C��i��m��ȗ�3ݸ�>����C�㴷#c#s'$���I��^%M��wnw\�m������n�.��p��0S��qj+e�ų�יM����h���X�ȯ;[+�:k�׺-o��R�����6�Ь����쭹Vz�N���N9�F.�hL���ǯ�۵f3��~޼����h��}}�)!�]W?9{�S��kn����Q,-uI,�{�_W����'����~�O���"L�OC�2os����F���[&���0���6L86Z{��N��;�Z���لK��w�I�� �k���O�����5�r5�*}��2�Sda�%��T�R��nd]���euqv��8SGN�h���vy.BB�pG�a������}V��������|GLQ�lkoLA�}�/}ğ~R势�E�m'��X���;f�+�~�ĉ;��{�r3���0\�{��:����r`d��"�[����E(e�.Y{�n!_k��]T)��<XV���+;Dh�������Ve=3>]�:Ӿ^nAc�h�NGI!rי�<J�w�ƭ}sp�������?9�~�������߲ܓ%��~�,�/A��=�>
P����j�tw.��R�Y�3����6�6���S%�����lv�^=�:�{H�ʭ(�n�d���=��w��}4�I�A�%�n�����Y����d�[/N����BCZ�ӆno�~j�N ?����_p|�j���v}]����j8�h$ˋm����^]z��k�`L�uuq��2硞�{Cm'4ш.�۟��Z&o��st'��3|�JK#�K_9
���42{9�+z�{��"s���O��[!�Q��M�QP}����o�o���ࢃ݇
����5�/*Q�1q>����^n�)7�9`o�v�PP��ˆ`��R0�UݞS9��!��
ʚ��p��O��� �tF�L��;]���Ƙzn��������;�"�0 �0�M��q~;C����?D�Yk��{�yln�w^�u�1+��}eʢ�Ot�}�閽}�t�1�Y].	F��i�������L����&�,ɡ7L������"c��Gw��N�V웮����Lez�Q��,�̎i����s�]Ь���J�RoZ4�/�}��ǻ&���[Xka�$�aV��IB�һ#��"�8�+3a�/�������
�E�(ɤQ��s�ѭQ���2�0	�kv�yf�t���$�́��vۆ�3��<�ݓ��C�u���K��!ǃj�X�tu�nL�'e�����l��p����>�"Og��]r��q�W8z�۔�kõta�;�;:܆��g���Ug\풂�B�מ7��ަ.��TΥ���n��r�uتv�.nS�n�u��ˉ�w�Y9���.ջI��#��^e��3�;����4v�pH8M7c+ӁCF��;Ɓ�H��U�O5?~3H��;���|�[8DU�5S��b�cػ�gy]n���"۟�n�nC�nK�����U��y����/_�����
�7ܫ0�x՘��S|���vq����{���q�q�!P���� W����չ"�ďE�w�+w�R���1��ޑ;��c�m�[ƫ�z�T����5�aBd$8I�~����y|N�NI�w��=��q茚ȝ�y9O6-��`��M�DЇ��<���ʶ�8v�!1	�	��qX�'���f�i����cSӵqW�׿O�=.3����mԬ��מ~5�����tDɭ�+�=^[��ۆ�m�ښ:i��DA��[p+�,��+����f����u��[�����M�[=�Z_�������}�Ũ�x+xm���iu�y�*g��b��v^̢�Ϩ43{��qb&�(���^��r��)�ߙݺ�>���;�p��0�Yh_����*�n%��b���G9��n*�RW���5ޓ��N>/���	a��Φ+�񗞋�O�Ө�CƫkV}��2�%�P��O���s�'��]l��r ��f���Ք���D0Jm�N�D��:=cp'K�]�8�ā�I�{�hzb�m���OAg�ǒ�CE�q���i�1ȷw��#-w��N�{�9�]׎�֮����C�kb�U�҅���gί�%��蹎�g<7+K��2�r4Qb!��!�![�þ�u�G����x�TPʙ��)��n�r�9��ǲ���;�
��9�����_j����s�$�m�[ۇF�鴰�uMi�H�[]����*��`U��o��>�-���}yYd�~�s�ѷ[�S�W�t{�®��]~��	Qq�����8��p�b��Q��$��\\����yof��nɌ�LVw�*�ݲ�_#�T��7�`Ż�����shj�=rG�d���f5�ng ��\��i�Ê�<zv���&��=֖׍/�\�=X��B�Gw���qC_'pe����~���ڎ����BH4[A �"Ob���6��,�J����y�.f�!�7x�eryWK0����4�=����Pyx��si��r�U"�x�����I-o�p�VӚ�y�̅����ro �F�H �Z������3:�
�ݻ�j�m�}E\F��_,õ�ٲ;���-sT�^^e�fN�}4�����'9�8\�0.�ۻy��O(X��C˓�`̃JjY�G��W.����mj]$�O*�p;Ks��T�f����l{Q��2���R'�һ���7V75~��j�mcȳv�2���iԫh�#�f�����*i�=E���w]
��h�j��g���ѷV�A��+o�W8�VK쥭P�5���|��V�f\�r����%U�}��=�̕�u����g�Z�6�7MX�6yK�Ŀhj^&�+<�W`�P����ˬ#�W��6*�h�l��a�����[�2��45��=���yy}"I����k]���X�~��%"���5ov��*��l36��ڴ	ݒ�8�����`�W[J�+�soF�D>H�O"]�K�t([�����a�n ��Ev�et���)+�PZZe�%��=y9S�m^f#Q��JU�a��[X�	òj���mk���эVt�(1����;�",�-B��q��ֺVontY�R7������>���	���X�(�ā���s�1u�
aws�J�.^R<y�9���IzMw#6c�gF�@�G�����}#�o�ӗ���ain��!�V�N�\^��o����Ru�����S�~���m�;+��%,��J&۬�o����czs��\�W'm�D�G8v��6!�\{=��$�[ĶLB	L�}U5�9Iؑ[Y�&T@p ��i�ʼ��(��޸�a�3��w�Q��Z&=�^�;��f7���b.D�u��S����<=u�J�F�M���go��q����n���� ����ocY�ۮU���% ��JM�H��5�b/;�+ jcw����Q���*��L�x����/|�\�_�q⢯z��e8�6�b2�q�c����"��[�y��{ ZW;�x����\[�[��y���dN���.�l���7�Ԣ����M�M�ۆ���6j�>P<E]v�f�ӝ���[�2;��2s�پ�ǿ*��WO�K�p9W{~�}Ю&!6e3��=�=��ɫQ��o�LY&ez��e�)��D�,!�����thOO�����~}���+_�8��#�fv���Z#2����X_N2X�g,uu�G2�g�E9T�՘੡�{>�&�e�-�rL�F�n;�>�xf�S>�H�����Ӊ(u��I�A �M�Ūf�&�o��^aύ�������������;]��9�Wʶ�k�y���B3}���2,!�Q�}[�b������:��=Tr\F�a�VYoTQ�X䭺�ZR�U$��\��^���PE�`�e�7ݞ��ľ����q�Q#�S_Y��Nr���Bۤ�?3	%4Ґ��yY���}Y6��!��=�rnt���Zw}�����w��_�V�����ݪ���/�!X2�є#��*�s�n��uU9��E��f�vw���eG3��Ty4���v�ފe]�����\��Z����_�U�Ao�O��C����_N��S�a�q�q��h�N[�Yw_G�?A�N�%y!W���Ko�2"FD��vF/ �e>������v�9@c�g�1���
���B�\F
�J��J�-�?ܴ�L��5w��3��m���<��������3�e5-��O�WB
��(a��gi�E��zN��qu0�hh�4<�z�q:sM
�!נ���;��G��y�!:vQ7t����I!�f��C��O�����;��%����ps�=��<p����y�D웃=�[��s۰{s��\�*�y_<��Y-==]T�N�ۮ����vúWh�������.����Z�,�ݛ<�VW�D���c��;%��L��j�&�3��"��WWK�;n���J	ڷ#eos2!����!v��gN��+�:u^k]lr[t��h�x��ێ����P�u�e<yg���q���Ϲ[�-rJa�m��0�����!�O~ʃ��fD��}���<��O���"g|�v�5u_��򩑞�9"���<%���,L��n|�I0"LOu[��>l����[���.}��oOzl�>���Cz�Fù��x2(��s�+d,!����U�%U�al�cy�\���=�����{p��FeM?T�W[[�x?d�Uv4�ߗߌ_�#�S����{�=0�Rz�,�Æ�L��"7Z}����3{``�9ϼ���b���c���1�ow���T���;���m��E��GD�~�Y��-��I�1����E���D&�q�T��Re�tg{����B��+�l��G�>H6���<�^���fG�@��cz(���f��+�e	�_eOEe���A:���!���Vu�U��v�j�e%x��r�uwn�ҩ� Z4[��8}���#�2��z��.��vE��r��y���ݎ.�>kj��`]%�1�!{�e���8!f@6~F'QE'�^�
D��ǖ�2
g�c�����N���^�^�mZ��P�������5E�h�v����7�n���c���a��5�;ڪ�4&�Tb���]���F�z�k�Gn��4x�u���	�\�%$OuSg|4�u�o �{~��!/PX6K��@�e����ɏy�Oz=�Az�?D�f�'�WΣQ7��]wBń����)߿�X��{w���c�ڐ��*��ŋ��cb�˼Ę�1[9у��잹
��$=@�O��)�dZ��r��G��w#=Wj{y5��7�9jN��W�ӈ��D�B���Ec@����\�x�/r���>ժ1�0*_��ُc�OԆ��g��!{OYٝ��ƕ=�7��Y%+	/j�N��nX��ۓ�9�{�K=��n�v:�pFYM=���K��ⱌ!��Y{�*�>ߪ����o����ɘ,Vu��N��l�x{�e����nf|�?��8�%DoC��I�Y$��[�}1"z71�o~��\P��3ׇ��I�Zhd���_u���8קw�>�&ɧ|�xo�;}��B ��$ڐ�䛁�߶R�Y��`Ur_����i�,V�cMxQC�T c�q�_�h�Y�N�yx؛yylu���@$��䗷��E0��pX����)"U���S���+k���o�z�2��[}}jg�;�2$E3����j�Qh��P��g���р)��w���m�0 �h�-�>q"��0��ʘާ!Z#`x�`�w&�f{���:+��h%�1����j(&�7�m��MG�Y�7��C�^$J��T��GoJ�9]7.<|�����4%L)�����>�x���* i���Ys���ʧ�Va��%m7�m�ݮ�W���T���kԼ��U�i��q�\�Cϩq7�]o�a�.<��87�[%���H&mS�<�����݄|o��E����W�P�ث�[�\�B. M�!e�\����f(����۽��=�|�9乌�O��(l<�z픧{�xe� � r��y�D��u�����՟�]|y��M�BBj���se�����jo�.�e�C�~$����G��|+�A�cq���Q�}Pa}q��g��^-�tj���w�T����u4[�6��F9	?g�ٻ�1Ko�=X�,c��A�4��D���BȨB�͗^��A�cHW�{�4"۾�y8����f��%���e��yx��zO�iV�����C��g,���a�+��5�b%%R��"��oG.���+%��v�.���d��:Q��e��t�Z�c�����p��?9#��G0�ϐJ���֏O���������3��I#����"ǘ��ǋ��6�T(J("A�}tn}���j���Z��t���*�;�a�����mn;c���ؤ���;�wY���L�߶j�׹W3���F�;>����u�����@���;4��T{���3(�@�-��yYr�Ŝ��gؘ���T$s�H�=�>�����2>[�����l����3k��k��g��؀�2>��5�c��H,+���L��,�AP\(q�n�<�L��K)x"�r4̎<�	�!��#o�����8|@���-A07�F���1U2E���*����]g�h8i�R���c��[1�Q������J#"��qP�}��gr��V���(	��Χ<Y=0�Y׮�|�>WAp�mgݣҍ���i�~J����=�	H�z�������c�ƛR@a�Vy3�`[q�[���0l��7�mĚ�T!FLHCs�K��L����@���t�]J�g�L**>^�.��]�=6�#�no�uV��f��kok�R�*&���{�k����n���t��]��S�b�᮹^ܻ�7��Ч��6H�($��H$mG�2��k �<��k�n����|�ى���ۍ�uQv�(��os2���(UY�z6U+r�ݠkttM�<:I�q�OG��x`g��Kk����;,�G"��j^ q÷k!�T�<<�P[��K��7"]�E�q��m�N�`^�M���\l���W�G�5KM�������a93j֠?ߜ�s�^�c!vN5�4�� ��È�	�e@��k%��"��;��ɐ�`�0��uYc�C�Id%c��0��������܋+@�u�ƾ�d��$x�?^�D��^?�>�`Ko�Z�����A�}�%�b>�}��}0�?o쬡i�<�?hM��V
�]�&�(��a9M�5��#-�iB��?���j��W��Jm��r{��n�
� ��G��lK�2G��ڝ\���V#ؿY���K��qF�@�aD8T0Z��7R���)�� �>�-����� ^b�׺s�+{�B�j\�$~j@�_>T@Z��`�i��=h�����4�&D��#r;F�rc����m�x����0{;��1`'�dSp)mX������|J��wF	���W�*�d�v���iٸ���1����Õ�� j��Ȩ��D������_�_��%��Ib�F(�O���|[�V,�j t2"/�2��~*1�n�c�-�>�YE�qp�Q�.E'���x{��� ��`"EO��Tq�_T��L�Q���H�n���&8:SF:��1�N��\�����@�6^@��q�z����}�,t�h�.�j��H�l/�|F\�d��C^L��?w>��'qپj�z0Sǌ_Ls|��U8%}��p[�LZ�)�OY$�ʮ	�����7�EȚ޷�������[�{T��}��w辡Vy�%�oqfU�5�3tb��p��Z�v���k�]sO������[@T��0��W��U���k�~������s�*���Rd0E���]��w��N����\�=�ܯ� /��٩d�n�)1e�p���s�6M<C��e�2�����b���QAڞ4��d��^����kݪ��9�]1���?x�Ӟ��~ �W��I	�@�be��#g��4.� ���<s�q��tEr��,z z�'ڀң�A�'�l�����i��.���P��A"=�����,Dc.ZO|����,��XL�q?Y����)n�y_�U���:{}{�)�ى�`Ot���l@ A޺sda�l/��@��	~A�L0.�6��^�h�<��1��`���O�/�yݞ[��;��.���%� n�:z�4ڂT;)H�L��|�x^�S�/{ZY,FO�6g���v���D6���1���L�k��ņ�����T���ܪő��LkQ�_(D6�E�$D�m��nI+�c�6!g����op���X�b��1�|�k'D��"zb�,�Q���/z$�x��+V��	�Q ���U�So��B���$�	�llu�j���itG��׬Z$�usWS~��4 ����#ܧ�؇�~���'����b]x�ꅞNax��v΀�c۽鰇.�%�s]�<3��]����>s��AԇT{x��L+�VQ7�\����d9쿺�Ꙁ��K����r>�B��\���P�J�%�-��}�l+DX�KJ�LL
��ɡ�'�����A�B:3r%cf��o�U�3Q���sFR��U+}�쯅�8E�\��~���cp�����S��'����Ǐ9\B���QKa"�W� ����4��������DZR~!� �EIÝS����ߥۀ��A�K���0�VUi�t�^]�ǻy�w��	�}VEX����G4�_g���Tn.Y(����D@�]s͢�����U6�[u�@v�%���	lv�"-��j)��xK��Y ���fx�ݞ���굯�0(�� e�ĆA�IBj~#����~��m���BCq
 i[�r��n>�'%@'�'+��M^�[�s��UE�LB�� Ȳx*ݶ",����?Q�H��9�1�v��.�?\MQ��8~4׽�y��1��QA��Q�ԟ�h�<+V��A�]�4*�vIfp��(D	��sB��R0���!�	=���O�C� ����7��.2�	E?�_e���4�*���ף=^"�4�4�,�T�ξ���%v*���Y����j@:t��#U�8�A]:�H3�B*����U�X�܇�1H|L-�1�~�nCf-׵s�	Mb���Ӎ�35�Yծ��۫�O�%w���]=t]��cU�
8]X�3s���:]g}����e��wgI�_�O�\���R������|0�HP��f*����nZ�[H�ч�(	-N׊��tn��G��u����*�&�U"ѩ1K�� ���ܤW?}������[1�f��E�	&u�c�ƅ�=�O�צt&��U���&�N���=����OE�筞�Ɏ8�1`�ڑ�i�Tj�D�V��~��X�Y1S�����r��\D�L&��
F1�1����#��^H�W�3'�~��ꛉ �H��][�r����*_T�k�k��8A*a�楳	gz�"94�CC�ʳ��%�K�Ls���{��X]>����ّ�|(����i|3*�H�W��ɶU�-8s�:r�M��|6L[t༬$
?�L�?}g�5��;=ao��:g�ď�*q4�-6KJm�E$��	pX�:�0�a7"��z��K�Z!?k�4� ��N�9�	6G��q��<�$	xKB�6��,��11��2c��L�;�J�>Ⱦ�IpX�7����1��"��g	t�� A���l��5�@���>�� >���%%�*,_}�\�-
�Ʌ��LXƧ_�yA�.����.�fanp���d�����\�����g��b��${Y�wؒ�UU��n�1�bK��S�/��v��-I����չ�}?/����~�R~#�� ��{UmS��*Y��_����������_υ�����0��<�T��@��`"����D�����@k��m� ?ϼ��b>��W���!�����z}>�^w�t��*fQQF �Y��U�"U8e(����� 7���|5!�.��O���@m����9�� 9x�҂���M-�sז�Zڐ���:p�mԄȄ��۝����o?n:��l���;���p�|����e5������� �s2}p ׾8      T�(
        � �       U � �晴���BJ(�(��JD�
R�"�U*T����$�%T)E����UP�R���T���RB�*��"RJ")R�JRI+������=5J���j�wi����ƪ��
�w����Ѧ��^a���]m
�{z��B��T�:��\mj��0[h�ڱ (;�����É�
+�Q(���V��z��{z�j֮���K�{z{Kfw��C�^յw�W�mV�u�ȶ��צf�y��T���(Sl�U�*UBUT�H��H��[Ur����y�R�R�Ƶ���ڵ#ު�޽�X�Z���[��E[*��mf6�����SMވ��ך���=歪�y���P(PB�C[W�WM�mw��c[l�(���me��{��j���m�����j����l�p<�W{٭���ci[�gcZ��΅�j�=�Z�چ��
�G=H���*��� �TR��)E"�\��QG=����(�3��S֏=��UQ�R ���w\u�b;�:E锗zܥ�ye�.=������s��Ԋ�fD�*M5QPPc(���I֫�w ���D��D��v�겕����i%��m�'�˓QI%N��U"ނH��r�L�J�eJ�l����R��qh���aJUz���(�
I"�%*E
(��UH��ܞ1�U.YE:��=����w��R<�D'��EU��JIE�r��R�۪�)�k�n�*(=ޥTU��W&�T�{4�&I{@�@��]뎪�^Y/=�)(���!�)*�Lm/T�UGyܢ��I{�:(��+�h��8�JSzE$U[�T��Qw����"�y��U���QQ(y��UB�/x%D�$�)@	J%$�EO="��.��y��I޷����W�!�3-��t�1�<<�U���풥.��^,��x��ڋmoz�JI�yy�)B��2�\��.U 
Q w�Ӡ�X��A���HD��J��]��\Yր�z���4r�K` �$��� sy� �= {� i� �:=��; @ �? 4�* �T��
JUA�` Si�zOTb~�  3*�%J�41�j�I�{*   4�&�*�@4 �Ț��3���)� E��I�&&�y��ֿ�*� UUW@���U  ���(
 P���U  ����@ *����P 
��5B�@P��"� *�
���|�R/�g1�]�8ƙ��o0�/!uv� �}ע��w��Ŝ�@�$�ܝ܌F��==����o����O�D���:(6���Ŵn��.�Fr�2���t�Gn���BK
v����*<��;�o��b!��wx�sSq�.�ܯk2v��ʹ@YoI\b��nd��j4���)��k�q��c���*ݫsl��WY5wv��_!u�N偾Z[���Π�gu*JsPԐ�9ܛYn�Ujd�.W.7�n��t��^����8��0	��Z�'w��[�u#�mɇ#��X]��c8�{���߮j!�y��-���B��ٸV	���M���\����z���8]�D�uD���yk�T�����
 ��c_�=٤���E�w��Qs�8�f��8-���"�RS8ot��0�淗�6佨o!�!J�Ët�-m�&������GK�YK���v�T��ݗw�6q7N���e���v�ss�W�c흠M�tot�v��c�s9�'���P�z!;I�jW;�� �U�}�l���d�G��Ynu-�� ���]r��fܸ��}GD[�l���c�	�\� Zl$��쯄��3F��S7��Z�<�3GQ�J������n�:&���m� `O��4�6gjx�K��/�;�>����d�n�@���{I38`Fo1��0A9���k��T�M�Xͦד��5�њ�f�se�Y�n�鶒�c�FiWG$f���a�r��Y9B�Q�^h܋+��a�����a��r�~����5E�����#"Z�r�\C��͏�ɳ�k�����i��צ�ꟘH'��3&k�AZl7Nѽ���pDp'�l�;����Xw{szTfLAhg���gdFj{��"�&�ÓCZ���u�9n/e܉L����{pn��kp�n4
}���N�N�x��om
��󫲣�^���9���I�d�kV�Q�6�m�\��8���C9���ퟟo\���S����T�br�Obq<yْp�Ht$����8v��]�yo-o��9v��ν�� ^�_z$Ms���7�A(#�����;gk���a���<�9�;�F ����1�	���עqŽ���V�#m�&��ܹm�z�:�p�v`�y�)`wH��PC앜��٣�j�x�~K�ÿ�N���V��M�@�4�Ƃ1G���.�Ժ؜5˝���	l�	��k��^���n8�طi�s9�i�3���釕���fuy]Z5���iz3g�Z.��c���~.�Ǐ�F�E���<m�κaG�d�ڐ���״#�Ɣ�F X-,�wZ�;�Z&�q6�3Nv��z��Qz��Ϋ��=�Щ/����$b�1�ɡ�
`�����H��;��孌7�ˁ��-ɖ=�٣v���WJ�WF�"܆^������z���]��=���M�m�F	�g>M0�^1fdݷ��r�&!����"6��wk����"�;�ŻF6�f���+w7.��n�Լ�҅��El1bָ�� c׏�����8��zFC7������˰g	΍e'���u�۽�vqH��E�UoB���f��z�e�wn!�P{xU�;�sn<w���N�'jo(�Kc�v.9�B���'�nh���� � � ���2��\�b��˛��T	���O�4���Y��1��n���Y�&�ڛ�i�Tq���Ü]�BKl=�tÒ�@���h���SA7�g���f^d�v�z�᠔N��f��ʆ{O�9�#�d���g.���7Fr��yBrc�\�ُz��`�@ԇT�,�a�Ga֎{9�f�+RB���.��Ҡ��[7�����,�]yE(+���;�ܠ�Μ^:.�Q�ѣ����RX�@��-���l�ԍu�*�t���0�чⓐbv�����nrc0p
ik�b6���lQ��4� ���ʻ�fLF9�5';�ե`�u�+�&�`���4�]���dW���YH:7l'f<����9њIto"��&)�Q�����sg���u����U�nk�#��\�����i���8�*R� :5���	<"�{�͖�}Y:M����f�p�Gty9�c��7:Iʪ��� ��H���*�c�:���d�ާ6Q���O��s�3�v�W�Qj0��o-=�}z��é���<�BoQ=G(�¢�squ���tƣ�reS4q�=�S���)/
+�vWs�M���w��>�w�ej�F[�5i�F�1��g~�
�o.א��JӠ%t.���\��9�٪̿{�@s>�	��Q���Kc�\�,d;�˼��'MTR.���iq	���G(e?�SB`�o	_��Uǹ��IL�5�EQ�����މ��$��ʒ8<CC�� ���Y�Q���Ù���{�j���Ž6-�E�[9�b���a���@�ר�B�^�8W�#U��.^6��x�^7K������L{��r,��}x!�Tq�N��;�!����F���,��]ZZ[��p�m�fk��BV�X���ӝ���)FM�.�^n[݋]֦N�.��/�".L��R�����,����I��c�j�R٫-�i	�;4i�̽�[��ܟ �����ޜٚ�N�Y�ՋA�:�:Њ��V�SM���ӎS���eiZ&5����c�%�R«hI�9�5��kk�HǗQ�v��\�޴G��z��ǒ�t6.�O^ !BG]�Z���ջ��1;7odq��9�~$�q��xM_���]'[ޗ/�/EeH���ϐi�7��ްؖ}ڇt5�������D�׃f�}F�������*q|�q�uE�`#f�F��S4��u؆2���}��z�)@�&ŧ��];	D����4WMk'6rD�;�y��n�)H��g�T.H�Eg��s,�,S1�4��o{�'�v�I�~�M,s��sNk4�ըB𪈁�Y[t]��rT��۶���w��������ʷ+���vtqZ�����X�,�lF�5'+g����ۅ\�7n�94>�����c3f��dC/cf�[�Ś�s�{�7��e����wu����L��Uh���Iʞ=_a�j�{qc4��fz��CG#׆�,m�+��))_�9V��5�[�۹m�z�)�2� JO�Bܜ8G7:�x`����D��j-���t֛�d�ɉq�c�68��vu�������hGQ8�tuPHB�U�Oh0&�,�z���T;ݱ�ާy
v��v�>�F�5&��2M[���Z�P�#�KiӮt�}���)YM;��u����4t]����Y�Uk;���f���nh��j��F��K:f�0M�u,_����:0�v8D�Q���ޯt���A� ����nn�+��ٴȲ֦���
��Z��筼�,�#�3n���ת������9�^
�J M���0�Yp6�;�7tw^�\Z�X�D�f��J>�#�˯��IS� q
�����s��͡w�/��UU.��vrwFp���@ȹ`P�"z��.6��r�m 4��|��oGc)o���P�Ŗ���&X��{��b�g7	��ncKj�q:���D&vr�����%Q��l�:$��s`[����g�US��\��l�X��/�tn��D���b>,}V��[gh�.q�nn=wk����,|�������.1�V��9�����!#�égwelZ��ǚ��\��A�w��0�y����v��{e���f��]�lї^]�q�t�Ve/a%�J%���� �M6� M��T��YGy
D��k�^��!i���9�����ƊV9%�q�3`iZ�(`l�ka�&�c�Ժ��D�C��
�U�_W 1��r����6%���fhȴ��=R�3ecF�J@9xɕ��;��H���D�v����U���[�m��r�PKWH.����νs	d��v%NwM���t��l0s�cUb'H��f����z�p=W+:�bCxh�"[��]Xtp�ݏ^�Q̴:vw�gt�إ %�N��\/,�]�u�	�j׈�/J�0K9,��B-`k�M%�Y�sK�ѻ_PA������(�%[�;e���ʬ'e�n35��]Ӝ/���{5DAa
����{;����v��Zm�{��|���0�EUJ��vc-nܜ
�,��[-Fn,Y*��ye`L4�fm�Nm�u�ƜplIK��1�d��`.�T����]ɣ�n��Z�����sLo���di�0r��a�5F� 6�DWI-�枬��t�;v�s�I�_*;F�0�K��� ���K�ҳ	�ҭ_��£G-O�4�g~X��������q2���a�$�/%\����Y���!�����p���ZyG�T;�m����I�UùN�x9%����$���ҹ�z-�s�bO�Hӛt��F]���'u�-�4�0��>]�j :\�69NV��os:ڊ��4W�z�SM4qYA�T����.�����7��G��Acv�eV@��\\S�^&]�׆q;�{sP�N��l\r䊌U�9�8���\+�tN}�SV��i�����,��:���a���ɼ�b�X�	�8��ǫ��x FQ��_c���QT�ҹ1�\�Ʒ8�7��s�:�+�v2�%���o�<b�L�1�d뙫op�x���\����e8�Z�܆���C� x�ӌ��w�;�5�z��u�xpL W`C_5��Y�o�u�g/	�M0\��%f��J�G qCi�pS�^@��4��� �y]8�3�T-z�.?�mC��cy��[	c�j��w�{lY �>Өء������n��]���&�7�ky�"�0tW$����f�⏷z~��rJ����H!��@�%��sK.S�
e�P��( c9ĺ�mI�q���E���MSHaC9n��WP���n�A�@��u�6�mOq)!]���#����C�vv'P�nE���Z,���/�s�JQ��2���
��qð�]�̯.&U�ɻH�������Lxm�Y4^a �Y��b��~X3\xq^�&���otld����A^��:p��DY,]�e�k.g8S�^%1P�:Is�Vt��Q#�W:�е��f�e��v�و���p��x���곲�"Oe�.��-&I�X�a�����e��;�i�Ous"p��[�*��]U�Vmyk*^��W;s�u�xbL\!'Pe�ݐ`o�o~';!=
C�jpf�
���[�r�Ks����;�����Z|xvI����U�;���{\��[q� ��|8���v�D��}�X��p^����<�vh�<.�����I��+�Y�.m,�0�H�� ��4YWr~�*�l͠�40���/p���'v����kcp�n<'J���yU.hf��Rgsi���
�[U��F�[��+�l0&�v�N9ߦR�ٷr���uիr9F����0M�I#$�6�:u�(���N���8R�����"{]ɧB����8���7��`�7��3c�k݂	9Q݁�{�=��|wPog^]	]�r^9-=uH���eYka�CP��3�ҴCX'��; [v�n��(Td�/���AǑN�Օ�tC���-���{�N]yu����t-���ƫ4�����j�x��m����N��VT����9���Y�#9�N��}��yR���h��X�+�N�Rܸ���FKug$�[�fv�;��8E��B��t�zgd�EM�+t��V�=�w�����惡����i��ԭd���æ�����,����I�e�9�8�{9b]���.p{p���1Gè�V&��z0��c�wPݭ%�+��[��>����m��F�n��:������i�±��.g�rx�����w�@L��_=���sxf��\7�[��c$���ዺ���C�v�d;e&��ǳ��sL��sD�P!���q�&�-8.�Է��1̓;'��r8�0��͑���.�c���y5J�j�8i�.�mM�X�κ�[@�y���Ţ��Y��D�����cg.�����	=;��1n]W9��㝼�ˏD���v��٧O�.�y�G��h{6=�Ժ�1z򯡺jdO�O'���D2*c{�3�ؒ�7��@��bh�f	o#;nnp������GT��;;�h�M�ˁח��{7��q[����)����N��_E�LHR��>z�.ٶ��g.[�� >ݱ��-��I��	���E���H���NS*��Ȃn��u����*a5�·Us^%{v�2��N$(�+��k&�0����P�2ѫ^�E��v��(F�\��w�X;Ӆ놶�ͤ .E�U���N�.l:{v�:嘴��G�y=��a�(�6�M�3]��3�z�=�΢d�ۂbC�<J\����;AѝF���ٱXP�)L91g-w�e����o�飺t4Cf�KsW^�{
�^�l�1���U����׮�9�sK���{��^v��(��܈#.�{��������a!�O�X�v�Wq_ݦ�)�h�{���$d��_�#�gі��f>��o>�C��:4z@����˹�3��i8LvR�~ %�j�o���I��'���H��,�Dr�D4���(���IƮ�зt+��OMGe�m��mB���0��Ƚ�$<����Ǡ��iVat���_�뽳@�n�i�a+'N�y�y �u�a8��9{ym�B����bO��5B��Ǹ���������*��UUUU+UUUJնʪ��)�+j�hV����`�UUUJ�mT�UUUUURV�������Y[m���������UUv-�j��@+``n4��\�D���4F������rL[�'��v:&l�AP욒�hQ��Z!�^�HG�1��6Yy�GiaR�1����8�����P���%�ńk�ѰX�k���vػ�"k."�a�ͳ֨�/��7iU�׭��[W�@�2��K��� �MQ,�%�%]������ې�9��V�%`J�A��]�ʛ`�r�Dލ�����|�ك�;��v]�W1�.mV���}St���ш�eAt,�[t1�؍c;{{gr$�c��q�癘9"wC�m�Wc�pL���T;k[]� u�M��wm�y�.��J&����E�tq�q�)�y��]n36�����q0<2�Xf�Z Pu�]&Ճ�����*cssc����z�du�9�����X1����ݸ�����(؎:=k=IX̾{T�
�6�	��:)�aY-�c�h�����i��9m�;IBa�l��4iQ�g����{���ǣ�X´]#y��z��s�V^����Q/9��s�����V��D�νHA�s�z���ac��r��@U��K`)�]��R-��5:\�XK�=�Hq������	��������B�m��,	u#Y�m0f[+4ٶ����|���
nr��c�k�o+���%=l�g���ΰ�"��;}�cn��ܸ�-�m �����ɤ<WR8{m`�l���zdAv��qYM�]\�l<���+ε���,l�b�<G&æ(iTԪ�[5L۫���۳m-Rv� �Lӝ&�t���Tcn	N�ia{dn��d�D��}���t�g�A�o5�n�����.u�Bite2�*lєM�RX�S���#�3��Bʡ����	�����ny��:㮬�4FbބGX@�������.��6��Fܘ��(A����f�cJ��J��s�n��6��=�۰6{�c�|�E�Yxƀ�O.󕂣6�\���s�ۦ���v���DX�k8LH���<�-�]z���[,��&��]���!K�a���m�����wB\%��A�B[�d&��Z�:�3�gRt����wG#��s��ƫg2�-c�F�I{��c9�4��ث�G�sΝ�|@���^u����K��m����2����Y0��n�RkfHT�JJk�!��t�\��8�K��v�uגn;1�Zp�&68-m9Y�Ĳe��5�b&�=��V�R(�FV�T���$�k.@��nU���v��g	�	��gy�-{u[�s�8�H�I��.+v�u6�qG�i����K[Il�"�3�k�Vn%Ł�f"@�Kp��=�uI`)���X�Jު�ez_N���������!�sۍP����� ���//+�H7d�n�M�uϱ����K��+����m��X+�����G��3��K	v �+��V�m�n��PHL�����%�
�XU�������ºG�/c��E�n"��#����P{��A�� T�l�@�6�����hW�s�Mt쇞<`=]�88cvx&⻖.^���!���6�Nsxm��XK3�c���E�����oo�]�nlY�< \��iY�H%R�{2�a	J=P�pUZڱ�� ��	��v4��[5��2��N':pm���Gg]p���v񍦳#���E���n{z��ħQ�s���=�/K��:^�,/` ���Ҽ7�p�2��_���w�r�f�s���9�`Gb��6"�͸Ԃ�sq M�Uš�S|'}}�=<�ٶW���v�-ҤP�������78���t�ҳSq���&��;W��Ǭ��me�.K�8$p�55�G�D�3�q��M��Pc����n�w�Q\��D��8�.�g����6�
�'!t��3L�> �)8뗮x��K��:�i7:Y�r�lH�+u6j�h[���b!<�l�P���7g\p�����okl��bRC��Y��Mz��A\]��f��ܕ�yb���D�`]'��U�\K(��F���+��`�i�Y�&��;R^��O�/?k�,g*^�f��k��ӫ�c�3��8�<.q��ЯH�fhZl��IcJ`i��Fm ����J�d&bn���͔��۠kH���!����CJv�YjKw%�jU5��"�Yf�%�Tq]cX��6�/$= Mq��`��`�R!bmF=�Uܹv�G5�g+v��NVBn��6퀢,��ہ]f!0Su4�qK33�E��"-�+c����Cf�@r03z�(4���6�L�;�f<.3��<<�<�2m� ��</�)+����f�R����|�x9���Y�/������ҵ�mZ�cf�{s��Q�����s#�	�yH���1�<�8-�KR��Dڼh2i	� �ذ�9�r	��Ľ�uP�脏f�v��xh���I���Mc)�����;���vs�N����U�"q�'y�2��3�.糥�:�p�a�3۬�z<��l�\��|�v�g��y����]�P)5��9nզ�EVۉ����쬌��X.y��M�#��2sW�u��ه����0�u	 ��9kX������j���C;1R�x8(�$��A�x�P"��+�]ՙ�,�q,�v�]�dj�@��eH�GG�jR`C=B�gj��ؘ-̐�1c�(�:�a��}�y�N�H�� ��ں���5��"p�ɍ3�l�&qڒ�Ck�̑��z��\��=3�v�u��k�=�,wd�\JK.��x����%�pƗ@�N��M��WXc�%��;������N07E1	��N�F���-��R�vy��ʹ
q<p�q��ɒ�>�㼾Y��Iic�ٻ2݃�Ӊl�^\Y�5�g�Cu�nӸG(\E�pp�ob�+�1^�l�����P�.��G]�WR�%�n��%�bJ�7P�`>#۩�K��F����� p�<uϰ�ݳ�*�=6�6jc-&Ư0�2�Eg�@�g��&�<c��js��)ە�������˭J/Uϛ�A��k�%�0]�n��A�.�ͭ�A`),p�.U�7�GQ���r�.��[ ���k�t8l�T6�Z�Xڢ��rM73�E�an|�rkb�Vp�E���@z�e�#)�;ih���qj�#H�f*�=���d��bn֝���\f7�j ch`^r��B6z
��xl�.#qَ�;r�<Gje��6v�w&+���&��9ݭ��72��qWR�ja����Z�bL���Ch������q�m��!Ĥl����#ɇ=FŽ��oV�i�.��.f�,8����gFy��\���M�,��'R��1�a`��#�X�?����7��F���N�͖���ά]�pj�=�rp�jxS���+�Y�������+�f�4�,��oz���hCb��u��vG��9�ڝι�]��ف�x��i�qѸ���
K4i�t�����S�VQR�ԙ�����@��f���Ps l�d�KIve�5m�e��M��V-Lmt�(nM�n.i��)�n݀�š5��/'dلvK�FZI� a�V�M̳K�6�cۧ��wV%�)���05�1�� ��]�=�FYa�ҧa����J��J���[/]ôK(:0��.mFC98KI�mt[��z�<A[�o2Ÿ�srNbwXn�Sq�;p��8K�7\��\� �ݹ�u�O[��m`ׇ��g)ێi
YER٨q��k���\{.7��;q�]�fw<�Լ@�t�ń�"�IJ�\��-��Jz�����	��j�X�3C)y��I凅��|�������i�s�w#�xM rܼ��6�rcn0M�{S�Ůdz�2�1q7Fz�w���ۑr�q<��b�X��D �R����)�(�u�a��vg�ĺ��m��j�*�9s��f�7��#\[�|��>^ق��1����� �ۣd����ܽ�m�{J����# 5�e�z�^;6m��������J�h�K&c�h��o�av�7'�ab� 6_e�{#�v�;mpkx�[�t�.�4厕���.1Ƽv�N�ɶ�Al=�x5Lsd�&�5����Rk���5�J��&���p�f�M۟C�����0y*�x�>�[����k�k��M�R8�h׫����rrZ��y���\�kd�+L��yc���Khx`��� ��pQ�>:w��&�R"J�����ll���ht;�ƶZu�.*'��rk�%�.�c�s��^�Ɩ� �Jbip��SK�i+,���N8�Mp�D��� 1���v��ȍ����et�'nkh�7wh��Mc��"4���!V�e5�u��:�Mb�㾾���XunM8�tIYf,��e���	`�t�8��ԴƆ1,p,˭��e������,��8�y�:���s�Ճ�mpX@#V�QƃԘ��5�h��R]��Bf-E�6��#%���ĸw�]��e�4Vd��ZF�����ڲi�v���nb�sn�4v [B����WX6����]�;*6-w&#f��1��@�������M�biˉ��Ѷ�w���!�ʺg�6X\��ֽ�B�c�az[��-�p�\�[iZG �dG�
����&bU+5���1���1�ħ��w3J��W]&�\e�t��Ƒ�3h��B�1���%��Tm�Gf�S)S�Ck�]icm�jL�l Z�q��`�3p�n�m�[�ke�Շ�#�ʹ��[�B4��z�e!�&c����ޜ�9���lѲB�4bS��ʵ��ڏ���A0��.�e0�J �qݍԧ�N�w���%��Z;��1�ϭ����5���4!+	M��i]Rf�mp%·�)�[c�J¡�&������1���v��Ո�YD�9�c!e�ֵ�X��]�;y���n7,p�KkI.�pŕe6|�珂L�q�9��"P�Y��3m+qMi���;��<�����R��פ�$���	��Ӻww���$���gN������o^�ڪ�M���Y��*�Em f6��M+iM!Mh�8��mkm҇(!�%۶�2�Eź�光Le����u��mְ�V���J���3�)l���������X��l��6�ɢ�ԃv6	�7Q�Vx黦��#u�s����K-pS7cYd��ٹ!+`������l�ʞ�\�wX,Lv�;��g�&���v�\��R[Iulݹ�V�Nɰ ;K5ńFZ:Y� �\V�GJ����ִ��:f�9�z������sщrn(��ͬ[�p�{dVS�ۛ�#�����s�{n�$��� �\�6��̉�k��} �&Kn�<dh�	��L��h2�(M�sa����썔e�.t�`b�9{��p</c�KN8JC��T:�N���*�u�����s�Q��C�gq5ن	Yn؄���f��W�D�M�e��¶��5�8r���]+�E%+�	���bfX52ɷ]�7n����6 �Y���:�Ӥ��ݻ^"շ��06�K�� gDm۷�oVf��VJM+�3�w 7jMb��
SXE��I��	��]��Z嫛;� m�1>���E�5s��t��#�mx�FC���gl��b�����&uŤ�W ��c`���6 �y��W&�����ڳ�tm�
�v;[��ʦ��tu4��'���Ɲ�P�#�tɢ×cKGL�\].H���.Jb���Jb�5r�6�L`�S���=�mI��g́Gn���T��k�B2ˎ6��dZ���1�sZ���hز�;X�	EZ��m�lPJx9؋D4�&����[1h\=l�-��r\*�:%-csClq/`��qIKo&��P�k���x6�w7�u<�:��m�s�*�Cd��:�v}Յ^m�	u��ZG�o�q�n;�lm9��p��id&V"Gj1����V�k��ݳ�yA�#��q���S�jْ)-F��+ 6����%7LK���ۘ����:���m��dHZ�p�m[�N��ӻ�t���y�9�om�����*�)��t�
[�n�S�2�N�,З�3!lB�&������k�@\R]Sd�*���=�n����g�q���n1������͠ꎃ��YFX7U �EQ��v�Qa�� ����G�e�S��yW�y����u�9�zr��1ݶ�B2#�irl2��]ٛf�:��1���@ie�8Ѷt�h��8�r���g�7/hP�[15����H�@%��� �b��O�b��Q�e�`V*^rwi�أ���ͮ����ɥ$Q(k&�j&dFI8��rv�y�Y�q��yU�u�ބw�������O����n6&BJ�9':�>��s��|�� ��k
'þ��??+�?(2v�Eh~bTtaq��ݓ�L�w�i���?�5x�Ϸ���'�%&��������j&rB���9�|���Mۻ������{6�����}˽�;.:V�|}G��;��v�?[B�&�e�C,(
�k	Ÿ��e;�<Q�<�s�D����kv%W}��wy��2����d��Mh�_iW\[2��'{|��������"	�R����}��m��Sᛤ��P|8S����̹�=�8�8��脵~#4��,9&(Hѹ+}�h䩖�	��Ҏ���v
����XX�
��2g+�!-T���oi��T|g}/�!F&�D�cL�����O���{/�#��SM���y��{���~}�f�-vz=1FT*2Yq�S��so���{��]���^�������&w�q��F��%�����w7���b������r<��;�; q��q�)w���n����}�sI��!���O\񛳣�#�vЇ<�N˓={�.�Y��E*��Ѣ�.�-�np�'��<�R�}�\�J���o\�I��m�eL�G�.#9+��~������$IБ�3���[�>}Vc�K�q�lb��	�}���)�^��2�. w:�8	�|��C���U���D_��/�P�k�$W�w����0{\�:�*�S9�	�w��al�0��u-�����"hdf9ܝ-�c��dRn'�.��;u�v��("7�'{{����a��ԁ&G�e�/��}���ݪ�X��.�=ݴ�a5�C�}<8#EJ�$X�3<�������������v��-�lN4���y9˹&8wy���$$���D��0�(�A/J�M�8�/i��>��C�}ǳ8���-������0��� Ïo'NO����K�B�2\�9�ݾ��-������8�fW)���z�L�p�$�����g�,��X"�#���񏇽�-t��ZW�=���Ε�Xf��fY5��`cfDd�f胯�gs<,�w}���O* �Z}�;ȗ�%>�\�s��_| � 9�xI��ߦ,{��fO%^�0r�*י����lP�o��.K�My�x}R�ޣ�At��y�������k�9�	}Gw��n������\Z��(�7;'uٹ�uąn�Q��T���E���A�܇�s���c�ÔgϋЋ�O_�u���3I�ӆ�A��o� ��.��I����i�15��!,�)�	u�z�׮�ٵ������mh.���8��A�l�E<#6�������!�6y�����aؙ�}�m_b���-@\�f�[M_z��f�V�y�+�<2[͸��SqWUv�x�lB��Z�܀��F�Y�=�G� �<A:�־���m������>7x}�~��dE��/��>���{�s�I1M������3�x��Gޞ��n_��$��D= Y��=��?��k��³�p_�����D�1�O�Rgy���j����r��&|��^�ѻ���~��� ��W���ym��i�S�x/�����)�ۂ��(e�=}m��\����}�ү��(����}|�sC�4sT'c�(,��{��10�^3�e1���rl��K�9޶��s�7W1���6����	\�e�,�.������pn{u<(��4*����/Y7l�,�k2=�Ξ�j,�lCv��\��\�m�]��� d0n�[eA�Fl�p󞛝��7n�7]�rNk����{f2s������0��i[s�HN�m���)��M�"���;ayN.p�nlK�qhrCV8�;8��s��J���A�F:
��YN#���ݣ�	j�[�`""�eÂ�W������������m�J��~��x��Hϼ%ƾ>wU7n����C��O�i��{I"|��g��q̥���W�Vz�8��������!��k}%��\�F�@`��S�7#�g��.z�'.���x��bOtY�ڎb"/u;���>8/�g/s���"��$l6�R9����r��Nv\��.�;�YT�E/�#)��¼�*�ӳv6o�O����;�Å��? �N.ܯε�v��N߼���O�z����R|�{�r�B{�_^�B�V�-N,)����^]9�#��X|��]���j;�76\�gn�8��+�p��G�>_|�BBbC���S�ObY�ы�n>�r��޾�����M9
C9��n�2Os��K~HD���I��-�E�8]�nb��s����G����!�Z�����碕�\c�G���}�:���I+�zXo���������M�y�5���c��'�����U����(	Q��q�uB}K�b�Z־?|aO�x������fu��ey.>�e��vb�������i �L�^k.�������{���I��rn��+W�D�C"��yZ�dA���۠���	�aS����V��n9?O�Q��杻ػ$Ck�.��,w��\��H�!�%h��I[�rS	����Iu%�G�x��r�,;��j�C�	"B�R+ئ�v��rǲ����8��G��0�@n���+�z�Y�{�s���̇Y~B�M�䉹&͓Eˇ9����*���mNm�䲎�{v�rH̬�����l^�P`��0û��R!g�ui��{nZ��\/���xlc	�fÝe�6�G�ڃ���K�Jü\al��	������ʔ��'n��?��s�â��=&9ِE7�|�pD����%$Qq��BTQ�C>��b��vdqR۶r�36E�$DSp�A��j.!��p!!eE99�v�}s���d+�y|w�Ӿ��;U�1Z���8̜>���\���/X�&d" �)T�A�XqY����]ɗ
𧠛�t��됱�E$�N6b2A9y'^�<�k�q)��.��5f���?͵JS��i�J�b$�/u>_����o�`��0���
����*;tNVL��x�.��s��z����h1�FH�Ga&��>�l����,l-r�2'�r�*���#c�����D��$$�wN8rj��D�o�A�{f�?_)��U�s�����n�W�� }�� �"}�q�\�^<�zi�5��L�[�H�.���� �9�7�6�-�9$-5n�AVQ�b`UV�Fmew���������h�D3������-��D��FdTN�x�X&�bn����_*�����`3T�E�HS�-@n���
�9��u��n��%�j�W�2�V�YM�NT���7�N�˃���}�c��^���Of�9��< �����<\��w�l!I$�R��T�w<>=rӿ�����Z��k�r�Ϲ�.A�0';KO�?b\�(��4��r��F�+���o�&���y<�۳z��f�v�!@��"!l�
� �{N��w��d]8�x:�M�ڮT�W~Ȝ�Nm�\Gf.Մ;�HM���8��󓯹g��s��P2zu�Ɉ,�{a�k'ׯ����ɖ��y��:����N�v<AnɈ~<3�4>�C�;��Ѩ�jnzvq��Cw�z�ٹ�$����̓�s�W5�Wyֺ[�n2J�u�:�A��5���o#���Ϸ
��B�u83�el,FÃKt��Ƶ�cV]Rꑉ2�6ma��5�!\n݉�uH(:�Q�U	�Τ�����]ͻD���`VTEdc��sn�ڼa�ѹ����)C���¶4�ɣ{@����a�m�	3�nv�>��"M�˵\q�n�Wnzim&lбUX��XiB�IH-k�4#%ƯMqmxԫD��&���E�e�@���-�F����ǘX4G-V�'��]~�G�b�l��g}���^���M��r�Λ�^2=��O����"�2��Hc�vl{�!�MG
�����7�C���=cy
��3���c4�.s�����Sj)	Nٖj���{�h���(�e�S���\�<���zl;r�
���;Ov��8sA;��c�ߏD�R�����}�6"5<t��'ׯ��WI���8[���1H��\�ɞ�ok��s+�绿��ߎ��%��l�X�G��p�}5ܾ������n�(�`��ZR3�`�R���Vd���5#�݀UUl�G� p5Yn&[����'�i�>��C��>���z��p���xˮ酼.o9�$�L5��Yy˵�Dz���/r�E�zl�m}�t|��i���p6�76����%�^:v^��=r�`����q�v\�"iyއzn���MZ��Js	x��r&��ڋKY�|�s�{������0��8c�q���BR&�������_�&���ܪ۔��{������sM��ݽ��<�&Pn'#���8�ۜ��?7����W	Jy�êN� ��)%k�i�RY�x��f��4v��8�=�s�C9���~�M�"}�ؗKvo�]֘J��3�{w{(_"H�#�U���\�۩RZP�5Ȏ���a�"cA��ҍ5 :�8&9E�_��ש��+P�������V4y�#.�Y��f�� [}e�3�q��v���0��ˤT��}+G���D�^���G{ݕ�Z��[�'��8�tSHRn�s��<���Q9��n��0FFNkpC�4d�X�D��d�'���59���1�n3���y���ӹ3��=�s��,���&�{�;������8a����s��o���s����"�+Z�}��H��O58zmܾ#Ԛ_D�.�f�;I�'��ׅ{�Q��<�_�zꤧ�ط�
ӥs,��AسF�oxᏤ�g]�|+r�A�l.ְ��<R�g����#����#��Qn,�vn3K���]�q	a�������z���;{ܑ,]^G&-����CT�Q��b��5E�����:���hK��\����	�׀�{wG�H��9�����v�5H���Y{7�S74�C6K�������m<5�t�X�̈́9;cL\���RnSȹ�׶<^i��\]
Y��5��Dwr��(t!��<����ۑ#KaЭ**.�-�NR+s.8#�k��i�v�;Wq�o��������;ͻD�t]M�rkM;������:o���_k��[�:|�,���쏷
��K�=NMn�$_kQq�OS5i���e�q��FSq�*�.�hѕM3�	 ��
�ʵ4.0cz���A�� ԌU9t�Ǔ�Mo۽���u\�g\		�+28�����睊x�:}:�����q��}�������v�V�=m�y�9��ٸ*^����ީkE��?z`�82�\E�<w�5QGkS�[�9��jn�>����;���=䡝���5���Odm�������ۻ:���r��cN���	����́�
�����
��I��ϩ�� v������9�L�~��hD�+����浞Ƿ/������-÷���G{w�'�8�U���N��������J�ރ���5���B�p��8A�s&���V�3��9�R���m�vuZ� �Xc�&��Y+5I���h��B9��ymv��|�������E�!�����Osu��%��w�Nr�&&l�?�9�'��C��˺OB`(;w��Ĳɜ���-�y��ao-;3��"M�w��[$�)��2C�滾��&^I׶�H�	�Y�ڌw��>��y8���g�߮q�2�
�~~�����a-��[�������_�O���Y� R+��	H���q0򯯻ڰ`ǳ�`�`Z����	#H/���Ix`��!�Sp<v幊�� �7YVv�Uj|{�rUJ���b�wss�$�g��12L7tp�� v�h'a��|�筞����Kwj�n/�o��/���e]4���>-���ep�^&�瘺R��U����;:��MX�  Z�v���,:�h0�6��f�p��;~��|{�&qؗ�ӈ��O6�}�h9 �����\��χ0@[JB�f=Փ��=��9Ύ�Y��l��mn���c�:�~�"ob�>D��y��	���8�*9^�O+w�����?o�y�/�rE��ڎ��qQOf��~=4��'��"N�8<t��IG���[�[�_.Ǳ��q���HaX�|!ء�}Nz��͹|<����c,���R;�>^��pϓcg{�Yc[�����T�_C��!��C׌�N��������d�$�{}F,���cگuf�I�Rs/0���������	�q��W�mhO�=³��Vk�۷|<�k�J�b;��;~)�Ԣm�(�K��v�#���V�mXe1�c²uG^�<u�7)g�r�4��x�����:݊�v���sQZ{�C�q#���ǔ8]	skRU�	��mA��f�����VVc�3���f�.��5��Xր�H���-v�i�-��� ��V=����s��jc�ysn&�̶��k$.�^1�cl��I�ņƗ����&�#]i��@�c,`���%{�d�ɮ %�A;%��Dtp9�iΚ�b%8C�'���}�����x��̽>�m$[�>+��&�d;"iP��������ǽ��A�8�'���(��~�Е#�ͣ����q�kO�@��;�;)M��K龔��thDF���IL�2'm�x�{��}����汋�-�k4u�VWǶ����3��^_n�v��F�A��N8f��K��F)����yp�����O�v�;~J��8C���w����ΛK�&D�aw�����>�I�nj�ϯx��������c����}ә��'�gV-���(�J��J�rP�61IH.�$�M�e�ڒ�����sp���]�n"����'|�z�l9!C�x_yO<o��H���͢T�^=��}�8���\�݄$I�c�i|[���>���2p�RCo]��=�ʻX`�� ��ǝ�i�Yq�����܀�;TC��ͮ�n�D��0l���4u>�����]��M�a�K��I���n�s8��C��]ʹΌ֠l�$�!r.ze���G2s''������6��'�7�=�7^{��`�vu���]2b,�gx�!��T_�_|wLodD|w����asN����ǽ�#wq��y��۝�D���LfE!1���q���N�^Q���Yâ�j�j�����r�y���=&�m�%�MH4�A���[o>9/=���qfln���V��j*�(��D���1�.C�Z�ou�s˻1No?�\���?�>_tj����93S�K���m���#��ˋ6��p̹��ޞ>!�E^�Z?u|+��m���³����L5!��7�Ξ;���qQ��]� �3N�:O#�;�z1�!���w�8^�d#ۭ_�X��̑r�aZ�nSD�v��zp���N��*������<�ֹ�^x;ܝDp����{|��G2��7�i�q|��{����#1|ߗì��v"�s��=�u�tL�B�"�M�^��ޯcﲯ���ϋ���傲�f���.��֦z68��ϻ>�n��e�6���$��C5����WpJ`�sإ�!rm��Y��CvG��w�޾?O>��$��܇�|��us�Sۜ����y�K�x	�<%8�Rr'���Oh˻�+D<)L��y�rrOyg���y�uN>x��d�h/m��F%B���NU��-�c{]הX�Rc�-x$����Nm��,3a��K��!-�L�c��%7=���ه��WB�����|he����EoY��������&=Ֆ���"���q=�{��YFN�#�u�����]d��~xC��H>�~B�Z���H��E��n9��|��{ޞ��p9E0������K؈���]̻��e�q��`_��T5�����ŘE� �u4QP	lӶ���XK
xΚ^y}����۴^wH��*<���b����ϟ)�,Í��!d�d�����FwQvu{�����<������HRB\�3S�,T��ڎE^#{fNNr����Hy�;r����b	�Y<m�@��I$����;�>����^b�����N386��<�l��o�(C�G�x��M�6.�����9���8���*���FY�F�����x����:��6�.�r,c%��o{��Gf����*�"NRx��>�κ�-���p�Ezk�i$� ��Wc��_cGf�ݤh��o���8O`$������Xt�s ��`��]��wo�y�����e���������"!BZi�%����^�)�ղƃd��h�ꨉ��T<����U��e{�986���zʖr�p�5�eH���4�� ,4Ғ�4Z�ɖ[h{N�F㋩V�O*<��76��[�n����Ӹ�קs�	y�9�<9�����G�X�<teK^Ր�U��M��M.���F�n�r�uR�#�3�L1K*��ct�i�"������_&�Rbhy�ef�:WU)����,��ఄlE ��*Y���lZ�jp�~UO�?'eV��}+�22�x.OeK�@��4S�����$��f���v�  �p�x�%�t�V�z�-SK|n5^N79�c l��J݇�ũN�l^O�ANF���㏋���s<��u/|>}���l�/�I��$N�7�[y����~\�~�oI^"�����Ŝz	ql`a�;;��{j6�>���S��u���N�R�OH���b�&29�0H�,A2&�o�mspյ�9.����I�ݻ!˕yٵ4�T�Wuq��y�ǋ�ٌ�G��%�t�E�#�@�7[�0eBǆfـ �9��kg�WU��1�f#��d�		-�|�y~�w���^�}��W����s�G�V+�ud<5��;F1�PM4\n8�Ü�w�2���Gmo��'�J��b��y�l����n��=rgO W���'^l;�9^���$�Ĺz{]B�)^��K}��/����'�N�sȋ.�2����B�c|��;�����K��Rp#8�DQE�7��0�"�!T��oÈQ�w<�흨�¤f9ڭ'�AӐ!B��fH�ió[\a#܏[����gmu�Q�%me���+L�c��u�:�<|��)T�Cm8���ǹ�,��T���̬U�|*��e�>��q��#����Bѳ��f�Mi��P���<y�GD��R��e�3\�dhD�@t�np��Ҳ�a]���&v��PO����������a�G�;�g���t�s~8����=�y�h�]e{��DڂF�1�|_�-˛a��l&Ho�4���Gs��חњb)�nt��U�E�e$�"2'��λ�ˇ$G����]���;�����m�ëo3*/�F�5�[����o$|�����S}���I�H�hḂ���-rfH.�S9X��S������di�����0�6���ΜS����k���1
T�*fn:�bs�Da�3���Ocnͮ}�醜�����'+��o��s���x����'A��m�R$���9�J�
��fN3R2�"�Ӫ:{7����W��E�� �����A�0BM&�1q 5�qe��<��l����X�8�Kk�(F5:H� � Q�S�0����]���7�ہz�8��0w/..�(�eD}1��{Oyɾf��2�a�<@Ɣ��\�U����<b�+�}��A���Ӥ|3�����aڗ��}�( :#�2�J\s!��L紦�������/����4�S�r���@������
"fRS2ky�OD��l���c�����}��v���>2�����;�t�'��k���%�ⴷ�܎�:�.Y��&� !������<}�A�>�w"���W�͍^������"|��;���xމ�������ș�w�a��m�R��.Z�y�z�����v�-�d&i�Re3tj�M��LG(RZ�=��QӀ�rn[m7=��3L�GVUF����>���_G�Y0�r�a��I�|ci� �Z�:y�FN(��x5Q�Dn(c$�'��Y��똁s �Ӝ𾗭l5G]þ�qOT�sf�k�F��__B���yq�zfH#��q��`��5'�^r�N>��8(𛍀��E�NK�{���������7�c-�C�����#�T��}�#�:�˪Ȣ����-)]���S79S�{�8jPL�0&dwoq�4����Ǒ�}�>��xy^K�=s(ogTF�f���u�F��n#���UL[RKZ��l�[��<zL�	�W�����<N\�I�5�Izz���M�Ch���s���'��9Y/X��!+�`Y�B9f�۽�n-�om�;|{ޛwU�z��	�X6XMT�qp��_fూ���jl'����r�����'i+�&k=���^��~ [��zί�h_������r8���c+j�<��Oo8���yl+^{ۅ9�ɪ��^�e�3������vf��؝[�*d�S�x�i�L�M�"9�t�w�	���~��`Z�����޾���=��t�{&��e�Ɏ�\�|]�9�l�/��w����ɇ�����#��o<��G=|�v������l��MK�n�&C�͓���5�{��x�X������_o��	��c��Ǵ-GZ|z�8��/�
X�uk K��i|��侌�;"(:�$��BI;MbI��r㴠������ě��w|X{���yk��޹��mp�{=�]��I���9o��)R��1�p`���w wǼ4ہ\�g��ɇ�5s�L�ak���_>{���Y�?\�̰^B�H��Z���6���&r9̴Fm]7�S��XT���,DNʋp��ŻZ�N��DN�H�!�V5Ʋ({.{<� n�=�<y,�S���ZxKO%4�^�J^�ѫ���n�'S�Zkuh�DuLX�H�v�cfF�͸"i�[���h0���<[����%�yß��=��֘��zݓ��3ѽ��	��[b���j]oU��:�{uW<`���|�c9%�=]���UUu]��Ȁ*C
� S��1h��L$,|�i��u�Ck6�9x��r�*�� !��]��z�n��z�s��^�fɁw6)�F����tF�n��nR�R�\ZƳ<��e�E�a�1f����Vޠ_*]vv�D���3��8-s������4�Ί8՚���2�J^^�qw�t�?x��!�.�3k���P�i�G\=���#���sv��a�Pl����3��c��[[��1��s�)�t��W�nn�`�Lgv+��k��\��T̠:�`�	N*6Y���Wj�b�Mm�-�[ex�x�Yq�8u�P��1�r�.�l�����3K���`��ݺdլ��q��y�s�f�ث/e0e`�{�y�8����V��L'n6�Χ�J�:r=�����ʑZ���mv����C�c����X8���v�<%[�VJ]�
�,�v�!�ˎ���\�C��Y[']����I��9�8vXnI�F�\�'�����hc�M[�(�I��o)Gb������dі3[�q�nG���d�D�M)pֲ�pzҽX��هl��q���fn��2�(�[���X�,�uw(�K�`��R=v�^�[3�ل��[-4��k���F�˻r������v��v�n�`�#f;+-m��e-#R���L��v�#�2�Z�B냜4Ƶ6��;��7t=l�u\Y	�0�SŅĖ㲷Lb�X�#�7:�<Wm�L���J��T��^�m�-,l��<B;�"@n׳���It;��Lcr���]�B���w-�,W+wN�l=jJ67��Л�|N��'Z-�={kGF��jr<̢YX[.k،Do��f��v�
d.��'��G��#��6N�c+���k5��X��󚂼� ,�����RapۮR�b�erǨMr�fe�5"LƑ̀X!Rc3B*�;��u���4r]�v�";b:�H��b����G�M�]5�\�g��Cc[���?z}͞��k�r5k��3�l&��i�k��Ge�7� 3`AيgK�R�x�7,F�x{^�=K� �u�3��Y�hbXð ��5��XS��eV*�f�P�ڄB�\Vk�]N��2P�yb�|��A�����iㅝ����'m�v$�*��۳q��s$�����.W����%�f���i��lͰ�Bf��v��YV �-���;X4��h�qI;!W'�w+�q�:�E1&�vg� ���lt�2�I�1�X���W
�
���I����~�Ca놐��hfM���z�EG�<w/%l�|r^En�b����Y���	Yz���$��}������l�Xe�nY�o;���Ν\��N��}���;*����T�/��}`w�x�um��[�#H��(�pG��}�j�Z�|~�^w>
8ύ�α�E���D�ogD	l�0�HJ"f6�|�<9e����� ���ů�x����n1��g=/��`�-t��i�F�iFMI9��;�<9�Ƕ����q�]%dt�t�"�k+U�Z4���-=��oF��p��|{�8d"�q�.�6�y2���냵H2v�x�g�C�F�ޱ�N�@�RH$G)�$=�pz\�x��u��Z��϶{p��+�_>��>Jy:�/�Sc�����h?���8�9�����;�O�r/5|w��a�'�p�xq�^�����׸y�1���*�%��թ�b���G/l��NM��=YOf�d��E�5ܳ�f9']�ʗ�_?}��޲�j4��=����;�wI�ĂN���-����D������}�;*=���v�͖<�a�.��o����с��0�qrb��3���Οi���o��;���7�.���s.pE'x��㞋�8y�����K��nB�u�����bw"2�۽�>V=>�p�j�Gܾ�B���]R�}QS�����x$�s�
�Ck��l���Sn맣��+KM��/B�遣������p��΅9�oYɹk���������'q�&�[�yT�c�2{'��F��p�#z4�#�����on9�S��S���C�;��w��:jg$r���w�\%���
rl�i��}��зf��d|:(���ozFF���H~�\CX�]i���٥�r�k����zB����!��lA���wVp�;�z\����仃P���>V�$����x��Se�;k�=�ANH�h��28�/��g�t7i_4/0��"��۾�{�����(�-�n�7ۚP婧���A1�1��p�A�Hy7��/�ơ[�;m���_�,��}�w��>�����}��s�����%��l�M�h�)��m4�a&�	���e����j�ن�5 �Ҍz�BQ���؉�6S��j;zs�=6_�s~�W�%M�=�S��c%s6�K��}����q��T�EHS�&ۇ8�:��
�{�J$��ɾ|�=�_|i9�V@�r�g���H��U��Ò"aHP	��&��t�v.��Uu�\+�#.�`3��r��e��Sܕ���Y�$h�����(�f�3 Sw� n�Eu>��ggm��S6 f>o7�5��^}�Y�s�g,�&t(�c�'�!��1\b�F�f��I������Εcs����V�yd�S�����swS�;�������ǢB�>��N�$��G.�k�.���)~����ϝh'_e������/}�S���nɱ-���VDcq!-
�4�%��2`�rY�ՃN��7;λG;�r�L��Q	IR�L��T�N��r�sՉ��B%��8��܍�o{���%�bRT�`w}�7@'�`�<H�D��v��y�#2Pʺ��h=�vo�$����⫬��ε�6N=�*w�����xc!��	��/�|w7���3��^_.�B3�ߎ�t���J�%BY�N����\#m-��L"ǔ
��C��(pN7��ݚ"�֔�;��I��Hn{,�θ����b)�@�<�3�O���4�)�_�
\��'�u�b����a�^_+e�7]3�t�h�}`�Vyܩ�x�ڜ���<��/�T�'�||�m�r�N��ۻWh�1���gt�,v����ƹv6ys^���y�G�x� �3���Kn���0�˞���\;.�1ڬ�+����-�lB6��E.&�d8Cj��n�dT42���e
X[M�e��n� ��|�w�Ɔ=��Ѻ+uQ�rvDW��l�nv���ck"#7M\�˞x��m-�]���l��n���8��oB�����2�16˳q�.�ֲ����Z�oP=/F���o6��f�Dl \hY�]ZnD�r�'We�WZt����&kHƳx����8im��% *7)�"M����ﱯ��2��me�{����/��=�YHg#�e���m���0�w� l1Q�ّNy���?�Ϛ������ߕE�P�s]�.VӸ�/6�
&HYm�#rw�F\F&�r&�o^�U�Ş9�l,����P�S��3�C�p
���d�w~\���<��rT��đ��nLᇚ�{x]�|&b"n�5'$�l��a�O��w��Ȉ�>&��C�~cwF��;��qx��!���]w�Bx�%��/}iLP���(���f���v��ox������RQ���0�A$�^-�n7���v�RtPq�n%D�ݳ�/<m��F��&&[�z&�~��6-�B߶{/^��]]���Y��@�tr�z<��x����]yC-(�1��Y�9�f��ӱˎ)�Q_e��.ƪ���7b����_
���g�N�����Oآ��nÛgy����{��$���$daS��An�=��gr;:�h��]�t�m.&��_�r��A��J��9O t@Q#!9$�6ۇ6����xw�\��	�W���
ʌ���;��Tm��d����uf���{��&�,4�$'{"��Ϲ��<�l</�Ǻ<,8v�&������y��Ω���m����K�����;����Z�����,�@WDm̱��h}yj��������kP�9��Z>C�>O�d�l���q>�lAW6�N:m668K�;vJ�a]��5��=$�F�g]�Jkkj�͂_�;�sqgx��v[����G�qcc�5H�-�qZ�=�f�ٻevH��A�1
����Y�睋v�B8=@�;OMQ(���x�랊����7��=Z ��gu��r��
L̔I���Z�Z;\VB��\�ۂ&���Q�VRQN�����ɧ�� Ɛ��T�x��I��y��b�ۻ�7����60J�H�|".o2�9�9�}6n��?��ת�5��x��bؽ�?*�=�r�|Q��m��<[�u{�߯�����#����f)����5��
��1�|ٰW
>Da�J�N��k�-6X~a*�)n,�zn���ܮ^��5��H
�%-=���g�r�˨YJ���7��7��3�^�w��l��$m����3.<�/\��N:�%7%�b�X�v�\i	.(�E��L8qw�{����o1����>[�z��ݗgA���"P��ΒF}�ݟf��F�i �B�����N�I
�j�Gw�.!��Gku�o-�{��1��ouگ�o�K5tX��!��!���3\1z������1�?���_�7�;�T؞���r�+O%_w��"L�I7"n'�-���*&gA��V���x%aלp�u}]����Fm+���DNX��ݺ����ͫ��>�����%�y�;P��9�~�i�P��֥�.�v�F9=��*�����6�'}��ֱ.���u�,��<�����4�97{�BOv�*!a����mŧ6�����p�����T�Ǽ&v;��<��~ﱎagV�u���+�6�ܧ\qg�۩n��k��Bfca�Kv����#4\%	־�̏����i[��r�ߘ���|t��8'=}v��AΈ��6��IFT�Eqg�0Gs��g{��".=������j&8�/���F!�����m���޾y�'�@ѐ��	��y�uWd���E�Ͼ0'?�ۣa�e��.ʌhV��X��z���@�t�
q7i�/-�vOM�Yq��x����t���y��r��Q�(��9�VqҶ�y��q���þ�'�C8�e�0�H��x�?��~�|����뎚c�.S4zߵno��'��}�웗�|DwC���ו����\c$؃	�����ރ��=�?C�=wۖ������`dg.�f\��ҭ��ү� �SEC;3���=���s�$ܑ��$�D�v8�E�%,�)�x�5wɶ]�l�u�X.�\�,�3ͣMsc#��e�\Y�����F;/`,q�i����[�ǅ�m˅��`�x'���8ޟ8wc������h�NRz���r���p&�sņ�
W6E��H�v�0��6�g^ݠ�)+iH���Is�ὶ��tŕ�H�w-�F���b�{mF(�ڶ��{�ހ���+�q���n<]�����;�g����+����En-���hA�Z����o��w�?�?��r��}��~3��-f��}, }�Zda�Kt�Y�s��-@���t#��;Oi員������3�T<\��ӣp�"%��+|���w�~��lѢ�7�r�]p�GI�&1��r_�F���ūqP��!��Q��������:g��'��|�L
�_�
!�q ���ױ�%������g15,�_�Q���L94���L��_���}��0�M~aׄm	DXI��T�����bB�ﱷ�)5�w���̍ۅݪ�،ڜ��u̚TC`*��c�j�]+j)���]e��9�Tqٜnlp/L	���&����5���=���p0�]t��2��o+���݈��[U����=G�7Z�8�y4�r�#�p�����g�����H�)�7��y=�ztmI�x�}.���l/:<�7'��x)�<��擅�����.�����W I��X04#{���w�q�g[C
���}�7�n���S=�cװ�=�P���8�2L����[��y�9�/���+[�����M[��"��f=�����ێE���c2ؒ&ی����6�?wy���)�Y?{�bD�����z?��Xc�yv��b����{�.F�nI! �)������_W:d�����;�حWnщ�԰�ft���`��Ț<�z���E�Z���^r魗#�v�9ڐ�����y=��OAb��Y�ۭh.Z�lP�-�c�w�ʰL��o+�l�����)��}R�S���?t؛ӂE�܁��)"�i�����W7���W���Z,���ǽ��mF��wN�{�(��A�
s�J����m�O��ȳｏTFI����'1��wǏp23��9�峗�F�����tZȪ�Mc_�G ;��'7��Yyf��< ˽�B�R������{�ܜf���߼������2����[l4�i��3:�}8���o��v�])�u���iQ�1�®\��o�no�Y���As8�t`(q�L�S�m�F���WB��\��e%���N=����q����]-�+�6�o�ʹR�2��L��3�η㼵XfN_�4rb۸���X�6b�P�B�#ɘ�{Ǎ��+��<��e�wx�7�n���a�l�޹s�$�tlf�ݣ��h�y<�Z4���}_��J<��o>�~��*uxˏ�*�������	�kCs
�l`A
��wcQg���kx�rL�	vM�=,����"��(Q�/{aY����0��f��m|J~n��;V�P����ݼGg�~���>�.׆�<W�Ģ�/9C��W��-�ȯn�Yt������v�J�gc�&����� ���5pرdl���������Fdf�bU� k�fg��r�c�2���ʰ�P��KodX�m�7x�q&*�²M39����8�ܽ�^}����:n/c0Mk� �7A�n�]�0�n�JM�aނ��.��jުu9C�����sn��ۭ�5����CB3�gd��nOt�T�[������m��*ʽl.z-k+y�+:=����Um�7pn���"'u�^dKcb7Jțį/~�h��]77�ݞ��{v@�'���5���#zI;G���px���Lh�j+����K�������vNsrS0�~�|W���w3�}CP�����O͡!���e�9��οtep���{S
�/������z��b�?�T�Da�YQnclw�W�H2_#h�0�QI��ۆ�ݱ�i?zs�r�Lv�+��]�r^�����W����{���oe�z������e ����7B�v��Õ�npX3=���6<չ)rư�jLR�ɐ��I�b�Z��!{�������z���ު/%>���w�n+=��J����"<�09�H�k�Ç�n�g�{6j�����~�x�J����~qo���V�n��w�&A���a����=�ǰv�����e��a���|5���>X��u�}��H�S�O��t��E�ّ�̳�<��J#�����_m7O.x�b��2�>5�����4u���rEiUR#)(�1��:g,#f{��OWy{!�"�oo�-�"�	M��r��D��˿�̕)l\	�"�,��tZ����!ӹ�[�I�,>Dq�c
CmI��c/��	:]3������F�V��.��5��93��o�a����AJf�B��՚k0���^^h�mHf�����q��.޼����Rq�E��|��g���<�ْm�1\v2hd^��zH��rE�ӷ5Z��W5���^_J���$P��ؕ?L����A}���%@�~ay@�.Ȯ�n��97�r܈�[k8*�cz��hBP�
�`�"U�̳����9ٟ��T0�!��V�u��nf����zKp�˿c>�$���1����gkJ�N_(g�b�{��;��5=�������|����k�O��$U��6YS�a�0��lE�����{''k�,�����o&�?D���\�,�Uc?�
��.k/ԇwWsߙ��"3�D�GF�W���m��c�S�[��$M�k��r�j���ggc��i�&��x{�p����Ś��}��>]���9\�Hk�ٜ�MamT�H靊��k�0��,9�S5�/���=R[</R�fv��l\�.�f�Z$�Jd֞�W����`��k�9�������ٗ�i�:�ͨ��B0���lXoʉ=�G��=�t	�W�lP�nv��#M���u�$dԽ^���Me����׳lF����:׀�x��^ۗlFq�Bd����rd.��p���@�>��CG��դ�c����Kw&�a
JA�f� h���J�
+S���w�޼�Y���t��!����6��B�%��A����9��^���q�"*(c�wq,�w�0���ɝ�Kʽ�!{�}2{t���ln��s�"xE=�44��囈�qSe'#�Op��1j���W=��Xf/8��
B}�C��s=Rj����l���CA��p� ��֚���c��G�4��z��-|�uE��9���Ur0H�S.ɥ������I�A2$[i7's������j>D�9���y�«w��[�6���o�|�9���xO�H�M��nM�̈́sY6��(�nJ��]�Ӝc���7��b	[�\@��"\��|�<��k�D/���u�A}��UU���ǽ��uZ�s��76e؝��P)�Lm(��8��U�_@�A�Gkݹ-OͺN/?=�w$��3��$���c�1j����ˍ���
��۲PD���}�%�%o.y���uj'Ǫ�y���E������hA��O>�1��=�1`�Q����OxM˜���/���2W�a����
����ќ�]ш许���ZE��|�HS)vp�p��o�rߤk���.?�E���d��qh�
�ȅ&�NK]:��U��6��H6�q��rs��E�_���wUüͬ?=S�7ed���ŬcV��_�����qw|�F!	�"�RD�=As;���P�3ӌ;��� w�ϡ���	��E�"2@�*Hw�.��s�"Ҿ��U�^z���j��[�~�6''�M﹇� ��Amqs	�S���KI�tpb'�D��o+��Md�wVq�?Iԧ{��z����`�����"	-��q2d�`���f��4��n}�(L4/��.�s̀G޲v�;	1`��w�j`�Xd��ɠ����N2�(��2��E�{|��3�珣����v�1x��v�{�M���4-"�{��Ǳ�{�q�Me��R�����3�/�9�`���^i윜��in�B����3����AS���ϊ �7�}�H�
�i���1f�����t��������O/�rj��I�u�i���c����{�dR3LC"��Wq��l-YG@�/�FShs-���Ī�<i�y�JT1�c`�"HH.��te���ۜ�	�z~��\^�δ����/=���3�5%�g�����@���4�Q�H��ד�2k&gK�.�븥�$�O"xN����������5s@:�"J
	�nMs�d�{��{��|�����^Wi��Q�*�oغ�?��|�P�,������NB�9��㓺TEMF2�;	no)U7};�q�tf�{6�e�uŞ5�UFU�b2*dzII'NVn��T���t7�A���L��-q�3Q�ј�c!��V���v��p�����1>�=�ʾ��(>BQ0	fD�<��l�^wÏWɢR{���'�l�<���N)}=����j�d�`'�.��E�"*,e6�b��Qd���Syz��k��ȃ�ղ��v��(�ہ�K�0�I7%�w���v�s��9'���6s����p�׸�/t\A�����7��lG�4SM8��o]ۛ㊑�t`JVSp���6NNA����˛Z��D�7��dĈ�!A<$��,b0��i����N�^%;��D��N�Oe@�S�s�g��Ռw�W.#j"��	�����}�:������3��NO���˗Gfa�Ƣz3qT��Sg���b"f��1�ok�_-��
���v�@��<y�Z�5η�ns�~�����lN��t��bS_f�![R���i)+�l�ޒ��'{SI��v��ޭ�x��b8�x9\l; ��p^��"vy��ݞo�)a�0"��6w@ۋ'E�M���]nq[s.V�MM��3�n�ġã�rG]q����s[�=qӢ$�\��h�[u��l�/����Dq�mF��ma�}s�aԋ�5c�Д�%jcl��;hL�P�4pl`��n�铇V�PK���I��#Yl�2k��ԅ�.�81�v`����i��ӨLse��J�	6�-A��2l!�h�8��F[�.A3��T�&z����A�MֲT��,�+�"�L�����{�3'�;]=�u2]���>�;ݕ��osgj����:l���[M�#����8�����g��x��ٸݜ�Ѵ���M	�́���G�]��"�6dw��a d fL��1��z���؋�����&u�_N�ju�����;�����Z��+�A;@�\e�ܛ�vΉ�-����=�yg&��޿k�Es�{��l}����ژk,\�k�[���QPb"~�0Q%a�^���8�L!q�|��s�K��{��Hg��W.�����a��_��q����� ��79�X�2�][�s�3Z�����)�YnطEl�n�` �G�L?.^��E~���}zU�L|�(��p�gfV��4�lF��EBmD�lB������{��pa�0_�,�3�@�n�-��fcc%E)v�n�y�;<�����ï�j�|;�c��F\6\3��fޠ !7w��@y�l�����P��C�H��_&W����u�3y�aB4䅸$�]�]7�;w9�fG-ٞ�aۡ
��3}}��_�r����n���"�5%)�''+�$N�0z^-�����y��۫���V(�~��銫�Y�m�P`�Q	��e���zծ��,.�l�y�o�Z���'�^?]翾������iy��������"k6A7��B�n�������x5��a�.`�u�uHlH1*aD�jF82{�N�ɬx�������j��`��$��mņ�εcvci&y�c�<O��M������ۿc�O:���&��8B�}㳝��&�.����M��q�P��L��bM��ؼ2v�Q�]x�"�eTѫufD��bxTR`��:�5MCQ�C�VpV$a�2EC�{�ε��RΖ�^��N��gI�,*D����@ʜ��4�'�1=ӬV'V'|V"T1`jF\R.rr��6����Gr��*��&�p�ц,lU7];��]�:��s�_y����M�!�Hc�c_}���<�Y����|~Q���g�?����W�I"Ȼ�3�>j�:~��miiشԋ2�[m!�bGo1���+��rv��.3�<(�0�G{F p����P�3�>�}���B����'�(~�.w�k��p�:�����)�4ԎM������v�d� �|"�l�Q�z}��>�2��m?�NL[4<z�2�M��IㇸN�a���9��}[?��y���nb҇�p`�MN/� ģ������ԡb8ce��[&�����=��=�S��̓O����x��P��]�9E�8������5����f���;������������_���e���{;�����\��h��*UN���1�_
��2��j8SI8�x��}�\��U�_$�vH�ό"�֡��&��o��&sB��v��ۗ
To�
+4�1U�'iAJ�Bs���L����-��C7�֫�*4��#V�/�ߖ??z��L��꾥�,:6���姅S�l뭙3�s,����Ǜ�B،�n-�xj��>M|�y|�Җ��?�M�����K��y���ش���6�z�������d�!Mž㛁�f��C�׍پ��˨�,���蹵���p>yr���8���2cR0�9��	��0�70���u��kV }�L�U����LJ������|﫼�˞�ӥ�$E�L�m�w7�ɲ;��0�T��t�������'+D����$ȿ������M��ǧ�p�ѷ��iͰHĮ�'mM꛱�E.�j���݆L�a��{�O^9�ͦ��p���zu�l�w��^Q���!�q��s�Ɨ�t�=�ݞ��"Zlf�C�嶍�]y�;ѥ�7e�����o:�嬵1���^�t
�β�NiwA�����iU�DLx.�#�}� '��h���a������SÉf�}�$��x���rtkv�;
Z��_b�/y���Z�Cr�ƛ�o��n����^�^�� u� �{����y!E�ý ���r.���/��;�;F��x%<}(E̻��9�Q}H���6b�]v�7�ܲ����?��<-�����znf�^�����䕮���8v!}-�L�/!@��TTU��:Z��!d���]L���0��8ga�f�)�C�.&7H:���7�/��OJ�+ �	Z��N�,8�ueHp�Li�}�I� 9�ga���Sǝ�p�0�޴�<{����y��N�z���y��6{O���t����Ry�RR����٧I�������`?���,B?�j�f�1yf�n�m�1��f��܈�o��"��3GW;q���Ńb���!��z��L�7j4����[
�j����E��sG8��G{zK9�]h�8�c���h>�}���ȳ͹�W�,%��촎�ộ��,J-B��¬�m�F��L�Xg�_>��C��\�Z����wn�i�Z�o��f�-Q,�.h�y���Yޔvwx�I$�Oq�e �m��V�S ZF7F��\�{��Ѭ���\�[���L����b�t�[ZYk5��Ԁ<���6��㷨��y����g�h<p���^a,�u�f`�H:)SLY[�p�h�oZK,��
�R�F���D�;l���C��L��㠖��{�Xj/.��9ixmn9�m�H<i7w����n���+�p��u�uƹ�!�'�7��k䝳����O���8��O^R�v�f��x��#v'��e9˜ðMetZu@������״����-��&�"�V�W*<�;X���C�Uu�m�N�vpt\�^AS�tX˳̸��5�X��<��z�=�q�G�H�H�`�:��C%n�n�ܼ�v���tpiycp�88����n83�9���3���:Q/넄n���N�lN��|8��ܒ���=nwHsȷ4N3ٻ	6��3��1����.-���w/7`SK�� 쮅+F�{t�lG1�w��[u۰�<"����m�*�%���;��F*�OC�[uϱ#uUר��(Wn�v瑲�-�h��+�tA�X�*`a�g,�2��kΓ�����0�M�	�L`�\=�;v���f��L5��M�Nͻ9�k�:�z'
i����FiYv��5�-e�)G�%()1(�m��u�S��s2�J�u.��0�4�<ƬCL������C�63�;���+��i�̣6H<Q�Hj^cۇ���Np�yd��+I���mrGAz�ˬ��LI�Φ@�-N*	Ml6f�Miuٙ�F��n��!��M&��!��-�t���jk�CcD���%�[�:�c&m����),���i �A0�څ�`����b#<s�!!�L���@<�6:���Lj�1ǭ�Ϯ1���-sʶܝ�v���.ງŦ4���R�M�(�6x��0&��%�Xb��kX�p=:w6=��8�/Ti�s��Ñ. 4ᒰX⎍��э6(���J��G(L�܎�-me��T5��AD�vHD�ZX�@�p�q�J�nݞq�V��V��V-ae�@�0������r���j��X��X�[L�Z;���Ƒ���<ɠ��j�=�'Fҭ��r��(i�0�eI����c�����$mU����J����^���]�vT�a��^�,`�lf��r%�P��8�V[#2Ɍ�a�-�Ejm�۰�\$����9���:˒@ҀE��6��+���4��D1�i��DF�p4�׽���..,��t~��(�]�"�����Ў6��W�Gr�����i~�MY������	M���B�|#�D��q��5����QĐޓ�B�wU顇�5��"��鯙d�ԍ����p���$�=׈����!r2�I@�	8�x郇�΁Dd���Ml��ƾ�=�^U�4(�C. �22���>�ۊՈi���_�C&��B1�2�����h,iI!r�`�%���z���^�h<B�75��4B8Á���
��U
k�#DZ3 �{�4�F!�S�@�}S�m{��re�5cx�"�z}�.�ؑ�2��ei�k����wW���cőd^���`�P���Oˮ���(�f<�_�����dt+"=w�X���~<5_�=<؁�ɣ��x`t��$��\�K ��m����n#�WsnA�����5�P���D[�z��l�_`;5=��Y~�(���M#M�ag�6vߕ�z�⌟����(����/�l�#����~O� Jp��PL��ӆ���Y�Ezhiw�y�@��C�����«��O�Y�7$��_΂�e�ɪC��L��-0��2�fy{�i�Nj�-�T�p��"F��&�"=+�1��5b�"�Ȣ�^�43W�hs_a�^�߱�U���ĐC�����K�ސ�믑i�i��3�a�4�dO{/��,Εf���t�ON*�G��Æ%)�8?l��7�&��#Ԥ,����k�Rt��ȳ����ӫ��9#p&ˑet�kz/�x�#$/,lݍ6B�dqә��Y닲3����6l�u�E�aF�M\ᔳ툙;D/eb��ȣ��Q�����2F�p6qXӤ��H��J!<�����G���g
��Y%V=ysv^�"�▾��oʇ�j~dE����Xg���S��|�2n>Qc�hYa(�m�f�Mŵc�h��l�lX���'Zآ��J+��q�2*�>�C���-��&4$�ފ��!������6��F�!��*&/ӻpIG��Q�B��6k����Z��8~A�b  e�R��4�6GI#���W�[!�#V�0�9�B3�?O��hh:D#Hf�w��v8N��ƠH�U3���tm�G?Q�ȋ~�7E�ĐL�$�Mŕ���|4�C>\���:xGZ��)���}�В.}9��W.��]����=?E�x�>�F]��w`���S��������
c�Z >��^��A�aփV�l��>'���O�hq�d3����Xåb���f_�h�da�"�6�iH3�8l�?X=*�{nC��92��V���<#�~�XŃepɑ�0k{"h����x�0C!	�d����;le�H��ߠ2-.�:u��31�E$2�C>#�!�u�|���<���>�(�C�H>���U�$h<Ed!�~�'W�-��=�M��?3���י�гł���T�[�Xs���n�U�P��L�b[��Ҥ(E.��4+C�0�f��g���ճ� ���7��&��P�DugyPM}G��'$,��{H�4V�g�#3�(��y9��F��dG��ϭ��Q$�q��"He�0�����Pf�|���n��Qx��r}�.��5�!����cu}di6B�Vxݐu����y�fH��oA�P�E�bB�v4՝:_P�����e�":���k�d�8��0k�:�T/_Tl�*1qD����ۆ�栎C�MC�}�� �3N2�i��f��C���w.D�DA=������
>����B>��a�}˞v���Dv��WT�Gfn��u1�L@�j���"�����Db-hx]�	�r�>��D���!��K؋�\.�㼜��?]�y��u�Y۪kd*_y�8d����8ؒ9$��	I,i�G5p40����G�Ȫ&h?_��?F$S_W!s�T��E�#K1a|���:t�!j	$:;�3>�"SH{¯�"�B`�fi2e��W�%/n�lC�ݸ(�]qQɞX�2�.[��	R��#wӠ��3Ȁ{.}0����5��ɯ��G�d�]����tm�]x�!]�͘�U�<B��0h��f�d�"�
8����5'W(�0�{}�}����g]�2�N����OZ�z(q���~��^�4'�?ID���ECL�~V���l�3L�u>�AM����K�a��F}�ܙ�J����:Q|O���a:��<7Җ��+�D�D������Dǳ�K���!�:d�KᯣC��a8��Ƀ�s8�67qf����-[�Gw����d�x�c�ad}�;j�P���,i�!�#B�˹��FQ��6�洳���f,��4�0��'2�Y^"��!E���M!8����8�#�NL�tVE|� akH�Ȭ�TW~��j��������2(��?Hn����5�7�j�j�R�_a��=��w'����u�44h>��]9s�d�o!{�����:w}���my�Y�[�Lwh�c�A������c@-p`sVD ��w��v�[���he2H5a�e��G29��6��;��=h�ҳ�Aě��c�6�4jƓC��Р,plf6yx��^�nЭ��ŮX���l���<]�\�K��m��e��3q�fR2Ǫ4�M`kh�7b�a�,�2��A`@����Lk�k��<�d1�9��v�vx��h�"S(�n-�d��h���g�X���^0i0�u����y�i���{Cf�L��!i�$H�)8�>�DY�8��<=���N��(�E��=�CO�k&������bc	8��|d�x�`�#u}�ע���.�!����8GͤI�$�L��p�[����zh3��������4C!�f*�D�u?20��n��#�m!_����u	�;��ػv����7:WI�P6�)Jfj�!#N6C�g��e?{P��J��_��P�~��%�k�w���3�Ț鯰��2���|���b:Q���pq-pDѧ�ꭊ#ƒ&�d��H����}�A�v��j�l�g��F#tn��D��E}慚��S��C�B��SN��H�dMU�[��w+�a�jX�*5��{�L�:�gƱ��|��84�i�*[�?_���j����]Y\㾅U"��ٗ{�f�1��W1�a�L�i���� \�����^
��Q�F��*�_����=�1��{f����B��H��dWծ�0�4�\����cA�/���>v�2�B_��H�3�x?.��|b ��FA������^�H�_���y�%����DV{�f���`�q'"�.����h~�i����i�� ��L�N�oiU���5om� �C��wD��b�d��"d����ql1�{��Dq��ݾ�[Y��")�{&���Q�Gq�\�'�����w���O�H�w9`�Tq([p���Xid@O�_�I�P�5g�s���|C3�4�k֤y�4����f��>������]i�������0�I�"T�I)3bc���!U|J� �gR+��4,�$��Y�E�{&����,�d;�z+�,��Lfe{�2qg�>�%���"qYd�{�D��R4��"�I���k�/5�~Ȭ:zP�F����T[Y���,�H�^保�5v5�#�ZF���[�;璼f�j��������� ��y.�P��$^����݆��Ig�z9N��k����@Q��4���˅�>��!�"�T/��"��gM��k��H���P��Y����_�ƫHϲ��*�����U̽��Uaj��O|BФr�eHJTȿ����G��qa��/�zTM<|B,�.p;����
,�<F"�w���VG�������"]����NLO��	�)E$pX�L�>"�7>�&WAᯟX��9=�PZ������ȳJ��1L��C�30R	����w�����e<M�WV�
����qps�v(ju���:��.����Z�FT�Dx�!���B�(���_\���"�XF�ga���)�Qp����uæ��xz��p̃�h��qY顜�C?Q�N�}��!Dx��<59�h������ߵB<U�*<�!��~��G��>�p����Ƅ-0�-F�ff+�HÄi���{l��DBn�Eh��5�B�}m~����4;�B�#�{+����.j�hi��2�'m�����Ub�e�R�m��m�h��#�����u�Ϋ���J]�b�[e��$m���҄5����)�h���'P}_Y��;�w5�ZFC���w����H>'>�~�/6�׵E����a�߹�[NBR��q��V=8Y�=�vo�o�jCHI��~d3��צ���:~���:��"O�idM���X(i�>�3��p2���nXө�@�FF�)D�}e�?2(�.���a���k�:}�xk�hIR��:~�Vz(q�,�!N��w��a�G�d���/A2���Q��NKj�^�Z�����D�?c������!Ĝ3Ht{�-}-B7hM�� ��C"���<Ϡ{��EB�/�K$g��$�k�V�����c���!}�OM�ٍc+ڟQ%)!���8����*��N�2�f����K5��4�%�0pz��IF4�N"�j82�C5�B3�~�{烧�a�����f�|W< �&a�u���|���M��aB4G���#HT��(��s�sTO��X�e��A##A�d#Eʢs��yxwA��㲕�u���x��;�'h#1n����/B��_9ފ�ӧ�`a��{�B�}f��C��1@�tV��qf�Fb��V⇹W��g;~�B�0��a(c��5xb��!3�@1��鱤�����`dY��w+b��B��yx�2F��4��D"/��׊"�����+�C#ő̾喝�q��d��`�#��#����ȓ�jk�e{�A���[ձ!�"p\9��͠�������(���V?}���^��������m�P�&8�xl�{�؈���3[w�ņIBդ�8f�ފ��dz�"����5��F�Z�=݁}QNv�b�A��ij��$��9n$�E��p�������>r]i醴�;��8~AB��k^f�i��U]�>�W�äY�4�����b���0�4t�Mxyq�����
?�4��Wz��#���=�}4c/Mğ���eB����C}<��=t�z<�����#7�Czk���n����C�u�o�n�T��I���w��� ��vp�Ӳ۞��iq���8YʴrӞ2�7gv.g �%���f�<��mqz};�����1\�m�!l,HT���"f��i��p �]�s�F����P:*0��{n��k�@��6�k'"�u�^%��nC�n���qӓ�Eo'��s�vA;^�Oe�����H�=p�l\�k.ư��-�``+Vř��JQ�gZȔF¶J���E�b�]^O0����n�w@,�ٍiĸ��l�8��ē��#�n��S;��`��0����R��zk�D��?z��*��9g���da�3|3&��6W͔�a���%���i���:A,���C�g���q��&�qIֈ�~UU#ڕ�o��p�=�tq�RqY0h�(���~���僫���K+�MYF����DI��QE ���$!~���Ɨ�C?Y�Y��iF˥���<�g�5�\Б��0�G���Y�`�/����OߌQ�̅��H��:G�,#�v���A%Dh�ec����a�?E�3��^����������`�:��0�dG9��M'���r�r�힚�8F^��p}�B�-H"`08�p�\hY���d��$I���}�b��!�2ï^�+�hI->6h��^�~�C&���zk�F�M�#���˟{�����6CI8�܆ۛ�gl\�͸*ۣ�{]�v9��v(�\��6�Mb�\&_�������t� ���_�D��:ԑ��P�_Qe��7��B�aK�D��$fF�'u��g�̖�)�B!��>,|�D�!�܎ƞ��F����0��4_Ou?�H^����u�+s?�d��Aou<�k��6�^��;.u�)��]�1z���\CC�V2=x�
�d��fw���;��ɯ�>#�ÄZ������v�#���_i&���+�C���o�D�h7J2�M�cN�kfAh^x{b�dA��͙�1{*X�P���>߲g�7M[?0���a���H����f�k"!�?��� I��&
D��Ϭ���{�	��xR��������>��}�p(��x��eϢ�j��@db�o��]�"��n�:B�]=<5y|K�Q@Zq�
�'$��d#di�B��]�������F����
�tX<T��i�#=/��H�\��U����t���""z����I^���ިEBˡ�\1-b+5�k�6�-�<�-'���l7n1�gdR�m[
���H����m�P�TD!��d_{�&�����R6z���hF�Kč�˹���z�!�#���u[�04�q���DD�6�JAc�U��P�~���e���0���x<<C����^M����}v���E}�AGN��z�ދ�ˏ���Z��7�H�h��/f/�0)R'1�gH���?}�%�8D#������^�� *���lL�Jl�L�$���6,eSy��s_L�d6^I�0±�!�gg6���������^m�N��p���Y�G���v�1S^�l��c�$U-��Gv���ko�x�����)�^cƚz���ZrorQ���_��~�M���P9jT����V�#��/b3n6Yծxg�OVقw1Wj��R,.'N����E��t刉��0wu5yo����ܚ�5�!�1��lY��3G�n�)��{����A�nD��\���|�o>K���?��Ŵy��Ӆi\�ɭ�����q�}0���E�K\:�t�%�&���ټ����2e��Srѓ�$�qi9����0D�51��x�v��������Ruq��D:��L��ߞ�:`Χ�S�I0~���5��Y�F�k��q�f���&Hp�����h$_=�
����ڻ<R�ǖ�|�,�V��QF�Y܂v���`<�5�r�5wv'��|�E@�ܩ���\��j�'dYuI�*��:	Ħ�a�ʗl����Sj��֐n/h��c+�jбT~8�7x�ݒ�ڶf�����\|&��ggB"]�Uu�%�;���Zɏ������Үy�,���n�����9.o%G�0�W;�(1�y�f��|�3|����,�=��2f�E�@�y��o?;�Ǭ�8E�n.*��f�X.Ƽ8uk�H���hlZZN��&�E��d�g��~0��;�f��V���8,mx�ۂ-�aC,k�9k��o�6�鷧p ��9����CW:{��n����؋��y:��F��*p��Z
���>���ͽ&����Lt�����:�i�Xk����*4L�� "BT�H�ā��g��~�K3y����?&�����CO�|Y��	y������Pd+'��o>�nd���e����=�����&C2D���25!D#�!dL%�h���a�+W�w��͉u�U5��E�/�+�4+\}�"p�{-����b��oz �;b{_�@����L	Fь6��N.n��f��;�{&�1�����t���j2�}Z�>�V����K2~Z�5�n��Q�L���z�P��C�<���a��&�E�?CH�dw�xK'��2n"��ZE���%�顇�g*�EhdY�H���_`"���da��r⸳����"]��@e���Ѓ�9\9�O�$�g��P��
9,{�Y�4��r�W�4�dC�Y�3��p����v/T�ӄE�䑦�B�[�C'D20�ȱ���MQg�ha�����%�Ðd	�܂��G�6�:�'�_Hv��n��B&���u� ��I�E>���F��=0�y3����$y�V2бyT$��d�ҡ-J�������Ͳ���z��kqe�&�b�gel;y���4.�b�fgd�"�{����k}���I'(��,��~�4�"��휟M���X~\���ܳH�
��͝�`���,Z�,�=���4�?i\}�\R�REHH��.N���
?�Y|8�%:��auD�v�jk�a���6}�f���h$���e�Z1���ȉ����0����4�!q}&��ߕ}z�l�K(Y�C����vF
�gJB6h�領�B��8l��4��|h��I�$�����z{�9Zg<%WsM&P���~�`�?��4�b߾<�0��G��\�y,i��16tJ����p�"J����M��[�ea���6,��=��	"�Ueq_K鯙BT�d}^�4�!q^����d��:���!�gC�;k�	E��I@�NGc�v,#J�\�D��&"��Y���ȓy�6Q�^M��#5"/~�򡜸�,Dd��`�k�����t]���k�<��}MFZ%9.�zp֑d?��ϮX�VF}���OY�5�xW�"���(���E�ꀆ�M���d2�>�0�ǫ܄zzz!^(���th�����&��cb��=�u�Fh�I�8g�
.�Ւho=�N^K�%2����F���WaǇ=|���C�:�5��)�Qt�-�Q�B`�eڪ�Z�qG�É��v.�d���h�n��%;`�W�0xY|�юr�2�&��]kb�>p�%�ǭ:�g��7���KW[k4���1��ۃ�F�z�n����\�����d�S$Ed����[Nҝ�qG	c��,R�Nn�� ��pAa��<��8�Ӱ�mq�k�XD���%H�x�{m����lr�S[�l�y�=i�fpX�tNvn$��F�m"ĉErxa`+�a����V~�г ���~������4<�to��Ho���G4/+�퇝7gƬ�Ä\����a�$-D�p_�dYw�F��Ek��_#��"�WK�wF��s�X�!���3�},N*��i�#���w�GH�Νs�ݦ|p���C�S�
�7����dvQ�z��g��?Uuzha�|�3��$�1��2�O���>6t���ܗ��R��U�X}���K�TN0܊%	����4~q>��]s8Vh�<�D9��CM�Di�����z+�rhM�4p���o���Y�4�����nq����]i�=8i?g
0��7Bd���l�?Q�W�E�Q9z"�QwU�N��cӎ����!>�s��HgڇH�S.�v8k��Ba!�#�>?`�
���61�oTɧ]U�[q�֞�'W ��w �Ćw.�ݢ���:�sA=�����k�C����4����VX>���3�CH�ȳ�OW��Y2������#�d�h�����Di
�ik�i%�@�!2�v>�,�CO��
������,�7{�lMt�_�A�����w�*�a�/�퓖�N�,n��VI�]칸0��f��$	a����1Þ����G ��������c�y�buU�N�~�;*� ��|U��{�U~L�S�qM.�bġ`�Ώ"ԠЌ'
NL����i5n{�c���|UQ�V��H�<#B0Y�����A���!��3�/&��3�e���Ш��O�"J^'DN)p�S�u8F�4�]!l�n�#+�zo�"OըQ�w�P:������{�ab�P�]#vn��2��{�v�X�Y��Y	
@�1�.�C5�_!��2|�N�xD���w��]+�hIt�7(vE�P�C��dh8G���v"-}����w��=]m>�Y�������[#F͓C�/C��61x߱��N6��\X��fwl��ӗiz�̕(Bː|>#N�W��_߻2�~��O�adb�zX�#�������Sr��k�9�c������ϳ��M���08��L,��Y>��v4��~dȲ4�D]���Cr,�������Xᩁ5d[��K�#���V�����ۮ��_S�p���MB;��G��+HdI��������P�_Y�=�tb{��A�kU^�Ǐ֑��Tǖ��;��3�.3��!�$�~������n)�t`����*��lA��b:������D���?:��$�$a��C��8��lHmJQ�#���,5���(zMl�U�b�"���70�k흁�@:E�E[���xޠȁ�S����桤9n���E�=q�\ۂ0�����MY��.���KP�cOZ){�X{۱AGG�`�8C�ߕ�ȳ`20�^�hwe����ip�~�7�u�j`��,��t��r:t�3�uθCq�՗����RB�ܸņpA�#�eH�h�����8k�Y6�����a�N�h���RGK"�=�>�Q#	4�s�YhCVE����#�r�i�������ɱ*��y=��,�{�'�/�ǋ/�Ejޛ��ѓ����aq�/�s�c3�ޚdc��K��x�F�����g������w1�+���2A��Yж�J!1��gH�>:F�i���;j��ã=��̮��Z���rKi�,�0�K�+�����=�g���P�>�rW�_Y5��5��L�TeBc
2�4�#L�f/y�88B�/�ɕ���4,д�衇�RSJ5}:����la�6Ӡ�"���ܣ�*&�c�E����� ޟ��,����\����=���=�0n16���YP�潅�_OG{�@�!���Q	aX#���N���|c�/���Mv!����`��p2�1$��ޫ5�����ݵcLai�=]i�WB�P!�T��"O�Qd�h��H���g�8N�w�Ş#�|��K��Y�(��� �L�)DHv4t�� �¤�(�f���n���G�L���i����Dr0�F�i�+�N!/�}��kz��}�5�y��x��G&8y�9����< ��^z�����|���D.��4����>�A%#HH�i�_2��D��=�}�� {˺4i�}֯6;:�k�"��H����Ҥ^#q!��/�~b�A�Xs>g�M�9ڲ�!ϭSh �!�������͟�;��}�A�H�r#KΥ#�%�@G��~�@�V��Q�4�f�G���X�ڄ�\"���KI7�i�n$��]=���%��7cm��+5�Ȗ� '����hSR�����g=$5�E���qu�ݡ����M���/�V�1B,�5~�����HԧnH,i�#�������k�C^"C��U�Q+"����~��i��]�ޛ���#�]��ϾR5��4��8�xe�􌌕��Kr���t�Ӱ�`D+�T2)��g̨�]��@�#�^�ޢg�pw���>#�g��ܬj�%|�|���m>AQ�Ȑ�Ȍ��,�䴹ܧh��i�.��̣u�x�3mmtt�q�Eu�c�c��ܘ�rkp�v6Q��&�l��L�˦��(`	��Z�%��cKk��m��68G>��tQ�]�soF�k��B
��-�-×N�8��Ո�T�gh�˝z�
6�x���a]CB��A�V�a3b��A�VK<zd��B�c��������ny�[l
��7%�n��H�gm�n�E��3��U�l,��/�U��D=�;#�dej�#=��%֐�YxJ�S��Av����՝n�d#�}��+$i��5�3ı"I��1����ڂ��i�"�y{镥�w~+� z��>߼k"xA�_����<4���o�.��YF��^��;�xiC�!x�<�种�x�G�~>ބ�(�n#F&+�"فa�	�����z�����^��ȓ�t�P�A�3Y�A�#k�(>�́�>,��}�}/�x��������cC���d�G�O����l=P��Dj	dE�?
�H�/�B��ʯEj��~��x��Y������&7�&"#�^�S��K��������#�
m�M��W[�j��0���X�XF���!zfR�������@�q`s�qCH�Q�'Hg�z�Vj�?3�^�x��@"8t1k�`��E&�^fe]�,�s6� ��4^���A��+F���"�Y���������Y�p�=�xs��w�,�ė�˽V(i�̜?T!��畊�z�r{��`�g�� R��衧�CHg��~%�L*���T��N�l����,��z(3o}�m�ҷ�W/I!^H�[�wo>bq,?mb
�N^��\��<������4n�/�"��f����������x���m���Z̷8����+_i��W�p,�,�=�؛���#H�|������g��d�`����x�d>Ub����#m��1�ۂ�5}���i��u�t�k>�(����������~l����r`<���e�fB�����������8�i��|�C@���2L�"����U�"�~j�q�;i�����h��+�Y��"�W�]��b�CyB�7l�I������d<��H��Gf��e$�
$1�౤`8F���x�>��.�Y�\"�}>���ߜ3A[|�+�C?Q��(I�(�]
"���S�4�#�`Մ_>��fԇ��e������N�ش��r.1�� ��ʽ7��֚N�	۶����OZ8g�mK�[H����2~`�"�u�
h�"�}f�vߕ�ޱf�E���pX��N�˫#H�Ⱦ��^o�#O�a��I��MƢ4�S$���:F�N�#����/�y�p���|E��iq���a�}�r��v���i���?3e��s�b����Zǳ�!Z�Ni��Tw�(��IP�8�mD����f��,�{��tX�F4�R���Mi��<��D�*h��x�h��#C��0[������KM�XZ�85���B�h=�|r���T#9��ݛ�y�<�Wi|e���{�Q��������@M��`�d)_aK^��\c�6B��X���:B��ѭr���&D�w�ו�uY��0���
����$Q�A�sʂ,�?i�r��>�r���<�T{���\��a²3�\H���h� FB\��#��5�Y�B���A�F@�t}d�S�z|k�Bȩ^�0����
|�!��!���i���W�fa�8�sܪ��������cl����qÝj��(ش���:�W$�5!�Q&l��ZW9l�����Y����+��h��,��z�X�UB��4�g�累�d��������Fr��A���?I��P�JJD��m�����t�"Q�>�v8fA�r2���D���Ξ������	"�"�`B}3�����~�#��W�ELv6b���������:J����d�!-�H��VGs��̬����%��=�x�
�TƦ��j����ll^��Pdi���qH��K��)VB�?}�H�nB�eD�y]<��<�s�l ��<ş���Pf��+�_Y�r��ȣ��G܁�V
~�p4��^��r^!���o��iwg���(a�����\3E���n�8����/�9���Lc�Gc��se�]n��	��M�[�ۘ�T����F��MikN�������C�i�RH�x8F�p�E��߶�H����l��q���h��Y _�����C/�ib:�}z-��������j�w�`"K ��%iq7��+��(ʲ�M��õ�P�X�UsN�iB�!5����b��-�.�L.�ެ���CB>�ދa����J�����d^�E�FeuEd!
��F���]C!�#�{�u�=�H�K;���e	��p�h����8B�����&�F�m�nسK���Xm/�T#�r���"O�t�\|��b���<��ݪd<SK��f��cFSL��!R�NK�f��xA�\w�Kj���Y�?�.��#��8@��sIxDR���+����#d>���CH������Ň�Q5�6�!�#��#����������G6~M0Dw������l��w���da���g�2SR����v��:�H`��>e�(Q�#-8.����H��3W7/�cz���_Y�4�}�	6�-�_YD�Zx��=�b���� �Mi���ʓ�""��^"zB����q���#��gW����X��Zwp����z1�����Zu�%�e�V�ts~���$n����q��8���1���. M�V�yq�_]Y4Cʩ���M-��xn�#
���wd��0�w�{��٣=[����F�_{l�~Z��e�"�8^���������O�Î8T�7ln��|Fn�E�yEE�rc(\����'+�,�%�<��$h�6�ޞԺ1�X��\I�,����&2˫3�������z���� R���E��m�hB�WX\��EN=H���[�xڧ�c5��������x�ı4M�$|)=	�l6�Ii�̷�"�tSː���.��2���^��M��͚9�8�4L� s��f���_��Y��n��<1��Z��}����.�׈ќ�����;�;w��Z}����4�0�qU�\4����~�h]jpf<����r�2r�SLf}Ue����,5f��=�_�p��G�+讽[W{s��̝ފ��}�~�����C'_�}�T4C>�b�(&��v�S-c��n#�;��i��D[g`�	��oR��4��{g��R�k��gy��M�w���m%6Eޖ"�m�	f�K�P��M���^� �J����ϗ1�G�\���>�MIT�҈�4�K�Z�ʭ���f�/~Mǋ������\4T�
�*Y�JW�!��kp�j Y�We��dWfos�x]�=�ㄓ������`j��NMzx�ċ�8��ݵA-��6��翫�� � UR���(*����  &��9�f�nMx��'g�'�&� ��fVX5��]�afQ�y1��ɭ�tj8R�a�V��6��0�[fF�6x��N�e
	�>��i�h�)w8n�Ttw5�k=���z(Lz�{�s�
n؆,��дrL֗#4	��k1nx��%D�I���-��)�ran)X�n���L�$�L�t�Z��f��Rl��e.�m٤�2���h�����(8���(��3Iv��u]r]Vunr����κR�`&#�l]�zSs�s�;#'r��5�'n��;0���[
cB��Jf[.��`iX\kpi��y4���e'j)R�u����U����Dg�����0[`�$�]��T���apic���Ͱ+;����Q�V�������jǌ{g�������ɓ��(v�c;G,X�D�Z����A�ٰ&Ϲ���8Jɓ���q��6{$��g���>{������v]�#��
N6Y	8���M&���=�{Y΢`�u�Y�'Ov:�;
�.�u��*��RƆ*Zm�0I��ѹ:'&|��!�u�t��_�n����v�T`u׆1��{JM]�f�d̳35�dDBb�Ďr�Ng��v��+j ��nՈ�ٻ�b+���B\���n�����f#��6�l΄�6u�qh�����Rv2��k���õ�n�9vv�B\
+.�C2����q��R;�v�Z"�#��t5$��⺚1�ݞ�mQm����:FX����r4Hu3^L6�L��Y�`����{��uña��tc�s��hZ��%l,i���2��Ʋ�/b�&�{iB�ZÁ�f��,.���ɼҤ��{Ff��=����Ȇ�U	�`��d�0.�7�U�yxm��e���s��;�5t֋�V��̋I�*�M.^͗K�A�u&�u�is�s���݈��o"�˛ڭ�r�V�1.e�K���44�l��,RMsqDs��k��E٧g�wS���.랹��hnM:e�ew�9��V<ru�V%�1���K���G�J��F��7�!�5FH������Csō�L�֗W.7f�@�����v9����Gmj�ru7\�qtc�\^؛��eq���6t�9������m�+l�ЛU۩�ۧh'o)����oYG�gr���بZ��!���	����l�+���KnM���A)*�;�js�5�8��ٜ'@j�tonA��Eʼ�a�P���f7J�U�% ��H�px}�a�T�0����^�Һ*�~#�\�y9+�CYX}��7ˌ?Yp��8����ʷ4�4�԰��}&�G	8$!�r���7�4�=��A��V �B?i�]�UX3X�7��i�h���[~c����ɯ��W{���� �L2���5�0ڑ��F�)�c�a�4�!�O�����W̌6E{o}.2��Gm�E*؅����w����3�	�ъ�����@b!�a����@S�6"����pZ��H�R��5�G��:F����]�_iF>6r�9}�A���"�wzB�#=w!�8���8~W�V8aN��DČ���>�װi��w��˲����a<]��LP�����gя=���HeZE�[��4Ռ�(���sj�%$�&�O�L��)(��Kf�SL-�����о6^�mb	�5�׈�%����#��*I�gO�{�p�NOz(a�6����.}�(Yn a��i�v��B*ҞBq���H���w����4��w�/�����k+��eH�FGa�$`:��q0�#���u��,��ߏ�J;�$��5��Ջ����7�"A,���xt��_{}m|�b��Bۛ���vy���%�e>���:US����*z��F��%�C�m�g젆ufM:E���da�2_E;H�
1Ψ�((k����a�4{^4a-Cf#!-Ƥ��5�,���~���G`N$fTfA�{�"H�9@#ܾ^��+T���as]r4�}��ZF��K�z��"bi�%� ��>��#S��<�4�Bфw��k�E����O'��i�8xj����H���#�X@�ڿ��Ƞ��F���$T(��&�Q��	0�:���w٢ƚ����z����˚��DE=��A������^��l�"ψdi�ۛEU��5ޡ �{�X �j\�ݶ�7�5Z��k�� �س��,���]�$�rnL��M$�G��VG�����������X�`y�8��ퟴ�.?2#�kEq�ŰH R͛2�/����]�cH��C��<�_�6M���ȃ��(�|�X({W�����	��K1K�/Wz��_X�,�ȣ$R�tP�l}�i���w�T��T��Y>��^���A唍!���
���!`���0�(��z,x�$���Y�"c�(F/�����q�T-Y􉵰����[Љ^N�EW�)��yK���M�_�D���T�D���f�P�E��A�Rs�\`�����m�|l]��u�!�F����ע�:j���'`��!?�&QFS�+A�wX���t��zE�]�;5d`�,�>�E֑f��t���,j�#H�P"B#f���(�L��4���a����N
|k�H��BF{s�_=L���6w��l|.yhU��C�Ȗ~��+=�鿙d�tů�_z6�$�׈i֑������?����$�NR9�3��׵u��5��	Z�d[M�f��i�T��"R4�i����j�G_��ۚ�i�D#�U���{4]o
�t�4�=�`�����4H��n���Li��<!���B3�tA�]0�үC�	��A3!r0ӂ�̥dp�0�s���[���릆u��5~C��ϼ�_?9\#Ms��X�t�5�P���ܿ��i�Ѻ��Q�!�B�pS�(�d������B�y��}���p�ƺ����ϕ�V�dq�JT�G�_�$����ޏ��d.XE�צ�4���4l�~�a��iD`*A���qp�9{2���f����r�0��Ό�#pm!e�;����gO�Q~�(`,�5�2<��.��}�NM�_���.@���k�:>�.'��f"�q�!��q{�Ny�楥r]�<�<�w��[��؃�xW�w-�m�'�3��l饈p��c�����#��R�����h�Ñ�L�z=�(q�D"1�J�y��-�H��̟K���5�,���4����#�,�4��$٫��$�k�"�ŸI0K�]Ө�'N�LO�2���;]yѠ*�a6�gF!��qfD:�E=϶y[>�g�3xvh��ȓ�����O�P���ai����lX��H��L�?If���^�[w��CH��=��Z�N����ZY��ˑ�q1^qA���s�#H$G���UaD�6k��0��Q�A�NE?CA�`��ފ�4��C$��}fQ4���K�Ɣ8�l� ��6��YB�k��!�"��e��E����/���K�wl_�����5�A�n~��d�Z��A\Yp���@��A*"1)$7ZF�_�l��#��w�<�ő�Ua���]i��t�>!��>#���#��mē�Y�k�1�C�3]0٬Y=�:_
�&�܃�H������ϳ~�]>8k�Y��9S���������i��=>xhidY�4���o�Q]~�ZYt���D��a򞳕7dG�Q*��+�:C��	�~O�9��_�����7����yk/`;&D��"�8�L Ѽs�KY��s�.��8GS�_Kn7Dc���q�u8�6͌:vᳮ�h�#Ҽ�B��rn�v/����bS��Aa��ܘ���Y��x~9��۱ݵ�Ǯ��B�0D�%�d�*2�kv˦���^ƙ��'&�ѓ+�`���A�l��NZ��΢�yl���݆��a�;��[�G��ܥ�,ue�5b�һM6JdV=J@��B��͌͢�JԳc�J��hbl�Z�Fk�.�y���s[�R�^Mu�zۧ���`���U�!�y�hU����6+�^�?��jB1��b���,���D���MRα؄����h�܄ܬ�F4�����%�F4����xi:����(�a��X�#MY��7��:����/��g��/9X��%f���>�(h,�0F�M����(i�3���	j]�Ћ#�_lp�?|Di�$h�rr�w�xi��!���ƚ�!����Y�W�k�u� ��&�7�C�`�U�Ma���hܥu{�T���ZF���	(�@�P0Ԋ�uZ�1Af� |fk�GK���FWO(�\}c�O?�Xu�����43��˯����Dud ��I�,��K�$i�1��!�H���DS�뇧�U�Rp�8��4������hh$A��G���q#OHÔG�2Ս�Yb4�¸E�b���T��Sjq}����h#�#��y}_w�&�h����;Q����[Λs�!Յ�NX���TV^qy�n�ls�����,�(x�Ӟ�net�٭"�����C�2������"=}��m��wΐ�a52}�vxibj�"�	�����i��]<��*�CG�ϭP�}��g�oy�^;��ɗU)�T��8Z���Y�rg�+�v�q�
^!K�Y��V���n�F�/�I�{�cyk�yǜ\����߂�Wa����+�Dl�,��y���Ha����_M|��,��pG�h��ϰ��H?��+�DCD�\�5!�u����A�����w��M��>��9>ȦY�Z�����H�?VLU�,�Q�F�W�=�j���CH�xE�'wȲW�F�)Ee�+������g��g�h�#3y��?Y��:���,�#K"��>�4'�!pۋ�K7�{�O%��8l��Mnޯ�m�#L�bH[��"��4�fA�޵�/�pXt���a�3\�㔰{ҡ��|��a���BƦE2��g������">8G{/MB�&�R��4�v�H&� ��y9�w\��h9:.��,��G@��I�f���܄��!G'kN�a���0K˛�CK"Hg�"�u鯰�Rt�=(\e����)�gN��(&�/�0����Ei�p��ӆ��߶��S*&��8ʙX0�,�Ց���1_cO���$LtJؖ����aK��}4������1دE�ȳ�K(�/�xkx�?'z0�@���r�"Gd�j�_j
�oܸ8E����v>�da�t�����:1�՟�9'��vb3�>��86|\Z���M�|��f7���s��5��V��?[����vvk|���@��|�T/4|�����o��q�#�쬋�i�xފ��E������A$29$,6[�X����15�*�@B������?K�����u{0�m}&�q�%Ɲ������P�;�_��[��Z~�4�6Fǫ�����
G$��Æ�#���G��v(cA!V��n��d�� >Y�9�诰F�G�"�b��P���A�Fȷ��c��;�C�w+M|G���ma�Ż(l杩g�J�G
{V��uȜ�V91n��mh�[T�6�.��ş/�,�����+O�V��1�'�x:j�?R���m�ܔHX�6�Her��]�f;5�l�x�_G�IĜ�G2f`̋�Q���p��Uy�����4uV��:��"��eg>cCZD��Y�x���@p��ȝ,�@�yqJ'��=7�f�\kl�Y@��ɘ���#�t��f;��ϕ���,�VD�;܊��U�;�H�2�����@�I���YtF��:���Y?j�44�5�Y�|�����
rL���5��o!���D�s48��(�k�Т��Λ��!�oH�O�v4��j�w�5�nz}�D|x]�ө;h�&c����cf`�>�Y��W�^�J,3?#�4V�Ք����=�2�#��E�s׈��igw���J#��P@c���di�0�}�΋�:a/�a�3�� �ҾSD�|>��p�w�~�{F!�x�����
G�YP˶��}=��5Ty�#��a�^j:?y%>�=�	��s��V���%�l<Z3�Q�ڷd֦�P��&.������6k�5n~�X�����V~�}��!�YzP���P�xP<n>�
H�&e��4}��4EZp�x/��fB�h�NF[���4��0��o>�������% ;�F�Y�7z�k�9��B���п."��\׶h��M���x�
\�%�3B���bL8i��pea���[��`�߹nƖD �ue���٢���z�X).�!�"s'N��ۀ�Ȋ�M}�:_iÆ���E���0)�Hli
c�8W:�Ⱦ�0����dm�y�s�D��\1�dWd���a���G�����(�Αw�H$�@��׮�)��~�-"�u3�K	|�rZ2FCpeiᆵ��aiw���h��4���/�!A ٚ~����Vt�"h�FRy١C��9H71�g��58�"��d��6����棾��5˝�)�B��"�	
��R�L`�N��/*.؏���џ3w**\j&U�ޞ��M�B1�b����<Hgh��݊5;\^,��/5�@u��&f��-Yӄ��^-��.e�\�Fl��j���K��[uWh�� r	�+��#c�[S	L�Tw ʦ�X��e���j���e�c��r&}�p�uB�`��
�v���{g�gn�k+�z�G�4�Ԗ�J�\��,c��m�#a���f�e�a�<j�L$���������&���\u<٣�DI��x�\�tJ��]Z�e'�=�A��%m7]���E��4��$�>G�~;ha���.��B���0�ϟqX�UaU+C��E>�s�y� ��C��1衧�0�DH�?�f4�(�qɃ�ӧN�����hi���}d[\E�DQ�M�u5Gu�p�qt�ձo淚<�i�N}��F�U\+K4�m�*eY��5V�Q��N"�V4�!��A����|9^!���A���`�:¸���o�ێm��Z�}4,�l�47'g���M���HD4��\�_A#H7"@��+N�Xi�	m%��<=Ũh�_v��l2H�3PF�����_i~�$߂��f���A��m/�??#���)�#H��:g�Mh@p���P9$F2�dPdz����X������4~�8g&!onR0������,�+�&��g��h2H�_-B���ޚv?n���ZFg(Y�0��J,6q��i�`�͢�k2�K����Y��.
���4HBT�,&e���kM*��7�:F�Ç���������5V~gE�a�,֞�~�P�O���|�oȎ?Q�w[�BΑ}��oe���2�F@S�?A`�!z_��Óձ�(�i�.p�\c����#���ϖk�K�����6�,\`!��q�R@7��Z?�X�x8)on��<���-��5���w�������4E��Mx�2Y��z�_��Y`-!g�z�8L�LM�}�4�����G$����F@c1"f�Ϭ�d�.��LPg�4Ց���C�!�Ȱ��V��8B:D����FȦ�`!"/՞��~���k�������M��������XG�&A��0����]x��ZE��[��鰇��V�f�C>��XC5�fW�=��h�<W}w9 �.v"�W��P�aRG���}��c!|���li�"�U���\ϰ��m�̚9�a�dY�z�cOʲ�d���b��hwT}���܂
��1�5%.^�/0`Xk�ڒݜ ��d2=�M����&�8�M�9�e��l�do����{7hY��X���z,�drat	�k 5�����q��/�C���4��CKIX"��W����`�5��"�l|[a!�$��k�B��y����ݾ$����d8����_]lG�&E���oa�������=��z �ˠ� �r��5|��	�H� QB[������5�e��镧�ω,�9hy�]��>u;�>�$}�>u�ՇcW_���tC���3w[O��ޙ��(�#x�k3oL�tvw�Ɔ敷z�=�����_K6[핬����%�U���#P]��ޅUӲ.�k�އ�s�KQ�Q�{�Xr�l�v��ي_[������o�_l����x{="�������G���y�8��wj
�=�O�O�燏�S
잃��l�{'x��E��s�U���L�ǻ�U��������9�bd��ϳ�F�9�-��WXQk'�+����K��SD�8���J%�	�Wr���U����$����ܑ��KƝ��֖�$�@{b3vo`ɵ�@�Ĕ62�[y4��vv�Vx-��2�"��HH{�z�l]�G\���fg0��V[1:�'��:## DF��t��Y�����젓���5��$��c8ˑw�̬0�\�o��;{Ǻ�9��׼3�|���m��zjB�9$B�}�rԷJfVo����f�/�A>��Z7�Y���R�)��`��}�A�b�V2��^֕�"��7S��sh��I���m*zvz;&R���q=���|S�� �v�:\޿;x�wgC	U�����;j�F_��:���rx.��D��0��>�x%�3�/v�[�VD�ˤ����l����; ���8Lk��G_����W5�-p���<�����A��j�~�8�'/Kld;�k�)�x.F�rT����ȥ��/a���3ɱZ�.h�s��ɝe��w�ܬ�W뢋ar�垬�e����*U��X��
EI��N�=8k�sڻ�@8��20qJ��~�4�&��7���v�"O:f���C�1��C#z�%P���d�;����:�5,Ok��1�ԅ�Ri��z��;ϹϦ=:t��%�k�U�|��K��\�Q�WI�{�W̊,4	n>���T||�")��A��I��@d3�jK����퐞��5��+ -4�{$Cn��5�v9�ٔ�ɳN;y�Q��S�p�]r����O�*_/!dS
c�b�,��3�5��迥�G�EC�e�
��R�|�/��@�+f4��V�DdY��7kM�+�����*"��H�����4�!�0}}��]O�]�;��hI�B�U*#]Y�MfR}�4X�;�Q#/���d��g��#��{�H��䁁U��$�1��8��t�:Gx�g�w�l�p�2Kq�i���_{�Y?��Xr��R����g�4�#��1UӤ��AL8k����P�1$�f6�2�2*��&sZ �B�/�^�<�-Cة���c�]p��<�C��5аY`��x�����{b0�����&�����/�|`Z��ܼd9�j���w	��s�\�#p{�!٢Ц6.�e�I��x3V):��{��{���U;CHg���|`R�q��I�xGOOt�5w=��Ö�����0���6`�n&��{Ͻl_��~�T�މ�Ab�c�=�3�/x���B�Ui`٫�.s��Gąeq6S��M4��nVL�,��8f �3ۭD�c~����[�Gh̸�e@��vub,���?z��g�B>c��ו�ҳ\�c�F�J���c��ŇO��g�}43J�o��Ԅ�����}7U�T�p0�d��=�(�Sm%���Zk�!�:�ۼ�cO��a�^G�V�y�z.��F�4,����5}da���8���.������崓F2Cq(�rC�M3���y�"o��L��f��f�����`�".�y��׏�T�����כf������k�_�����,��j���Y�H"i�#2���t��i�#���g�9�0��#W�_�<�\Pµ�� lْ!w�����C�Tki���E�������"�f��#���I�$rG�H�ç�Ȳ-�]ϕ�,֬?!���P�E���l�����Al~�G��ء�����A�����pbM!�sP���{��b�����_�ʼ�����.����Z�dD2!���<�j�k. �g�qM�x�+T��!��bɧ��A��j[��X8�zݞ�XH� �=�����At�7ێ�BZ@��v��J�QͶĕ��l��&��i�JW�u)
�*���E��%Cimq�����G��sD��;� ���6�S���cr���i4]�&�� 4s5.�I���6�BOn���u��W�O��Nøy���l.�m����*d��nخW��t�7Inz�])�۱gd�7OA��g"@j.؄��J�.e��� �C3kMe�R��nv"��"RhVق�Սhb��{c#��K$WM��~��?~�<���,���"�=鯏��"O��>٭*��C*���(��t��{��#��A�`8io��Y�ɐ�L�AR,�'g�B��1_g.�{���>���&��X�����$��=�~��H�L�BX����g�}5�ń	��^�0g0�B��A�Ȋret�5��=2r��41��"ڲ0�u{�}܅[u�s�6�:r=�!�GӟZ����pD4��M�b���B��F$݊��!(�d)nC��ۀ4��yҮ/�X�$>����D�����9�^u���8��!qZ����,��U������w�o2j�)��lE��`�ip*l��06[��ǧ�p�}���7��ip��
r.�N[����L�"H��da�(w��;���Gb�+�nk���w���H2�$�s��1�������͕5]���i	yL�1��XK,�j�&{mj�%.<눬�;D��c�4�?4���#�A�}�>�4��V~dY�.*�M?Q�XC2�$��lP����=\Dp�0�x�뿸���Ӵ8k���I����0���+O8���Y����C
uٽ0v]�·�+��G�y�Q�Sf�UK������C3�Vl���Mٸ�qgO�
�Ca��/�s�`��c׸{����g��C�_Y��}�5�ÁG�"΂��h\�O�Q	�a�W5�y�
��Jl��7޹���p�{�0���L��d9,{PX��:aB�߾��r�D���i.C�=J���p��D��V`a?m�'�^�Y~�B�}ޚ�COުcH��G��AB��6Q�u�����$!�G�tI5)��A�<h��e��XY�s�u�!���s��a�VjhE��p���sH����lW�D��Hw���Q$��8��_�Hˤ�!"��q�>`+?_,0_����*�K��"���1Pc�H8���顴�~�,�}�T|5}Di����Cw�����6D�	O�V:ے�ev�h���i���}�'@v��,e�=�[qvo\7H�f6$eG'kK0׈�4������E���{��21�4D�*Z~�Nߕ��Г�I3���KB�;�s�x�;u��\5>���!�Q�����gg�Ç2��_^�a�P��k�y�e������?A6�PF��{�sC"�qA�V�QU�t��j�51���CΥ�Г@�`A����_U� �$N����PfAF���`�x�5�A<��`gN��n�nP�W������X��=�Lޫ��&�b�C.�E�,���T�D�V��Ͳy�_L��2����!��"��鬴4��%��Y5�o೴�P7M�)����Q��"HI
B�fd��rʳ��H�=�Ňa�×ۅ[�(AdI�BN�H3�_r��l��$�CMa�{�f���pHˇ���;�0����b��$Y�g�/��R���\�gCPl�#\C}熅���4��H��g�Ύ�HUj��lт�*�D6R��}�)�0����H+e���s����&�u������P�b�g7)�/`{[L�̱�CJd�!3�����'�Q�P���Pz��ŀ�_a�b��G���3����q�&ȿ�}�E/&~z�,�].�q�\JEI�'+�������@&��hiX�t\+��H������|�C���>:`�Y�4#V��?Y����i	���ސ��Iߑ��%���/BÁ�MF`�7��'˄3��@���g�5f��!���(!�i��|�"ψy|�mg^9�^�#�V��{lҥ��(i*ό���Qd��d�h�&������
O�rL",�s�C�x�Gd���{��|ȃ�4(�G�3Ƅ_T!�NR���Qf����ն7�V C0C��VF��|�����i¹>��I��`�H�T"�E\鼸j���G��1G�2eN��4B����0��UAH�ppa#z�#K���I���Z|p��7�@�s���l]sΝ�,������"�X��ȑ�I9]L�H]#L�:k�m��������,�ɓ���Յ����\�S`9[Nhq��3c�����a��+����Xj�l����;�4�����C�D+��̂�:د�|C"��h�<�g�_�F&�Ρ�z�!uۚ��g�t��'�+�C$�6䐧�#5YP���gܙ�3�P��3v/��z~dx�!�NM�������-Q�QbW��bH�=�]S�}�[�A�$<~��W������&�<nBTdC
2�|��ş� M� ϣ�P���7%ȓ�Nt_����v�fb'����1(/E١�㈸�Mp��o��^t�뎽�8j�O�!"p0 \)I,sPQp�7�WoD x���A<*34g�t? ԑ�dP�M�fML5��C���P��q�Xx�c��`�esw=�:is�-H�q����K(Jr6�F8�xl�X�c@�ﷇ�"V��w,\�8��A��v����=��4FWO�,2�8�����[�B�� ��s��{<G�Oe���T+���0��6�!�¼]Yi�.z�z�����7vR�}�Fèb���^�=��~	3�>~�g!�s��e�Ġ,%;�l��E�覐x��7�ֻ���ɀV�ךx��}ѝۖ97=C=ttN���;����l�<q����M��Cpv���c�:s�Qxy�S��N��f\���R���jHs57[יf�z�v�$�KKWM
��9�z�KY�xP픞ܯ��l��i�{�A5�9�#��Zh1w���lb[�'��Z^�J.y�]�]���ݤ��N�xv2�-g[��,J�,Ή-&f�-�^�Gy͙փk���C�5�v�y��8��=��j��8G�N!��9~�w�����Y�a�!{4W��G�l��^@�m�P��[�V0����8pdi�����>�d-U��}��|�j���Iɜ$����s2+P0�O���v���Gyw|g!G̈�v����QY�fD��d�P��됃!"��;����'t��v ��i�^��'O�!���NH.Α6J�+U�{��W����FH>�Y���Q��9�`J� a���?m ��%�O�ᅞ�X�q�2��KgM,�k${� �p�`����<0����d�A?�h�(���C�Q�;��l��_^�4GF�u_������Ń��Ԍq5C�V�#�^��٥Y*�ظiO��C*H�e��I!��3$i�d�F�d�o�p�$IdY��C;:��^r�����x�=����x�fPf�GMg�Gܙ��g�#7hn�F�_W���c����Xe�F\GNUG�C���D[�[���FLE�s��aa�W�rH#i� r��{F��"EO��ˤ2���2����6D�(a�J�s���f����F�#yV׎������t�/�h��F���"	QGrKäY|(i��!3>������=��O;W�m��x��R�cS}�,U�e9�AN��&.�C�9J��b��4.^��|��u�i�q����hgzݞY	bf�_}��u�h:e5�[,У�p8�:DUy��Y�&�#�8��pt�G���H��h��2!	��zC:�!�~��c-�큄&�3}{鯣�'/�� ��H�DL�rhF8���B8ho���gOF*Gp+��|zβ���00\V�G�Ohj�!����Άk���b���>"W���:��:�����z(:Z�'B���Ӿ�(t��^xT��4��Qu�mC|�"��33���6Fj���hq�/��]?a2�Oh�sq�(x��ȍ^#L��Rl|�����W�����B����Ӧ��4�3�����)�Õ	��R�D5�5� p�,�lSt��pS�i�,��ؙm��&��'n����*!d+#�>|����I�g� ~�4X���j��y��M�>��������!D_! �Ϡ�N��	��P�|�<�H�8I��$��j�G�60�k��(,�}���} �VBG/���1o����p72Y`��{E�����dO���w����)W7�ù�+�i_6"�E"N8�pXޡ�ȍB͑��?�֟��P"1ă��]>��_Y=��O�5:$���� f�iGƭ�qf�'�ƼE��!�;ٽ@��7���e��������fS�{�uHt-yɷ��znN���巍��?Wdnc�bO���E���/>x�V��01dd	��H���E

T(Ơ�ӧ}���ޮ��f�s�H�]���a�"H��������د��ώ�V��0A�;4��q�BE��)2�ɫ���8KC��ܰ�j�����$��8R�^�"��]�u���/�sJ��hYVGu����K�d:�B�t,�/��/��چ�c|DU{_�!�����7R"��ج�������w�ڳ$���Ѝ˩��vy�Ҏ���-�tSzmv8�x�
�]���ō�:�3)@�f&8x��Da����}��v4�l��V�}~�]<=c���p����3i�:2�C����>�|�i���4�@�����0(�Q9p�ƇJ�D������^�Y���?d!X�����?�z��.��$n��] ��p�gg����~fMb�{ۆ�騹C���v�":G>���CP�LH�NK�'{��x��#�Ϳ���E��6v�ǻ}�P�+�0����6����?\���ʱ�	�#�=lV	A�b��ӥ���iaS*"⍸�NA��]2��:%_�h@���~��Mo����F���0���?Y�ܾr������da�A��q�_�h���f���*���oN�͆��w^�>Č*\m�������`6�6ugK�DYa1;�Qgb�d����������8a;�C^9��i��8��dWX�!���&8K��Hq9�M���;d�>��d���������h�lLa��G��.��`����U�|�����|�t!��t��DG��|{`����LB�a����% �i��e�k�&�� �=u���^��9��m@�r �, rHz>#+�d-W�8Eϳ�WH�ZF�W����P��4�`���������(���mv �m}��A���?IR|EG$�&��2 ���nF0�|}���������/���>T� �k�c�M��_\l
8kQ<tȀ���n>�P��X��~�|�I�#�Ĉ��]����J@����IrX��-P�/{�b�f�!�_@hi�(z��Ѝ_Qz;���y��^��bǉ#�x��K�S����]5o�i�D�0.|�i�$�c�ei�#�۽��dBH-�"�(��l�,��4F9����sőf�äg��Ј���&Y�3�H�]�G���]x�EZE���ض����c��h�H���D\�b�p��D8^~�=��~b#f����OՈw��U�,�7��9B�}}��L���hKA#�tgK<j�H�ʯa�q#uw�zn��gwf���=j�\�y�^���w�J����������׽탭+���V)�&��m3ѹ�d��<���#]��`C�LK�|C%��D��r��M[�$��|z�Z�~Ү\��ɳxT�M�ŮŦ*�S�!�Y:�c�6��n9�M�J�T囅w�X*rx�x�<�*��?w^�Ǜ���G�-����~�O�Լ�CXݻ��,i�R�` ��U}O&T�Q8��y�@6����ՈuUO:z,���"�b�U=[�V�%���e����^u����2S/�5�����a~'w��V߸�������ǐ*"[�/!L(t�]c/F�aT=������o�D�wr/ns�Ǒ�b,X��ri�E����r��v�e��A��J���G��D=û�����gpP+�,S��\K��^i�Y��5t�<�k����w���y��X�`��el�:6*�>vw%�p&B&u�]��j���ZS����9��|s��h�2�9L��z��}|�4�w޹�z�ZR�z]4��^�����K�{���x����`�z��d��ۅ���S�o�����>�Y�}�R$#{�|L��r����a$���~����,W�"��PH�*���M� Օ{ޚKy���^!�۸�=�N�%Kjq9?D�u�[��ר�ihΣu�/w�->[٠i<�O]~o�2CÙB)�O�5!�Y2�f襬���d����&tm�c0�^��晢`AY�s�U�����ĒI$��I��B�M��+�ʪ�X�\��p��qu�.���:���[Y�0㚖ɓ'�b�vk�.}>Rzp[3�,�X��q�X� ��g��t�R^]�mq�����K�:�iI�i�:��`�e��`�ѹ��V]�'�x���Χ�n�q��K�̝v��Yy�$p�f�ׇ@������mN�ذqpgNl�q
N<��Nw;t�^��6�͎�`AU��0�f[aE����E�1h��af�qG9&��y�ݨ�xN�c<���7)�d�i�r;gJu���h��b��5�1Ѷc %�-���,��*����Y���9Y=[��'-s����󐤈u�h���:�2�/.*���P�-IhWH0؀�-� �-��n&t(��`�b��S	��W`����q��F�\�8�H-�	O/��]�����κ7+�G�}���:;kh�.��iu�@P��ꡤ8)��L�D�����[ז��z�n��[*��孑�NyUpu8N�g�B]�v���+|��+aL��&z1	��:�dP���er��s��*4�t��N�܏�v������^
��FwY�����t(��6�Ǟ}�h#���N�i��å���r���Ci��a0���qn�B�%�C�q����'@����wS�9�*�lӞx3����s�̘^A{��Y��6b��OWZ6��9��k ��A���/c[ٵ�UN��m�8x�<��]u�͈���j�U��`�4Jg64v#2��@ɵ������N�\�;R"d��0{�n��bd��]5�ҵ-�o5@+48z��3��lkm)n�� �N��D�1s�ncl�9�2��͐�͖*;�@4B����ah���Ի�:o(k��X��6q�4�c��t=X6kv�c�u{�Mcuv���qu d�3E� ՙ�l��S��Q���8ɜ�{����z�pD�U��u�d盲.��M��Z�޼�U	t��m�B����B�5�����3��[�ɍ�x����Qt;mH+͓^�|<4��2��B[��Эܹ�V^np���o]=�!oY��Gl���Ok�%��W<���1��uu:�nZ����7s��V����q�j]��1	61	k��utB���F��&q�=�[nM��:�-,�!���=
g���>����;�`����޺&�VX��4un:ͫ�yX��������#E.�9�m�U 04f�退v�����n�`���Ѕ�!*I�p�8k��cL�?r`��2 w�����</�x����Dzc<h>���|�+�����`����g�����]<����&�̆hD���!�#K"Γ﷟,��]G�����Ȓ_J�G!�����6d��G�U����dQ߈d!K�~�dջ�g�f�����I�8���ۺ�Z<�܆H������Y����Ys�+e����̞��_^��H�F�?��js#h��aU����!4|AzDټ�f\,t�;�],4�Ӆ|؁5q��m��p�3�i�ٲ+���C?D!M�(������di�����>����cUd+�_�gE��O:�-�� �|DU:��꭪�Z~�@�F�H���$R/��q�`ed\kM!�D���1C��S.~�js_�Wш� (S9���W�|h���,��Y�ȡ]nt���$��|d��{��e��f� G'�Ӡ	C�x[�	
0`U��H4qs�B9��6�YJJk����C``Fӄ%�S��EI7G�'���cH���a�10b�E�f����V#`A��i�1���(u��}�=� ���5yݱH�����"����"`��LD�ω=:p�XVp���z����7�n~B��`�l��У&�v�����DOH?��"�{����U��m�b�>}Cʷ���x2ٱ/$�b�{�7~~8B8~?s>���в�e$�^���r$㯲�@d!�&t��8V�8��z�<��_���N�3ƕ9�D�4����!�D���i*��g�}�uQ����9
���Q���gr�ҟ�~��v�v��^���|Y�!b�}�ݬ�Pb�H������C!a�2��+��<=#�s�g��lc_f��r��4�[���>�_��BH�Ȩ��/ý[#��n&y���f������m�	q����.m�W/���v��<}�f��3�flMs�qT��h^ӗ9�[��(o<�ē:����gOȢ1	iG"]HVٌ0�f(Y�x�A���n ��U�)p8+j�ꮖ҄c����=E����qݠi,Ai�D>�z%�Θ����m9�oˣ�Q=/|���������gj1!M�T(�X7:ڻ������?I�N�b���ӹg%s�)��k���0&�����r4������0T	�sy5;量b���}�S��k�'�{]��^0��l^�)̓������w6��7��]�_���Q��x�5�R�j��9A�<&yN�ڽ��69��'�d����j���S\立@[VT�QXC�&"�I$�%g{	�"���+E��;IM�U�Q��>sZ��B8AYX��y�˼�1� ��J4�nB-ȳyB��1{�����5ar]t񠉵GI��v�P��f�eY�����n�j��������� D�-܀y�Ǆ�n�荳#�2��O��e��<�uې�r�y���b�%ru��v�0@XB MÎ�ӛ����љ�(mc�|~��,ج6I ���󼮌�.����07�	M��{V�uv���&8�-ɹ5V�F秧4r���Bԉn[�oy�0� �tc�6֏L��\�]��h�4r��:kH$����ƈX=c�����L��pXየ��]�3��_\*���qN���4#Pun�T	}̌�Fgmk�����跛Ź��x�l�#���m8��$n�i���>��g8��D�c)��љ�OK����W�+U~ZlDV�r�Å����g%���P�B�T���쐓7�8���\�������=���kh8�=����� l���l{]ާѝ̓]Bה�"�i�l�,�D�阮�a�U�Xa�g˛;��P�eL�n�>y�侸�����ݓ�Vq��霜H22�y9	 ����ȑ�Wm�Sv�8�˰�!�<�x�b�
9W@��nݎ��K����dv�2�ch6���Uđ���C���tt�EtR�%�6�@�]���=s�;���9͜�*q��J��!����'*I��9�����k$oE��B!Y�Cn��sY�
�ʘd��bl�3%z���Ǡ���珢���>�FF�A�8�F�U~߯ ���"�����?տ<;��,�m_}��͝���g����j���d����$$0-�d�9�o'b��8���c>��P��N`�	h���T�Vn�[�!|0�L�ξ��rf)]��-�o�,b��(!�����Cdm����|/x���D�����oC��1��;��ۡ j��=���.6B��,����c4b;N��g�zm�}�{��n�Ƨ����-˗u5� �M�Vzk&A�@�窠�<����#>��DxMw�[-�)	YX��lт�k^z�LsGK V^������x+�dy�ٓ��!��A�ХŃ��!�)�J�Y��,���h&���\��`�Q�����f #lb�ir�"�����K�Ԗ���F5ٔ�挡ڇmB���ԥv	�Q���nT6��-�l%�+�sƉ�mu�������K'C����S�rs�a��]�9(�n���|���;s��r�x3��녱��{����04f�i��(�d,I �`��&������A��2��b��r�O=}��=�����fh�!�*ސ�\��s2�\5r����2�)E�9 ���Y̱�8����K�TY��.F�����c,I�`d �V
t�Sn_e�Ϸ�|�7��9�D�_�}�$�6Z0@�m��P�#7��L�Svi��?r��Cw	a������Z/;(U�K I�	\fS��U})������	o�&�Q$dX�8t;�Y��� �}��Y�+M[k�y���{ޕ�¯̜�Ş#g&�ڋ#Na_$��[o7����뜊��I�|�!2dr)$��|T�c���/L��ݏYůrn}�\Zz��jk_e\��B��*9@dM��u�2�S�
i�#'.�����ngx.��֜������;3��uҘ���ys�*�J:]�)�n�Av66�|��x}Q���7p�P��o�&�����O���#�:fZt�-��zW5s~�f��"n�gr������F"�[�X 70,�+�n=�cE���x�e�^+�D���K4�2c��2u�t�4�@�35�a��#�wvs�Bq|�@���]ɊO�1�SZD׹N�P6wr�wl��g��f���.�oK�zѢG�YZ<2�z,$�R�l#ܫ�u|U���͂���^����I�� %P>�B�H轺X��Ȗ^dp�����7ax��!mD���
�tE�;Mrƺ4[U�I����p7��b�;	���_=C���NmF@
��|��_J�<a��q��l��٫�E���[���i�0�'�jL��"�����1��ٔ�[�ɀt�|������5Q��:P|]h����gD�� �fz�2�H6�y^�`Wa�-��;��+r��e���2Te������z��]����QxP�h��z�'WwܶA�=�,����Nź��۳��i|�zp���nM���ԎZ#,� ��������h�6"�ha�̧dL@����ۍCj>��9�a+�A�wF�5�Հpp�	��)�|4����rQ� 8�0̊�ՙ����O+��?Z�tK۷����'p��W}O��'31ժ��N3_%�	���7W\⏹�C��ՙ�+1��s���:�#b.�<z���h���/�L�=�u`�"�͞��#4���dc�e`F>�-:�#�o3��=iX�G�͹�a�i�Ghk��>�vWdK��L�3���U�ʪM�@���f�����˞FX0�J`zi!EHۨ��W����@�0����!գ�L�t��1����t/�>ڵ�z]���g���L�e���'����ٿ����D���?�۟~I�\�ι�ģ�C�"[]�]�Y�c�v�+%u��<���͈�-����pc�]���3/.�?�J�c�!7x��\4���yzs���{xyx5;�o��+#���q�289�氆���K�|�wT�]��]	��}QU��j>��C4� ����N����}�k&�t=dWˈ�I�wO$�r�m��(�5��%^���Àf#�U����Whx�f����۬���kjF���Nsܞ�5}�b���.� qȯOo�=c�2dD~��2y�џf��dƛ���]SUm��q�ע��H���ó1�]��c -h�76ٚ:�B+��#p2A˖����(2�؆7��)�CO{ܯ�x����%��x�_)5�!��u伎@nD=����#�6`d�L����!�lo���`�"1�:���E��Go6渄r* �"�o��<���F`5��(�O$B87�fͻ��,e�iq/�����]e��l#�o�R�+u�+f�P�Y.��ԫ��4�:ܕ��j8�rZ��,��>~��#v������DnVZ����;f�o��=�\"�2c�^/U�;����YR�x��b9��'6*�4{=�;��f�����,�]��ӎ�g��/�w Lk{ۜH�:A�������&8�!��(ʑgK�C���A�Gq��W�i�Y%Iˮ��6�(�GF�1q������Sq�霚[TV�l�4h�@�`���-y$�1��n9u�Y֕?wuP��0�^�K��5Y���������D��6h�U����@�'Řy�k4�;�0�8,{����)��j7!��AB�_]���TF���{����<^�Q�8�U�H�$�HC���7��Gȍ@,�뮔��J�pP����w�v��8g���-��M��!�2�Q@�.^☥mO��v?x?ǵn�#�{�͟\�7�����خ�����׺�A|��v�IZkp��a�	5��u����2!`1n�p���=9yX8�넲g�6�	��Ŧ9a�Y��1\�a0m�ܙ�#�����-%
���ZA�e�ˬ�K؅��&Շ��ɮ�v��u��z���W2��9��*��pA�!��L�۶c]b[��X6=��`и�,����m6���lݠ���큒�!).Y�E�)r���Ks簯<�B[jw9"�dt��0�-�ͭݬc�+�"RZ4��Ҁ�������m�6���~O>�L��J���?*Yju%�m���8���f���%|M��M���iؾ�s]�w�����0[�`��A��)93o�B#aY]�}�?a�h�}��Y���`j�dm��~т����J�q�$9��`QkAk-���Ufqw5x�cE �2�2��~�t=-�.P�/&2�:lQx�iy��L�$�Q�S�w��vUGHp�C����!U�y��W��bfD�Ċrw�wmb$�2Ak�??f���<�觟/�-"��_��H����;!�ǘ,a��=4�-�u�0��8�ھɏ��h�����T��/̲�Q'PANL�<��V�<��k�[�f�ڭ͎o����յT��zP˨�}��G�v�����:��P��un�R!�:L�m6��=��f�Y�ő����SKܮ]�lb)���j�2�:Ƒ�ݗz��}}n]{�0_yV�Rבw�����kvc�>��B	vH1�B�	��s�|�#����`�)�*F��+O��HWTt�<�!t�!q�'�!{�0�W���ŕT^XW��<�}�Z�8�˕d��赝���gL^��P�����z�9ۣ��y�W�ӷ�����_D��jߘ��������`c��+oX�����9��������y�"�p���M>@aq�-�W���iȆ>���Ȭ��@��`L_Z��ܗS�e���z���]WJp#�²��ZPt�2�r8���*�4I��r�)�0 ����sʺh�3�L� ��__bspg��Hއ�L�0���x�9�c�	�,���[g�4T0т��pQ�v�y�܊n�Q���ޙ AM���ǽ9d
#���@�lг���6/�v��b��F�$ �:G���[�-��-t��C�	.٦�uw'a�V*v�5�0WMf�%���L7*���.��ӳ氌��u� �4��.FƝʍw�5c���W����,�Vt���gy����t4���>O.����C�I`9_;��FF��_w[�Cv�a`��/��"�������\C�a�'�ލ�{Z�s<��.���,ح�;��4i ��:�) p)#�<9�>���Sk��:�}z��m�m��m���N�wU�;ՠ5�'9����������ޛ�8lK�j���*���۳K.E�V�T0�T�8���c$ ��W��B^��Nr�{�eAw���2>�/Y��%%sU��v����ݧ�Ҧ1b6ħu>M��q����� �=��+=���9]���c��^�{�i�8��'�Mz�C������׷�Ќ��e]�W�=�gA�%�V��-m2��za�����zzY֬i���zw�i������?ޣf緃�������+�{��݃�~����y���@��q�5yw���[�\y�jde,.G�>�s��6;�*�^{N�Ɣ��f.��8�N}L���G�������n&��9���?Q�M����! ��0�u�=���މT��F�F�j1�8"/f�fp��Z'�����QӨg~��ݣ|�Ͳ����.�H��̫����w^Gct��y9!C��r�X&��Vl�vC�����X�'��l+0�ky�]�> gZ�z̭��ɺޗ2Y:���7��h�q�x)��J�<�
������MF7Gd�b�&2���tr���E��'Dދ����e?��M�d��y���X	����I��b�n\���}g����`^����R��<�s�<�6=�����n�]�:�9���R!�3{�8�Cs�(�3���l�+�/l�N����ު�����/$��(x^Nr'��������{��/���:{�D���Mޫ\(�D�_�ӸG���uC�_�����{wF
�H��ߵ�ݦ&0��kv7������oy��:F:Uů}���y��R��!N��H$&��N+��`�ԀZ��0.Yތ��i t�tߟ�eо#��)��e��#���~�d�ő�5y=�����ۃ
��i.��/��q0ԋ��i�.ac3�Ӂ��;�2��pI��^˩��f��?@���aM�+N�/IH�	����OM!k��*:���~߿K�#H��]cK���Ѵ׬<��C��b{=�|�BF�+��Ƴ;f��=\e�rbBډ�y�z1���q��6��:FOh���ֺ͏۾Ս�l����]������1�>�����@d��O/}y������B�Hj-��/��YH`�3�Y[כ��L�;jhQ| 03��E�5�V®�s�^�jj�Q�}hq��,P�Fo/��@�G��B�D6�(�:w��<Y�3��։���o�X#���9A�:j��0��xC$;�V�i֚6�;���\U��t�y�f"�A*h@�(�3x#����,K��@2�{�0ߎr�.¢��;+�.����i�t�cY�T9ك^:v	Ni_?��<}�S}{f��Z.��2�Fݪ
��ćO��0�mZ�Q�v�aӨzo��[�0�();/6���<T�N,q�[��r��0�L�HpȉNN�1�5e�_<oZ�d	���{���`&V��M�SΆ2��f�׼sEﶘf��?\vY�b	���.�mPg�4��~�nB�	OZ�t�U�-���<�q�A�l�:��׬J)g8A�١pųCi�)Fbc�?8
"��q�Ş�/y��9����UBƫh\����;U���1��/n�����˳5ޙk7q;�2DڑX��Z�_7��kraB{ǚ3N��a��^pw:��[�����+�0�E�7;�xx:�N��!?g���NaBwMW+��� 0�h{�:��" �ei���|��q�C%!}�Q��[�CC_Q��CWX�2��[����F�hig{�8i�6hi��{�Pƌp��Q�NRs�0Mz�:rm\o�;/���E��H�[���qa�y�������M6E�뎺B#��d��{9��!�X��]�P`k���\h�Q��;�,#�H���\#�"���>z!L�M�n�xX�$㬔��H�Xǽ3��B1P�ҍ���sӀo#�5��,	q���a��H�x�h��;=�`���QRn�u	l#���l���zy���R�8�"eBZ;Zm�R�����v��ϰ�ڽv�'s�5fA��ޤ�B�q�1<б'+�9�����Nٚ��5�m�s.��8!�p]��k��Q) ����F��c�F�6���Yut��a�b8H�k�R�5]\�%�f�d|��c4 vm:��ŀ�f!H\����D�A-��	����69<��{Sׂ�wm�<vN�fn�g=�s���m΃-f�}����v�a�F3a�R�,�KF	����RŖS9�jV���nL0>�]ټCe뭟q�N�%x�;15�MMX£���Mm@�9��V��� [������\��{;d��L�/��-)\��ٮ��\,U��~ԒLxCE��(05di�7��O\�4���o�50�i�CHtE����P��>�y5*{h�B��NP�{��\�
��*ں
�`�"�m4\M�$���k�Oeq��Kۗ��O	YT�EȺ��� Y��Ǆ�v��_"hf�*��0�}#�x�J�y3Bu���Ք�{�2�F8d	��i �F�����c)�9��;���<"��}�u2�X�li�ɜ J�����묖X���Y&��&�޽���4�*cM1Da��VF��q��NGc�e�0H;;��cyCфGJ�;���"gz^��#�ȴ�t��3�w�P����?g��:�\����j����>D�_b�8�mu� o(�5���v�r�o�����6"��Kݫ�.n�J����_��t�6�.fO��k*#�����Oʶ*=5K�0r��ws9wV,���'����Ҹu�7F�V*���,�V �6մ�1Q��=�:����?Յ0Py=�_na��7ĩ���V�㏷!F���ή>�FZ.-y����s������(Yy���Ƚl�������Ù�7�k'_;h� «���X�C7���`ap�@�����7�^]+��c�k�o0t>_�i�px��n�P�G�jr c1FNC�H�U��CC/�v4՚�!���U����:�Y��)���#�^� #H�uP���#��t����T��@Y�q�8abTI���"k�o}��Q	/X5bg���	j�Yj����a���!�_�|����Y�i��uӠ٠�%�Ԝ����k84�8@�sܿ p��DEq���|k�Uu� ye��_�Y�����qM�!��ϙ,`�a�u���Oէ�?!� 	����8������t����]W�!���A�)	�R$Z����e�L�u��%�p�f[b�.��9l�8#֭]v����ϴ���HI���7�2,��]��K���N�!��5 �6+�{w/���.u������m�!�H��?a��aI�Q"ʎ�
I3O	$�F��a��z���i�������#2�|0ia����#MYd��i����K�E���!
8@������Z�@�Y�)t�"Q�X�2��J9E�q$Ͱ1���-U��_�tX�pt8V�i���*�s/�n2B����!8;a�z��:<���.h��W���C�pY��ik,��1|$�F��S�T��Ef��FI�8&��N�{bL>D����;�����\`/_0غ p�UhW�����tj�H�i&!r6��	�,��;�[Y�|�PU���`4������`���ج��������d}��NeT�L�F&!�O����Κ���Zj��4��i{�q��Q�q�N��
Ȯ4N u�N� �! t� ���_|��I�b����X&�������縮�4����2��`��������ğ�|����SʀH6�])E���a�g-�Rk!���Х�83�fŦ��љ0�9#��0�[T�@N�!i<y�K�!� Mj�}�:9YZJ�uA Y�(0;�.���G��ғ(r�:D��`��m�L��xн��ar��0�#EĄ��\�ls���"��{�<��>f"�H���~���.��]Q�Os��x�u�0Mku���úV����z�#f��[6��7U�A�=e��}d$R.ԆMs��ElV^�� B<�Dj�?@Λɦ����n��&����h���һy�wj�ha��D�[�{���YCM ����9aU��)��N9%�À���̨k�Wۜ����T��,Q屢${X��5�����yTw 4ի�[=$��צg �SE)y"V���{3ǣI#W
�i�|$KF!,�,6q�k��"6{��z��|�[�p�������Gd��!p�㡥�t��c���ZR%h�&V�9D⽑WĹ�5�>�������_{y=��e:��P@���1�����.��X�Zu��@��p߶��Hs�t텤b�#����8�JTLb,�Qkq![Y��1�;1:�!a� �ڬ�cM[�ci`�Td���r����(k�@&�0g'�  ~d0C� b�H`�V}!�g�zZ�7x}[^#�Z@i
��R�曾A!V!Z]�A Mf_�L�gԌN8qen
� �ȂE���_n����(�/�ֈ��X�~�2��,��YM, k#賂Wy(:�Kw�/�j>��:�|�#'8� � k�`�V쨀�R|�����v���u�}��7�0��R�U�8l����7dX��7�8;�M��G�����M\.���V�R}"���uU�M� fz:�t�5a B�Ҫ'zÆ�(��R��pCV��&�VG�{�)`�/��.��"�� *�a�{�� ��4�$��@{��,:�5yt�i�ɡu:���m�hg��QU�����<'� ��fHn��a@�� Y\U�o�]��@����,��D	�r�v�,S�r 0ԪѮ��t޾i���t�J�s����]r���X����M��m��=T�|C���ZFjg�:wm)�n��!e|���g`-P������+�����{�4	�)˴/�x��=e!��;#Q
T�m��n��A�9ؒΎ:�K�V<%r�V�����9�M	���Fk��!��)yQ��y�{Yk�tɐ���Ԝ��
�"��{v�Ï;]r�	nDv�Z�o�#<��T6�[L�N5��R�7it/B�n@��c�yܝ@��撦�gkK�B�s���l4`s�3@֙RZX�Ir�G0����tU3���&6�F��n�+oNy�L�l�X�O���M��=6v�Gn�n��Y��H"Z�pJ�D�&`������Ѯ���|��MJ�!���M������!�4۪@��ӕ��z�*��x�B�*��o(`�i�5*��)�,���|�w����=��{G��l������V7<�|�  %P�LQ������a�]9�*���0 t�9�	zh,�c��L�l H�CM撑�����4Ђ�
��<h#J���`0���"�I2�MI�2V�A4k�� �*�o|lV�(29��pԠo����t*��٧��h6���!�8�����}��4��*$H�]����+M �2V�eB��@ M��ZC�$d�an"�+HZW ���
��4�ՄOrƑV,�ǽ=C�	�"�t� 0G����A}�U�TGO�MU����P5�h��K��ɷc�2jz_��&��
��+��"(� y���<,�l��LB�QǕZk�����@Y���s���45\! M"���0N�>�� �嫬�GU!�MMt��F�����H �Xi�4�,����U�4�J��P@i����ܚ2$6�2Ia	����۳��K�gP��cn?�e����;]	R���[����oΞ���N�O�z�)�L�X�<�A&��UCP�;*� _,�t��C�@ ��=��sBm{j�Wpx���!�C
֑Y{���T1Up��^48h�'��CA�E#��J)(i�u#XzX�����S�_.��p�DsٳW8v`�����U�F(&)�z�^D�E"�b�u2�D��b�3C�۲�QJ�0�|�;1eb-�.#�3��J���C���`e����	5��V�A�y�M�(��4Q�a���C���_	�����,�v�dȰ	�p�+��8!��X! �'�p��#�T9tӫ"��=����9ThY
�P�!�������N�PE>���r*[t���_:leZhY�(����C�g��(�) 	�(p�b�.�������hy8(��$�U�s ��j�r��xƉ8��D{p��J�"d���0H���K `��0�tHM}4��	�<`�h[F�� z�� ֆ�s7��	 ��T�}�t8E� �y�0��M�*$ے]�[b�<J�5�U��h�oۆ�i��"��5�0��4��6���<8�i��@iؤ%��E��	 �\.��5Zk���(?Na@ pЯ4h V��5�����y���:{=i3��L���LP=��rQ�i�9�[��hǤܽ��]���lf�R)ID�LȌ�ei�a��hC�z��t4� �j���dB�C`�3��`�y��A^(�����D��.����Ĭ�Rm�Э"ɫ4�4 ��N{����HB��K�����Y<=��r�s�ʫ��i�("l��K �iPI���pwz�WWX��� pP� �L+�ۆ� j*�p�C������D�:@�t"��CMS ����<l�@ M�`'��4W��VCJ���lT��S���
8�W	�"�DuAP@@���_��4�F�Eset�dd�I�9�+������[�;6��ۨO��S�9�"v�X;B��*nP��zomb��Ԣq�&�8yI~�����\tyk���rZ�FjJF{���������K��8E.���8Et�@� I�\F��}f:l�L
��TH�F���*�I��#pPT,����x�������I����b��Ea�U���4���b�UU��ĉ6@�	�F�W���X(� �x��8lQ��v�"CH�-�@����L
5\4�*��L@�5d��h�p�2���pȑl8�CMwh#�������D#�w�`��@a����=�F�|�:D�x`�S �@@�P�� ���:‐M�C�h �F������ ��+� �B���i��t�1�����c��?%J�>�%1�Q�G+��	���3q�9�RbL�mG9����V�X��Fc��Zk � V�&��@A&����uCH�@�a�#d!����5W�,
q5
El�"�� e� �I5]�睊�N���+O�"�FP$db��.�АB*]޻�F�UZj�F�Zie�"8� 9=�̥��1�3U�I�T5�H@Y�+����M�w�82��(*骡d  �g%��;�("��49 ���꬐hiV{ �:j�$
&�
�{��H&��� ��9
�0��0�T4���|����v=z�+�#��-�L�E+���
�C@*&����]P�8*Ъ�@:��(a��
��u��R�:hd��6T�o��}@i�!�I �MP�����5B����f�"�H
��pЯ=�Y�5@�CH�� �x�V2P�`p�R ��O�(H"&��T4�����ӹ����#E;��}��7��n
aM � �V�$W}��b�C��j�W��@�������� J&���:�T4�KZ��X������O?I���y�.���j݋'��,Au_EL�U���m�IV��ڽ��j��F�^^��[�:{��Ԯ/i����M�������~����~ ��V�U��]:D�I�4)h���c����L9Gy$�/w��'��:�M
�A @���`i� H&���� �ZE e��_�Ш<�k��U`�� ��� ��ˡ��V� a��@�5H	@���7d�5U�B�&�4p��9)E 
�>��I��:'�8+E�(�ȅd�J8�뵱�����M���B:�˦�s(@1),j�fl��%iX�h6eU�:t�d�,�(�E�
�T��\~��@p�)D��ֈ �4(aв���y�
4	<"� �5�
j�&�"�}���@�r�v��Up�� ��� #��T{�E��5@�B�@�D5� :i��0�PD�����7G�|����Y:O`im��E �{���4�x��j*��
�C
� I���� ���B j��*�:�"���xlQ0�+HVh:$4� � �᪡�{��PEP���Є�=j�uU]5L� ���Ǎ�zpC
�ӊꫦ���a�KUU��DU~� 5X1#T"�" �Uf��E
���� PZ��5Uǉ�� ���A��4 o�n�x�@��BȪf�� ���
�Ol����"�Ea��4�T�^�)�B� P᪡�*�*���90uX`�*��T=%�*��5B��� CUT����P:j�CH�*� (d��]CH U�T+MU#��J�����@{���P�T*�TW�� W�wo}�tM@�ŞwwOvN�gI��
�@T  8E
��xn�
�UT��MPf����0������P	f�X�MV�C� *�P��x` i�8@��  ]�9�>N_¨ UUЪ UU_�T( UUaT ���� UU_Ȫ UU_�
 UU_�*� UUW�*� UUW�P� UU��� UUj ����T ���*� UUR@ *��*�  ����U  ����U  ����U  ����  �����@ *���
� UU�T �����d�MeƒLC�f�A@��̟\�z|���T�6b��d��))II%�*�g`9P��)���B�)U� R�"T��BB QTUU*�@�U%*��                                      �       } q��e��=]�&�<�]7���Ӥ��Wx��lO/ y^�7wX�x�W�<�v��ݼosD�A�4Z�x =�l���ŧ����ɯ���A@Sn   �    @� �    =�� �r���{]��v�y�/a�^�z.��z�^6�SJk^< =��c�]�v(�ݷy��G���0�Qw��o��@2�] $h�         \�lh�k\�G�����j��{r��.����&�F��Ov�� �96�-����d�em�nح���&�-�� ��۔��3�^���7u��@5ݻm�<=�6�o-쥷�.o ���wmu���z��*�7v�W���x��l9x��g�]� 杚�W.Nkz;��9�MZ�l��޺�^N�m��2�@���        �T�ۗ.j�5�.��̴�R�,l��]7 ��f֜]�Km�c�e=��\��u�㚗i� w[T��e:jK�9M��ZruJ��r9� h�fڹu��.G�TRn;��mm�;.ZKp ˑ.]p��W-�m�s�WMD�Z���M�+T	7         n�J��i�[��$T�YPumNn�j��� �K#.Z�%4����i�r�e.Zu��� ��I�pw�J�9�v�Q�`R�R�uʚm��d�Y�� s:8�.�����Y���-*��9��Zp ��i�Z������l���.���6{����l`P4��p         v�h+�\#)Z�:/x�Gmyw4J������m�<x sֶ�j�<vu�d����ׇ �Z���{[N�nr)B�7� �Uz��..��4QG�o{p����ij)��yqUOko7G���c�� �+�6u{�E�.�=���Ǎ�e��T\�skL���� {/Zmf�,u�:$]������6���kOM;x�v�ж[/�����M   �~�R��  4U$���F����R�E&� ��~MR�  ���D���F# ��߿����_ڪ��/��p�no5G:-(Z�Bn,VZ"��b�tξw�Ν?��� �\3��������-*���R�j�H0Q
"����O��Tc��S�ʚ���[��j����DF�ֆ�v	���ނ��7-c8h�U�'/H�q��C��iR[�d�x5B�Pf7%5�Be]˺h)�k#.�ÃfJm�K�nf�R�r�{���Ӭòd�*ӫt򴈲!g^����ð �3k.�B�����"��[�[b������QF����::uU�7nRZ�!&��FDl����tQ5��%cf�zN^���U����i���QB��j24e���Ef�cr�v�͘��;��Gct,j+f��L�q̓i��Yv��f��L"eX[��_٘]�6o�x �κCe�A2a�5WY!й�[�v�ȁ��õ�W1vXn�ǈ�kM���h�GJ��Z�n�8�4��,[��M/:.T9h�n�2�]4���J��t�;�0�HIb����9
t9e�
�����U�,'g�8�v��/ul�%�o)8�ɳr�-�V|�������Ů!J\�pfw{aST!D�j�Ā��P=�����3]�����GoS
Vd��ea�&ةslJ�R��-U-���kH5u*f��(#��#`��^�,�I*f�xn(�qe!n�ȝVm����)�9	�1�u=KoM�֢"�R���R�voEVk�Z�iu_�V[7-���lر5,^Ǧ�E�Š]�ɧDU.Jǿ\�A�>�gL�n��>eIb�R�֫y�y�Сv)'FQ�&n���;/"���u_PN��t���x|d�*�`��U�f5���Ŧ�^n+;�m��E������A�ՐC�hŢ�-*�)��!Xt,S�;JQ�xH���3Yrȯ�������1B�H��<Ũ�Yӻco>�dKj�K,^Q��j�i����5`�Ҽp���ov�ϓf,L�6��5�ռ�ߵPa`u2����E[S�m��s,haA85nV�֋+��mL� Ҡ�����PO1AYXpݦ�`[���n<��j+M�Ւ�#6��;lV�ܼ`����E F'$2]c֍
�J��z�/�bX�ͨ�k"��8�ޅ��P���'�������q����n5j������e��&�Wb�*�e�btI�0�L0�6��ǳ>ʷ���@f�X�Vn-h��T�VE5i�.�-���<��e*�����L�p,8��c:�;Ү�P_e*4�	�&NK�'a�IzsA9[�e�Q��o�Z@�櫢"o.2��NV�ő��k��!RUsm[��B����m�q}��XT2h5����U���s/XӏZݡrP�蕏/l��������i��E�6�g���$7qS�"LGaZ�	C*`�n��R�^�3C�2�n*����{�x�MĬ�%d0f<f5W�Ft��wm�Ú˼WYz���d,�����v�KN�]����hڲwŚ�Q- ������tHB�wR�Cu���/720����T�r}iGuY,٨��I-���v�F#{�L�CY����2���ӽ��xL��-��%nI�ڡ
���Uf�n�	&�c{�P+%,�n-(�z��ܻ�H��A���ɑCE��)zvMj�Rԇ��C+.��V-Z
�S-[Z�/4Xܭ���b�P���֮�sm�2��C y�/'O>�%�]3�\��.g~�㘫�i�45�ׁ�(ܕ4,�f9d����!v�Ĳ�K�6��$ِ�t'�R�$̡j`:f!V�&��wl;�!�4٬��.	�QY ý�ڙ.��8�+���ËB�m��Yh��(�4� ���֛ϭ��2��6��s�b�h��Z q�rʬ�LR[kb��2�DЃ Fc�e��������0�piK �k3Eݫ9�EVq]�Z�L�T�)z�ۡN�Nf�3u�)hR	;
2p��3[�Iݣ���'*��������k1�s������v`C/��yw&����QR��
 �P�P��Y6>J��Ě�4Q�*"��oo�q)#D_h�t-"��	��,Ŕ(F������Q�U)B�!%���i*5^r�9$@�'��v����iu���B̾�*�@���[j������$;�"�vQ��g�e�w�u�h�\�^��n2X��N�K�n����n��޴��Jh��ɠ�e���6X9�6�l�A��e����mc�adٸ�55��hؖ�W���K�x�����ٸ��bv�D�д��Ya�9�#�Y.�LF�6f�P�)�8�APj�Ҫ�n!���[�I4g��ٔ��F�1�K� Ʃpq��L�'��%����ڇ	�@�:��UB����h-�z0L2�I�)�2#�n���h<�,���l�Z�jL��� ������j��l
���d4�%t�cO%٢�YZ�;�2��P�-�����'I�KUK��6B��2�#s�
B�0��jӗ�V�����.ҭ�wM�v���T0<ۏ,9	?:��,�ݖ���
���
�K[*�˦%��Mq��N3�������@Уe�Z"��mh�GD�(��T3h谊Y,n�{�Q`�Yt�a�D�.h5�4\��HQ���
�N��h�L��r�TwJ�4��d�nDv�])����ս��6���PvB���=���o7Y{#���
�*�l�2�^�(;�����,���q���&_q�qm���~WyV��A�[��bEۙ�:bVܘ�J-E�x)��K��/l��J��y7ꤞ�c��2⯪������n^T�ViV*���#8�Y8흦�p.(ʛ�^�,5z^*bSŭ #�wC�.k�B�ك̼zGk��-]s ���u�^�B��轍�d-b�3j��o5lڼ�+ ��('-�*�k7�yL�*mj�6M�܁A���/M��Mɸ�Nc��U�̹�c�^��)3�	��ץ	�6�ǻ{*9��Zq�1�c��]���۹��6�u�kK��Ɉ^����n���;g��VfJW�8�T9��,m���kh�jֈj���hT�=Ԃ̖qU1oW%E%ޥbC71!5:�LL��χٖm ���Cj�IԦN;�����6��J����Ov�!X�D�r�6��H=����Bdg+^m�CYC%��*��8
R;N���\e��	����>���m필٢�&A�{���ڦ�����L�A�a醵�a�2���B��;��	�F<X-��f��c]�4�UE�Ҽ�G�Y{��_ƚ��.��QD�D��ǟ5�eJۖ4Ά��+-$����r�k�iOI��Q��BV���^c�L�O�T\:�,U�q�&쎜 ��TV�\Q��=����:�q�Q������U��Y8�45
mFoJ�հ)ɘ���
�!SZ/q�i��(�2�j4P���jE����լ(�tU��,�&M3v^�f(Z�oqh��<������3���f����1�����B�ֆ`$�������,ؐ���y� ϑƔ��b�wH�ܿ�<#QXљ��p��Ղ#���)����F7�[N��,KZA�vJ��t�9M�є'���5�=��PBM֩���˻5&A���zF��k�C{��%�7m�����nFfU�0d�\ � yr-�i�U�	�K�BwHZ~/p	�/2�,fbٹ��/�"��iӘ��u+*EP��`n^��&7z��͐̈́��
Դ�2���i$elW��3-+�&� �ӂn%7Y��F�Ʋ�Id+K��4���\ʴ$��*FA�u�
��ơ`�w��d<±R�u�e�PdU�i��M�����F����ur5��3�`�c拏xE�h�U���S�]�;	�หi-��kqB�QDQǸ��"�lf����n�v�0h�(З#YCVcÚ�
ۡmZ.�B�����J��� Km*a�j`v�Z&�5k
�Z2.��FFS���7k=V"n��5c0[��[$�&�z��M���0L=�4j����M�h#@���Z0���J%X���R�i�A�vQ;4(�DY6@�U����KE�b��;J����e�NP�*��񤊥{Z���V8�Q������o�X·���]���Ðm)�Q�0���Y����ԡ�km��ʼ�3�n�vXzt�t�z�P楙�0�.wܫw;�>g^S�@�Ohd�k]$�W�-PLeT�~Y
��Ӛ�٫z~߯�Ya����~�h1�k,�.T�#϶��OҐd�&*a��È��R6�2�\��.�
�2��4��Ҥ��-
�CC6l�����	tSԈ"��͌��M1�gƥ@�n�B�I^��XNLIA�V���D/���/mA��^b�Y�h �bZ��ܻ�b͛�p=yf�E�:��f�[0����x�`�V�8w1��/`F���a��m�D͘�~�ּъd��I9bSZC�39p����4�AgaYn��al�m�i@���yZ��;����:eKQ=yF�-I*�^������M��7-����]�F��� uGHMZ!L�AqT�%�[�5��t�R�Y*��@���G�r����RE����7���h��G-K�m}�i�cE*���RY��GS&T̀���x�ҼXM]�"��:�z�!Mu>Y��۟0�ݖ�c��u���
26�˂�e�!ٸ�ba�Ѻ�1Ǉ99"�Ka�w��GxI7UޫC
���
�+�
��V��Ԋ��Vp����ChYz�P�������5�nB�ſ�,61F M���r�:���C5�w�p+Wj���)�D]Ց��,�ѵ��w�d56��%7ݥ�]7���f�d���cJ"���Q���4����D8���%���d�4�Z���b#i�0�*��TЮ��Z�J�4�J���ʸ�y�jf�*��fЉ�.^�J�݌�Fn��+gb9Z��2��Q�W�p��zF��������v5�,��5@x#���Z�u,�Sdu70U�C�������ٰB���46�/�B+l5l�-�*je�h�;4,+j��c2�b���Քqm"1�/iT�����m��ڇp+a�j�ʸ�v�5�l*�h�u�
*�D¦�Ԩѕx��̸�)�5��p6b5�.�����:��kZ���:6�,Q,�P6j*�Tki��Uc�4C���k+*dA�`�gE��FN���ۭ���QxWo`���Z�x���Q��,�hX#�w��2ӗ�S[QQ#d�9���nˣ����2nM�E-���ߡT�n[d�N7x���T�RY�J��TWX�T���\�VĠ�F�N�'a"L)Ïo(ۃ2�8�D��֚M��C�(�@��:c+n���W�q�/�F�R������8μli�sk����#�S��-U6�nݜт��D�3���X$�ˋ*�BKwA;�����Wp!@�(�T�p�=�ϳ
&2��hd�h@R6o6CC2����jP�:S��J�
�V�E���͉b2�{ի��"���a�,*\���x+h��+"n��8��d�����2�c܇j�5�eI0�˚��f{��n���R�;���xƩ������@6��՗�f)D�v΅DL,-Ku�(���H�?]��sۼ�26P}��jL�z�^*���Ä]w֫U[W�V��T�#x�Rl��1�Si��|�$�V���x�8ݼU���|uKm�_jv�e��H9��ܔ��9�҆J��Rb6�D��:�3^��m�4b�&�-ə�pHQ��&J�U�ʩUN,�%A��N�eR��!��n��7YZ���r�t�`E[�w�Ŗ�%n6��,��(k���en\�Z\7�D��v�t��kn����,*JA[Z���ֈDd�"w�Ulu�]�)ѐU6����ֳRt�0Ӫ7V�6�m�rAg2᧳5�9�5�n����|��'� ����G7Iڽ*����2����"ˎ��w�Q����c`(^@f��HXH�Vu2J[��I�%�׭�ctC��*(�0�N���GӁL�y�V"B���I�RY�h�l6��kZ��C�3�4h@�+��oˎ�bW��uM�W�n[��wJ��Q���\�G �4�ШiB��R�<���V51	3:B�()Cc��aAU�ʅ�%��ψ�@[��xu⦅M£
J^�r8$�ZGv��t�`ܹ�h�PK������wb��Q͸�GW���P��̥�-j����4�����p�nӋ�vC�܃$U��4#X���Ce}yl��/.��YV44�����{����r���;�%�m;YZ���X�^T:�fh{W�,�P:��z.�h�*TBa���V��Ji�	�Äm�=Z���X���b�b�Jad�.:�/�������134���*��G��/KċͫͶ
�d1D�q��;�Z�v�f���Tl���P�������K�۪���fV�K5��ⱪ���VP[�mF^4��[��l;����oP9j�']JG ���Ů������O5l{$�bSr�����j��s%��\��v���	��InMY"*j�r�c�i^�3J�Z]���ktf@F+ea^�,l5�����Ʒ.TB�A�JƲVϱ�#����Ȉi^�M+�{�1�n]��ճdbt�B����1^�aX�uh�i�R���Τ*��nb���sf5�C��'%'�+v�;��d�eû�@��nƃ�ۖ*i��$u�c'ٔE�9�-�:�r���i�h����� ���QS+�z$$蓦/���Sv��V\�����2���L�p�¨D+V�-��^ѹ>]�Q2I$�FےI$�K������U�V8*���JHī*�UUUUUUTUUUUUUUUUR�U6vv-���j����j��������N�����Z��j����ڜh����U����Z�����������g,�j��������������������������������������������������Z�UUUUUUUUUUUUR�Jʪ�<�]��!vPv<Y�|�޺f���U0z��3�m��4;��7T)u���e��.ܩ�t�6�&g�ݛ4.M���P�شu�0��qڴ�zW6�s�]�^��>ӓ�u�I͜��}�e��j���e���c���Dc���mn�q�ge�'�NG9۠b�9x�vF[U��.;7v)N�������nʑ�����T$k�l��]t��V�b�^�{<��]�u�=�筢ц���+����6�XN��c��3ks�=�U����J@�Σ�vA֍a�Gq�=z��e�fl�=�����5pm���k�.ܝiuݶd�.l�:Ý����Y��g;X��L�f�;vWA�'��ۍ���6�]i0�7�:x�c��퍽oU�M��qՐ88��4�g�[`��@�K;��\s�<v>m��Gٙ�T��������B����;M��h�8������V�8��f��-���Gm�/<q\�T�f�z<��h����̯h�6�ܧg�L�˭��\G[Gml������n�4���\b2�9�8�n�w��w.�h�opgU�m�&�nw'b9*t��玢��k�{`{gvlW��s'�؃;��Vf�ƃtp�3��g���5[�K�=qݜ.�v {
]���/F�y.9yO\���Vd��]�)gc�Ʃ�6��v�)s�cy\�zY��n�	��E<uQ��j�{n���i�@�+���^]ƹNڞ���K��������s�MR��]M���S���L�Eݍ�h����Dn,�܃�ݰ��6��γ1Κ�����Q�/@��6X��<y�Ʈ#u�8z휗;�	�;a��gwi "��;��;/]�����-���0��D�m�y!�r���'�ݏ3�m�� ���^��v%�̽^�f9{v��>C�c:;r����p:hwo������ջ����\���G���m��Cڼt��M��@@�sx���>'a�[��uGBsqۃ�||5���3��u�l���C�q�xݸ1���ñ�7��g���Lo=gֺo���]���&ڰK����%�[s���p��"'Wu�r����3N ���v��e�JL���k�
g�Ok��:g�#;��i�����o?Tv��v�9:��q����i�|���7=��;q�Ѫ'7\�v��Gi�盷k8{pp*Qpm��>�ü�r�r0c��0�s�(^E����WmuKv��=��`�u�u�W�67�7m�=�ú�|���mۭ��S�^�%;I�g��p��$�l��7'.��1l:OA�m\N���p�N�W=7D�9��<�dǇ�`�ސ���#�ϏG3�yݩ��{,qӵ����M���Vm��[s���m=ڙ�ڎՉ|
�6��&w��Ӻ�G�m�7���x�N�{Oc�{DZvе��c���]��=����n�s����J����}������x��t\�s�\��|l��nH6�[v2�q��m�ڻ���ȱ��ڻ��7�Z�Kn.� ��ݳKj�:n����^�;
Ql�ܨ�{y}q�7]����
�']�;���n.mo>���60�K=����V5����w`�tlh�N��ݸQ��{���]��t��q�vO-�t��tNM]�P�1�W���spj�k���Z5v:k�T�q��n]sQ�m�ûl�����+�ٵ���Ճm�3c]2��m����X:F磛r��U�66�s�j'#S��2V�$�D�Z;s&�`�v�8�x�k�<��=mX���Dٺ�����s�O[����'Vx���[YlX�<����gv1m��h.�]�c>�cd�vf��v�7�ujH\N��n�b��	۫n(�ml׫����+1B���$�Ϙ�60=nOu���ҋ�|�ݝ�7�n^�2g���a�n���*��'9��qn���'<� ��2 Z댍�Ӯq��nr��n^,�q�:�׌p��7��r3\M���vG���+8�a�(8���'�B.۷i���+����+{O7Z|q�v��c��˷+Pg���K�V펠����a^M�{rhxɞ.��z�7N�ፆk#�ge��n��u'�3wT��5�`�
�k� n��>�m�&�x0��g��cn�z��^�H0����c����<�Z|z瞵v��9�&�2Z��'m�=����W^��	�����^�)%�u�(������\z����s�
�Me
�=�A�絰���nq�:ہ�9����c��r�[�����u�[oU�oi��rc���h',v�۔=�wl��ևTgZ.��v��RE�
!U�G>��{|wI�>�q�t�h���������8\�}���̆�G��2r\(�3��tz4&;���pB�76���:�{'�Q�Rw9�����V��@�u����^p�\+��zFxhj����p���:-FC�x7��}<`cvKu1��ƻG6x��vSc��{��:��>�uϴY�`�m�"[��eݷ	bv�p'Rj��9�����6v����ݺ��W^�N��<��4�7-7euR�u�1���W���^>�E�+Q�q�ё:K� ��+ruY��a�-sk.3�Z΄#���mݷn�J�m�웷P�M����T���k���p��Ě�z�t�W�6���tv"�Qs��;'\�d{���w��c7ͷ��=�Y�n!s�ivN�kss�犤�ۯi�ܼ<����[h����jxٮ�3W�g��λb�:�^�m%��㍀q�����W2�5���9;�����N�]��M�q�'����J�.7�Is�,�9}/\v6��n���Fn�����[ַ:M׬��;����]v�m� �a��P[q���nq��ٵ]mn�ѹGp�="�AN�=3���hy7��i�8�n�0��,:fn$]i����td�����wuĜv1�q�N�*p���6s�%�\v���Y����]�b�;���]�0�m�+��n��S�n�Nm�n§o]0�!�n݇S`B��kn��@�9�>r�������=�Q��=\*�l[-ڑ7�wh��!��[.$�g��!>��6ݟv�g7��C��V��8�]��b�b,;]\�2���v��ӆy���{C��Lx�j"�7<�ON�չݸ^8��nx�ø7lw��Gu�%q;<!����<�n�a:z'u�u���}��鮵wK�������� γq\�g{vks%�<r����ֶ:Y�u�ɺ=�u���r=�sU���Ӭ�g)�p��{n�
�pvx�	���
�5�m��櫞�^:��꜆���&��lnƱC�lw����{�ź������t~�>��]��dd1�)��=]c;f�S�n9:ފܜG�4xu�ZK��:�/�խ�˸�G#l��Gm�Y��
҉��,�6�t��vy�m�; X�-u��<���>܊�2)�l;��b�<��n�9%�tU�&�A�e2��Ǔ����Cl)֗��m���Wm8x�:��:J�>7[�X̃�ю7	p<��Nr�������鵄�mA��C]����O@�y�Ki�Ӷ�t���q��M��W;���WY�'+��d�!q��4�;/�pG	�����]{4uǅ*c9�}v���^�	>p��ZѬ�t���M&N�Qg�;�u�1��ۮ1�ӵ��C����*8t�Q�q�^����{\�����	UˈM�v��)y9]m��utք��/K���[c^mb�<��s���f3�]�q����(����
1�Ů�\m��x臶�����������͍˸�q�<b��n��xi{��\m��ٱ�n{�1���6l��U�ܻVKv������bLy�ۓ��<.q�ݲy��fʬ�\sGN+�Ͷ�jOS�20������W�H4��J,o/l\n��hn�h\s��l�{.�>��%�v��5���d糮g�ZA|1׈��05��K�����iӹ6׈��ے���^�]�}�Y�I�]z�p筻)�C�gP�7lM�rFC�[��m�t��$G#6]½��@Z� d{M]�]kRt��3s�K�C*%�<r�)D���&�q�F���9+#�9z������ʏ�i�#��(��_*|�F�0+k5�)�v�H�v��7"��l������]�s�$�"�y�NsE�\��֭�L{qM� �D�M3�3�A�xE3\�^��E�ƖN�;e�wFN���;Nk�ݶ�OI������%��.�w�u��nr��t�Ǎ�s�ϳ�ۮ4O^�ӳ�lI��<�v�4e99���[{F�mf`t�K�G;���R������zS�pk�]�96l�Ž�s��Z��g�;}g�⻪:�%¦�����&�=�A����Лy����bI<��c��R��X������}�N���c�n�Q���;s����s�C�2]N��z���[p�6wm���v1�����q�U@�6�f�	�J�8mB�ڑՓ��v��;�yx7�O2��]�C/cr)�z뷍�:��NQ�<��L�t�H�\l�'���z�[��ر�^cB�ɗ�Q�f+�\uۛI�69�<њENS<�n���`:��V�^suԮ7:<sY��`xtr�M�a�Θ�ꦰ��߭�=�3��km�t	�u�G.H�e[-֡��t[OA"v����Gn:�+�ͺ9k��W\�k���q�[�k2]�6S���}�]vݶ{eq���v�u��%�x��<(nۉ٫��aN�O1`d�ٳf�sg8l��`�v#������+�ޅ��v���v��Ճ��Oc�x�쑵aϦX����2��#�#NT�C5][�H���Wm�E��$#�R�`4��������~�����%ZU��SJ�U�KT�uƦ����������������h�����8�tj������-�2��q�/]r����v�X:r�V�gpqء#=�J�n�������^csO��V:{s�
n��ָ��[�9�*����͡���NG�����I�m�u����[�p����9uqͶ����ے��q�g�ݒ .m�N]jpx�n��w1��_���''��Ǳ�<���`A$�v�n�i��;vHN��]��w"��J�;�ƻqN�\��vh��'�n6��Q���t:�1�]�vF�]���>�Hݮ�ۍ�q�;e��d$Ճ�qs�΋��s��^1ӗ>�W���,\v�7[��,�\�z��<g��,�H�!���3��;�/C��y�#���uѱǭ�ې)�N���!V8��.۬m�;X��<q�ƴ�6L���8S��-nC�n`;KA۝�%�9��l&�z���gt�='[m�2�� N������[��ccF�V�6wknT�����W��2������v�Ο[�;���E��:�N���=�Þ�x�w<� �]ǻ3�kg��mkg����9�����vL�s��=;k'Z|���tt:�1�zʴM����\�Z[>�s��\�r�n�h7;�O��VO]���.��kB�ncr[���{��swc�9�x{a��9�][�۶3�g��ZΗ���v�"��`�u�JoGM�9�n]0G���燋����S͈�g�e���d�rYc[���OV��ܔn,��m���]AͲ��n�M���ہ@xϫ͙<Z�	�s���H��vN�3�غ�^8�gr��yj���t�A�p��eޢ��r�ݹ�yv��n���+��U��-�p�s̖����I���k�$����!�k�]���Y���p�l��
p�:�L��������&����Ṻ���cź`⒔�4P�
I�n��D(Q����ꔗ�����f@$��g0x�ױb�[\wl�.�Uَ3ő�k:mǤZ緻q�v��un  �^C��P9w!���]��T����q�y�b�k�n9;=�˼tq�ch��=m��^���Ue�]��:pc�cl�pWrUv��Y�n�Y�^:�8	�wm�X}�w�74e�	�n�ֶv�
ݺ���t<���^c�"�x�2�{��m8ێ_<�q��]���r��8�6_e<lɔ8q��������3���7��N��5�!�Ps{J�&0�M_jq
��U�qm��Gmt��S�>#H�H�۶�@cMH�p[�#aB�-�=��(x��d[��F$(���}G�͑$C*��	�:�d<�DD��#bT�3��^�~n�m��7"
2�v4���"�����a��6��@���׿h�c�>A��|࿝ʀv�ψ�1 Nx)?cC�Op�b,�A���0��es�;
��X1w}4!�H��N�G p0�H��_*W����
�9i������}��~��+���p�#MC"����3���VN�).	�Fq�wd��wn�!��B��_CG�M�(��_�@m��L�8���u|:����D�"�J2���B�-RDhH#1�$yՈ���o>vɕ �&���G:��C���gtq
m�"�?+"���w*j���D��O{T� KE����Ϧ���X�O����N���t�Ha�d��^мR�p1
�#pX�2��m�![��:g�ҵ(/��<j�qyi��aa���t��6�E��I�ԙ��0�̫����c�)t)8���hn]	6�>�=����N���������E�Q�z��u�XV5��y��3��yBa�7�F��h�%8$j�G�HGᒶ
?/g�PD�D�A}r����3�Gj�q@��`���!�Ú����E��U?f�ycL�7N'$N,z��'p��z4�īE��=�f?o�W=��5ƻ��N4JN ��ӈ`�ƾM�TO�dV*!��'�E	D�@�Ӫ��<xF�酅{랫Zb��#���uEkٌ��-|	�:�j��P�@a�4C59�E�G�#�o��H���������3I$2�lc��8:���Q��^��enX�+v�#��t�C
Q�����a�>�s��,��jț�d�ε�Y���^n��yi�Me-̓�)#E�g�)��t'z���@�f3M&�q�>�!Ey5=ʀ�ƶ���66C>:���\��Z.cb���+�\�kKoE(LJ��˰)hiӗM�B����a��� �="�6)�T�Uo R3H��U��(�
����Q�@�2�u�G����$þ�l�yV��Y�7
�q�jj����l.���5"gh������bZڋn�\[)�k{6�cx���ք8�1~Z@-!R�Ү��m��Q$_�Zt@�ƢH	��@i>����������A�eQ��x�?�k�DV�\�8�F������L�DB;�P�|~��e�S��e7Y�	�D#}��_Y-}�*�,�'��)ϐ��q�Qb����ˢ��x�8�x���*��id}ia��[��z�Gdr6���S)����*�:e�l"����ry�����zkC�CGR&�	i��I�ynADLKo�(������ѻ��f���Od�[1���hYG������V�h��^+?;�^y0�"䉴�w�F��zu� 0�F㙎�ٹ)U�9��j��ㅂ���5�`���}%}��m��Y�gH��Tj6�����@a����|��ءfLL2>�������ư�c�7�-�W�glV^�ܫV%d`���e{��rbE`��m�������7�:p�uI��;��U��ۭ�_YU���4�5i�5q�]�!�U��X2����@m[Z���}���f�_���kó�bJ���eHT���7�31QF��^go>��P�ou�,�0誘{a���CD{=B��L"�%IRL��>��熪;�)���D�9F�EF�5s��L_Xؘzp^�L,ࡊD�7֦%��S6��}C,\�胜�<\�������[���];s�Q��Ľ��n�Z"@�O�����"u:@_&��_
*+���.�i��=�K3��-�|)5�`��54�TWG�����E�~)p�"d�����Q�p��j���7}m֪�gt�*���X)�8C��aB�}��� �?I�_T�x�X�s�1��V/��y�L���\�8,a��?���o�4p���7�uN�A!ѩ�ܩ.�f;G����F�C -���է����l΃4��0��&9pL"���-�[���Q2�������D��|�����B���Wk�/��5e5BU":��^#�#��(��q��D7��_�tɄi���M7�J\2Ǆ<YXY���{W��n��f���_
#����}�:۟Ogj�?��6ОX@c�XwUVő̈:���95i���ܸ�+Sv��ӗ}a�Hh�	4����A�놷.�8�z���ez���Aކ�ԮA#Q@䪥;=G86Г�8��Sv��q/k6��Ҳ��֛tm��0�4��u'<�۶�v���D<�y�b]�t�n=��m�x4`�Vs�s'�׮L��q��x�;����q��u�Q��o���s��B9X�j�m��p��Fy�<����*��z�S�s�c�c	Iۣ���&�1�7f�˓)u��@l��vѷI�7l�OD�e�=�A�c[=7]�A��\v�u�s��ŶK��.:�8�m��Q�S�͊�F�}����-��� 0��ދ��]�衧��$zc�[e}�>�AZdEE>�	"�T�A�`E�#"n��?A�~myQa�Ñ��_�da��G�Tqa}eȋ���W���en��$t�x-8��).	����O���_����z�ҟ�"�i�(���N8�㧢�i��z��B<��4C>�`a~S�ʾu��#✵\wWӳJ�SN��Պ|-	pV@�B�2�A�����&E�䞊w��#Ʋt~��~��A�炃v�}?
�����DaH�J�r霴	����m����w�O��7�{1��㆞X+#.f��v�h��h�X{����u����2{����A���H���l���ZE���Ҿ��DI\p�oVOi?������*c����:���s=<��潮g���6ն:�]$�&�X�Dۃ������Y\��uS�^!e�S�e	@Q���b؅��UY��]��\#E�𺗄�*0^������YN	RӐ/�ܳ'���{ݐ�3�Q3ʞ�ئ�{��Vl�A��wp�	\v�+���o0�� �v@ ��ՠ�!坽��d��uny�P�3`N��1�z/��hsˀn�ȭ)=h6���?�u�:����96G��~�wy������ik!�D�$-������l�R��p��$��:��jq�7�o.9���͔y󉫖ĺi����Z�_j��R,�HUn��$�%G&S���b��e�S�FgruZ��jPGD��V_�E�kH��C�@�u#����wX�����E$�%J
�(��Vu�UDȝI��}|�`���'(�I��@���YMQ�G�c�h��^C�u 0�k�"��k��P�4�>��yg�ۗ��[����($��q��C����4q�Ą�z��[�M��ݭ�lg˻)$-�~��Ȅv��ʔ�C��B/���hY�� UO*#,?>ɏ�ͽ0���^#�}����E\�i��BI%�~da���#���ك�A҃�~ƄO=�&u��X?0W��&��HB�Q�_}X���?{*��,�f��|��!�JaI x�u��ʞ��B�}�a�ֻ� ��/W=1aM�'D`'�̐T�S��c��n��m�ÚJ+�������{S�]1��|�j��du��ڽCA�i�� �|�U��iP��
��#��#���˩���}�}�r�k-(\�8:��g��������UcHZ�tG����
:E�읱�e��0�wAda|a�;���i]_WFJ�3Z�~gO�Q2�TB2B�����GM�,���!���D����_�>:Y����w{�K�UZjH�*���{<W�Q�&Q��U�4q��?L�o�8c�+73nb�O���3W�l��b�-�Z�S\�[�W8�.��'ݏ��$q\
\i�sU��[�[�����}Ih��^;*	�t�����J��C:l�[�����G0�����M���c�-��e��Ԡ�f���$r@<z(|G�C�_�=4�c{;t^^oqQ9�E�+!�u�o&pTF߯=X>��?2��]A�t{�>I���������.�-�Z��1�cH�"��r��2��ж,� W����u��s����B._���8â������x�p�����VzM2d�i����B�\z�<G�nPk���Ф�C�.�X �tR�<Z��}^2fÜ/��{�n(w�-Ǒ�4��Z2�OV���S�᮳v�e���/��8���R����Dw٧���5;:��{�����M�L��d_n��ize�:cuT�!�	�����N���@OE�1+��}�j��?�E��񃎐/�G�}*WJ��""�W�ri��f�F�U�yv�7�kv��u���i�ױ=�br�G�y�X�`�>h9�S䘂�`a�����I� '��Vt栈��l���?c܀��%�H_�b���]�z�n� B0�����آ3��_Q�������e��r8�pX�,��Њ�ټW��B��.���W!F�78�� Y��:��d�#�Q>C>�r�����T{z2���nm|2�j��^��&4cG ?Q����	�n�)c���1n'��dA9�7i�Ȋ�\��7����\N�P�w�S�ࣆA��U�2�M�@�#RFӒ�Ĳ0��%�b0�A�-���"��p��W�P�����9;�7�:i� ddC�5Իd�۟7�@q%���ԉ�u��,���� ��ܐ=�D������XҨ!D|�]Կy�!�Ϯt�HF��}=��A��@d&��3�R\V1"�f�,�����8qkf���mL��*��ü7n��&\8omh��̵ٽβ�D3�z��];�ZOW���=m+��;�וx���);v��j��i����j�f��pXp"�˂�m�<�V���t\��%{I&�v�Ҏ�x۪��`�e�^�P���s۝v|:���<h�rp�����ܨ���벶n���;r ���c{kj��.CIj�nc<�sZ�z�wbؙK@��-�!��=
��5vn#yx�,��'�y��8;&��u��o|wݎ���'T"�-gLL��A5k3M����]���U�lF�ú�p��Rue{Y�.YKm۰����t�35�T��uCuG��`	w�`�xf_�XQ�j�к��;��޽"�՞̟��u�wB��G5#�����:���ԛap2" �#J@��þ��t��z��䴅�z���y��QܸȢ��n�	c`q����-�.���&4\�k�b{�A$&	 M�"���q�H��
�Ӛ���4�2CSׁ���H��c@��9�@�F.ЙW�])Lx@��#�ZB|�t�2�=ߐb������o{&���F��S
(һ3�^'�Gd�ݟc���������	�1;�T���hv"v�������>�(�M��eƣ������e&0��1?3Q�~��K��V��v
����Fu=?@B2���#�,Ф�o�U�G�
79��]��z�NNB[����94�謏͠�/q8���C"z@�l����,�5�rM��n=����C֑eooj�?klB_F�W��@pi�"q�$QPN��[�<wn1��ɁŤOUM�!��h�Ǹ�-�)"������da�����<�a�a��Y5M�f����
��P=w;�ܲ���X�$�Re��V'���-�#ū�r�
�t��g73�bU�t�ǥ��o�!��b�hCaa��Pdm�}������^�I��C�_q�ߜ���H�����N�ഋ'ﾞ�Z]�0Zﴖ�����w¸}Q�;�/��ʚQ�ʄ44��H��p �#�}��@q�8OBl�ِ�aNK?P�Y ���a�+]�վ�#�X�J[ϵP/%*8h��K]秂����D	�].��/)�EGQ9W:��H�5�3�P)�ZQ�$�4,����qQEjR���/6��?3k4���8��w�����W���vt�d^.��4�~æ��?ks�Gs;;~�hd-Ge�X��μ����m�*�M;>�uG=����p�nwprG�˭�Q����FH$f�� �3qG�a�p�}x���6�����t��jt��E�.��[����Y$+��!�KAn@0�O�9|,�4���Q�&�g!�����!��5��t�0A��T>G	�1�"�EbH�.�?&�[�3���n(�R&�8Q�S�P� ��٭�pQ��0Ffz�qE��u��E��<�엊��iڌ����ܡѫ�O*�%���)6i���f���&!I�WB����}��q�r7�70<�������E��dQg�Dr��r?�Kv��-����*��u����܊h������C�>�'��:e_ݷg�8����F8�/jA	����A��\��yP'o3��^=B�7Bp�U��%Џ1���-U󿯦�ƽ�ץ?Xcm͘��Z><�f�ᇹ
��U�wR�hc�NX=�9ֺ�k$�{D�Ҹ���Q�k��/�S3gn�� &�e)��W\��2k�W22Q�g]�Y�C���!*!<1����2�o\��c6&�\�f�&e�I��ݣ~�����a�i�ғ6�Yb�f�R?1ǳe�-�Nr!�֞�t�h�3�3&��fS]|��L�i#��s�*׺{�c,���ɐ�-�Wh���wp6��!�^a
�j��۳fp�KE� �P��O/DrL|p��3{N��۟<$^@�j9�}tҢ��O��b�>NϮǺ �5��a���*�
e��]#c���]YwK���ICL預��pD>;�fo\Y�ԧ�ȸ�b쓳;��s��9��.D���U��V%W[*ef�cu4rx�"u^���iT-2$�a=!�������\��uֲu�&ە�)#W�յ�RcO&6��o���	�{�1�'t?s��2�Z�w���o�Z���p��z�نDR'�n���E�=�a�縌D`�<'���m�/$@U(k�Rv3��f�*�L��lC�VJ�ٺ�q�#\i���%�a�]*mB!P�� P��vU�@�.����.7�p�P�!1E��"�� ���ndC.����i�@��4$���'	IHLP�B��7���Cd�QN��V�@�,!1B�ڄ!B!tH��%����#�!�1F�P�B[�}�ii�BL����TX�.����� P���	�}Yj� P��Ti
E+mB�qB� P�(@��2����p�P�Q	vZ��Bd,!sܫ�!
BS����]�O���/�LP�B߶�n�O� KǈR(@�P�B]!1D�1B�� P��W�|}ES��U3N\�r�(B ���I�H��m��(b��Bb���^�U�@�Xt�"�ﴒ�$�� �r�Bb�b�!B���3��qBO���p�P���j(AHLI11B�����"��*� �� P�(@�.�HەMB!}����aD1B��H��(Rڄ
B� P���|�n��*Q�@�sB(�C`�W���V����M�'A�u�^�����̺�v���}mJjj��*r�j�u/(A�&(UܪP�� ���� P�(@��&B������\ P��GmĊBd&(@�D� P���
�/�
�
}9��B���
(B P��LP�B���IH�'��U��BN���b޸��T� ��KP�B�ҡC>!&B���+|�eZJD���� P�ڄ
B�{��R�B����Xż�&P72��M<��B[P���&(@�K6�E
GE�)!)}Ɉ���P�BZBb�f^�s}�w«�/
� ����B�
�P���I����n��.
BX4(@�+!1%TԊ[P�BT.�"�
���j(�iIHLP�B�� P���^�j%
(A
�w<W.6��
���]�����
��I�B네��&(@�r��̡��QM5Jj�1B[��.lʄ!B,K�) JE��K<5$-���p�P�B�q"��Bb��Z%�i* ��&B�8R(X��ʵ K��
E.6�T���ȋ!Q	�(B P��Ϧ�`�HK�� P�����@�P������/>g�JD�!p��"<�q(P�B]!1F���[P�B[�/)��C	�虚sO!pP�B�'D,!1B
�K��6�`�)!1B���[�� P�HL_[IH�[jD|C>���* IX�*�ʄ�7��XGH�B]=-B!a	�*!
B�!`�� P�m��@��iI�&(@�P�B]!2:D1!%
w9ɹ���"f]L�ɟ�gI-gmp�N�;ؾ�61[Jޓռ�瓤{���c�����Z��3�	�}ۦJ�!���|�p��&�'<�x� P�{�r�
B_P�B\!1B[IP��+!2���w���j����@�B�� P����[j6����� P�%�d)�>��, P����(A�&%�(@�.�IB�sݮП��\�"���(�BQ�% ������I1BJH\��! Qd%�]$��%�|����\"DB\��C�����c#H"n4L��R���b�r���������0g�km��ԏi��9���TԺ�]��P�n"Hd-!2���
(ALP�.��~���b�
%�R.	&(A
�LP�Ĵ�"�
�������X(A	>9 P�LI}��+m.��.��IS�}6�����{}��/}�!1B
[��p�P�HLP�B ����p�P�B�� P�{\) P�B!Y	�#��u���Ҏ7
����&���/}wJ(@�/	U�6(@�kj$�p5$)�ݛ���
DT��o�̣���,P�����	\� ��!w\)'�r�B!i	�(Tڄ
B���(@�I1BS߾������	z��
B���B ��d.���?]j-%�*�!x��"/���������!1E�1B�� IxL���5��Sna�t�UUd.
(@�&Bd*!1B��@�*!2HLP���M�@�Xi
E�$�[P�B�
Eࡉ�*��*���p�P���qC]!t�Ė�uoy_m�b�
(A²$P�B��x��@��L��>�(A
�LP��LP�-rZ�
BϷw��\#�!���P�$����Li
�H���A�$�L��./��sC��*T�S.j� P��-!1Bmđ-B!h�w�E{�/fȡ�
$��.�uZA��
[��q"����`� P��I
�B��������%�J�!1B(��D2�LP�B�k>�JJ�!mW���\ P�B!Qe�@�6� ����=��4�$&(@�S��6���BZBb�"�@�-!1B P�]^o�$)�m�L��, P�ڄ�B� P�-�9QB����"����7�ڄ
B�	�P��"Z�
(A�it�B�
P��|��UƎ}�ԗ�d*���`�%�W�b�
.�����+/�P�BR*DI�b���j/��!p��+n��¡B	|B�B�ґC P�Ϲ=W�!������
H��(@��IYD,!1B�K��i����y|r5U��	uL!8�F�.���܏�MK��|ѕ�xVj@f]��؄�ʚ�85���+�[IBv8Im�$�H���6^)����	�]���g��'E���#�:m�Ŵ�������m��;+��q��T��юGm�ovŻ`gY9��ˠd��s�>"t����)۱#�[�Hu�k���v����^زf��m�%��]���笂��s���.��9M*��G;�ӳа��ƞε���-֖�u,��:��.Z�k,����kZڸ�퍞�<�v�Q����X�2
��l�7'�봷U���nc�]��Z^$�� ��	��mR�!B!|%�ݩ P�ڄ	/��U��ʸX(@����!Y	�(�]������L�ȎS��*� P�+��
(T�I�������!X�b�����X(@�
s�R�{���a'��P����m�(@�P���LP�B��ڝ���P����E��Q�dC!��Bb����4,� "�9�%��bI!-E
M�O!h��!B\�L*!Y	�(]m+2��RBb�
}�j� P�������y;m��Kj(Ar4��(B.Ꙅ�Eo�>W!.����ME�Y�O���_}~���{��GW�t�j����B�AB�4c�Y_�����Iu��B����L:�=�<����$� ������q��P�R�q��}�"RٓG�,�EC+�aH��rG#n
p� [�I�ƌ�D����I���$�?V���Ҳ�㋡�Z����\#E���!ڄH��]ԳW�+�ȶ� ��)4�HdN@���� E�};%#��WȺ�1�[ Pg�i�}�FX�����kXD�xT"Η�4l��;Wm�-G8e������d�-@�,��m��w���]�����j�Y/n����[E3u͵��k︦+��L6f�^��?n�h��~|�Ŝ[�<!�r�{+���0�ʘBq�̤N2#Q�[�r���!�i�&g��K�F���Ҙ��`��&@|�TƊj���U�K7wpt��6y��3s"�0c�n�v��L�fY��p���0�3X"on�vrD��"�yՐa+���O�	�-�x5㹵H"M$����o��avg�!Z|���u7�X6�%(>�P��(�iE$-�C�kQ?<lY�y�I���!��u��wVv�;s[��w�褎q�4�]��VŚ��_��:3�#P0�r�K�5����0��@�ϳM���ɠ ٴ���a��bE�U}t���K��5>��󲊺�s d�:ඛ��|�0��f�1Ĳ�,G%UM�/��"ŝ���z�j�AJ낛vxV�z+���-|'F_D~��YK����$i2������3��rLP�EPC�M���&���{u#n.�/;���
ZM�v�u�#��#����n��I�c�0���#�Nt,�捪I��>�`�YG�t�(�}�&g2UiK=r�;���������A�.�eeϣG����������Q�v0�(�@��0��6Cq�yR9$%	}>��{�L|���,�c��b�1)ns�ҿ!�9��W*ç�m�o1e[�:Fg�&D[�I"Q�Ԁ���h�{�E@uǆ�����I��̀g�(�>Y�j�s�P2^!�Z� �{����ҭo�K��_����u��㍝:Kv<WKb��;6\��E�v*�sVl��ZE�u�0/����a�v�?D��w��^k��#�8~����HX�&LF8�O�XB��+��eks��C5J��tD)��AE���_#�=#��ۨV���q�7�>�@q�0f3���p.��Em��p�?nm__���~gƈum�"���ޯu+)�g@��G�©� ��]^�h3��i��v���B�F���vzB=�_U:�ٸ��S.��)�Z�P���ٵ�0��ͨۙ
�wQu�n�4;�B�h16�J8�{P��+5�ТZ]��/�]N>��G��Ĳ�(�Ϊ`��>WU�p��$a�!��?2�S�KV����a�Ƃ� �ЈH�m8۫/�H�F��CCC~l��]֍hH��ղ��Cq"����,\��U�"��"�OW��6�9�Z��7v�HV\ �6~��4=�`1Iȕa��Y�4Mc����*?=@$����]���kD�I,d=��Ht�҄Rƀ�CH�~�=�j�V-�XKɔU� �t�t��:��4�[��q[]#{�pkv��/E~P��ӛ�� �@�%��`�k�1i#�w���F�Xӓ=��wt�eu^Fwv��3sDW&��������ډ�W�6��u�Da�P=Y��W�M�s�I�n�;i[����
��GW>�A��'�[H�n9pP�AG��@���?�kOą�dQ;�U l���nÐ��h���d�ҳ��t��q�FM�M2��]�(�<�5�C1�RM��ݹs���[��d�Ĥ2nn�훴[����W�e5�l�ۈ�ɺ�b��5�5Ǿ�L�	 �Eq]�� ӆl��n,�U�>��!F;�̃Ҟ
Uoz�/�T���7+�CM�eS�z����LQ#P��s��8�C��RCC�#��l^�`x�e`|�'�wOۜŐ�!��҇�ۖ���p�]�
�!H�=�s��wA��{�z�	{,�,�<�aG 1�Q'O�����I���衚��	 (���+���:�!�K�4�=푇��u�r�>CM"a�A��b�XN���^�[N|5�,@�>"/�-�ce93d�I�5>X_T�D���j�w�6P"u�C�U!�a��{����0����ÆY� �9�֟�/���Ǽ�-�1�c��j���o�4]��W^C���ڄ7����aB�2�h��c�1�Q����!3U�C��$�H���۳A�ej��b��G���ټM��w�6��ĕ׶����|r�N�ͤS���h�챺>����C}�WN��mzҗ\��rò_��h����1�'ܸ�q6+����[V��]r
P�����=&�zm����
n�vzf�H��ԓ���YW��o�]r���y��xM0��ݭ�3�<�۟VG�뇙�m�7�ѻa�74�@�ۃ(ln�蝖MU�b����j�:�m�#���Gձ�ssuԸ�`L�����y;v;\�r]v�uɼs6'��EN�������ԝ�����ӹy��mu�� �����rl�snzS��$A���^N8���N)�oý?DH�������{���Fp��-޻4�-;�� ��8���~>n�-���ȼ@ؾd{sh���f<Ƶw�mz[T̉@�D��O*�4-"7x8I���W;���j~�B���ǀ�#u2�8�=��f��(�<F�g-�ݹ!2YCm�y�k�ď��[*M�0��pP�{$�4N!veuo�4��K������Ma�xe��9S#�U'	����#"� y� �U,��L!Ml�W���q��EGR��_�����VC�-+�3Q��VP���l@f�6@�֚#iJ�`��x(LXE^�TT��~��x��?ts��@���e�|�j���:S	n$��f���ddB
U�`o����KuD�,�8��p�b�]����r��B���kud<D���D�z�� <CHg1	����!df�3�n�<�Y̹��g،�[���
ݞA^��[��t#OYd��J��Ok\��(��C���Q@���1A�:kR��iM&:�q_<��GPX����r*�X���.[��}�9�H��Ђ4�?^�_�_���=�L��˘%���X�?�Y�hVF��\3e+�x�GT���:L��ud�U1V�Vy�e�٣���9�_LS���fo"����h�r�8�y7P&��<����W;�|7��Ȝs�hq̜?l]�z��(�D��|���[������:����$%��^���H`	5
e��+��ΐ<Q��3�r+H�HЏg����R���� b�`������ �#��M
�0�=~v��ܳ�!H�y�i ��Ĉ�o9�ښ�b�&�k �I�4���'�c����q32Y��Qf�;�A�R롋����d��B�r��N�� 7e)GiT>ݷY�}�Q��UQ�M��\�7��FP��F�������@l
 w�O��M�TLo+��
uJ��FP_V�2(�u}
�hHQ�+1���0�<C�BwSI|HY�Gm�a���-�s2��5D8������mqٞ'�vܛ��r�����Kp/O]'Y����Hq6���U�j�;�5�5�R��0���0,LVx�l �	�V߼�﹒�҇7��Y�har��F�1Yƭ�����I-l�h��>�DRH�R8ar@l������C�]2�9��8�أ<|�2d��!a��(Ն�8���0'6Mu��CH�f�cx�
ߪa�]�$�ˎtk���E�`˶���B�f8�r*�@ĩ Z���A�����馬�	�lA|�S8й��D�]���֧k6�G��[�&ރ���	�;C\�/L�-F��,P�ʞ�lm�<��^v������D�m�Qb�j�B��Y��X���l��0�=���5��T삼��n�c3#n"Y�7 �!@��=��.��W�炇��2��"&����*����dY�+*�d�D�2D�A�QqcV2D��+P�d�6I�����1 �T�8"eK�/kh�R wޭD^숅:��W��%w��6�Y�@�3�n�]�z�M0���
�z�6�.����y*��
�vcݽ\K�>,9��P�Um��*�uЈ:V��u>D�bË���7�.ѻa&��_ӽ��F(��WL���q!CPe��w?��>�b��� �I�u�����-��1�n[�NO�g�n���	��˴�߸<�#��%*Fo�VF����{6���ߥU��f&�[p2{�a��=W���ʑۮW-��{��v��`�D(�H�d��m� ��zm-��+|���,�~�w�{֌����(AmB�c	:N�i^�(L��b�MPަ
 F%kZ���h������ׅ����H���јB�q���M���,��J�)��$9�IS��M�ĊG�샅5hBR�8-�xom��gwmm4��j/�'������)�A��҅�f<��4�*X�M}�"��{�8�[��#I�C>��]�{ˎMB&�][偫�jc.�Z��7s� �v�WW��xm�h��*p�i�@�D̐�J�O݈���")���f�c�DC�P�H���s��W`�L���)���z��Q�Rn�8��H��C=^�V�Z�|ڤ q��燂�r3JR�c�[V�P̮�]��5%;���.��ç.���Ѱ��9��rv6�ۢᲺa��vlf�˃I���^�rտ���,��<q���;�|m�h wU�H`��wqD�$	7k!|&��� ,IԒx��] ���َ&n�u|�l �ݠ��7�|���l4�m9�+x�?/!D���h��]�3��X��/�/L7��6�)IF�){-}�ј@,jei5$۞�ţE��=mRi"p���HeҚd$ȉ���B�&��h����hb���r��
$��b��X\e�'/D�7U.?*(\����^AZ�y�K�(��/�@0Q�$\{�`�$�f�R@��$�-��z���!�܆�D�͔n=�����^��׺�!�}uʄ�xH�t��k�JŒ�:	5��&��$����,K � �����FI��X��N�J����#K.�$��*ƺ�������Z��f\��޾xj�ٔ�S[L$p{��3!$/���]^��w=�Vc�M^N1"+n�j8ɋ��At��s�Ҭn��y$"�tm�J�ŷD����q����jJ�yC&N�Os��M�4ɦ�ݵ�MD�J>��gֱV�[��䞻��e��S�v�uvM���fI`�ZpK�I*n��WJ����a�H��"�)GIX���Un�[!�����H����̗Ir7�����⾹Ǻ��3&`��3,��s:�R%s.��;hRp#ل��.�{���V3@�BQڵ�O����]�:�u�P����d2�h�l�f����;�r�I#`ĺ�g(�d�3e�n��XXE8��L��o��]fb�vW�g%��7��B�o)�p����L{�е�Y*h�PL6�����F��0��5
ۑR�8�1a���Y�u󰊑n��m^f�*��cy)�$e��<}L��(���2�)���ږ��N�MH^K�.\َ0�ٮ���I)w#܍����;���<e����՞0`�t9����QqWv�qǡd����}�:��3T-O����\,�,63�b�m���X(��q�&�U�����`��u�+T��k�*n��*�_^Ҿ�}��h�iJD��]��t��rtd�Fʤ��O��U�X���Y�p��v���
�E��嫵j敪9���ZQ�B���w-3 F�.�:8Z�C��N����ۃ�!C�hY�^'���bo�z��$&Fb���$�IP
�Uҥ�Z*��v���������������=��7��>ܻe\��gȻ��O�E�n�"[0��uu��[�hwu�]q���z��w	F����K[�q���!�=nxǉ'��n���w:N.ݞ����s���]�l����j�s��#�/��&1N��v<S��gq�N���nw$u]�W kF��uH�x�����XNpq�tZ��<p��CvuVۗN�8�y�r;[�v�5x�v^M��l�|�� ��	��\q�϶�=X/ ��َۓs�b��S�]L�v�uúڼ�S!�;�m�u�W\x2��#��hG�&��-�#6aFs0�h��n3<=����Ѽ:\ޮ�}�;��m����%��c�E
�	^���Zܥ��kpົk[�V7FS�ԐknqOM'm�;^��ݩ�j3��_[���d�\�s�E�8��k�g�6��
������'t��fb�u�����T�7k�����1��n��q©ԏgq��v��^�b�5k�����vӫ�3���V�v�#��OK���T�f��f���n���,*m5*ޮ9%�ZV�<����ًÄN;	�q�n�6^Nײ���8��;���3�Ǖ�x۱4+��9�c!I���[s�MvC]ƈ7\�k9�n9�8�Qk�0�=3b��ř.�Q^�<*��v�k�:!
��obٸ�����b�c>��k���������N�A7�:b�۱fM7��oDnܓú��c��j8��U��%�ۛv.mm�d�-�z�xN^ܜ/k2v�b�n:܂��Ք]��W��.�q=��\��n���=\Wn�pYz͇�WG&�.M���qշl�]���_.��]�hN��sk���c�83����л�qpv�r��t�2Q,n��K�U̺�\ݎR�t����=+���w>�2Q���*�웑�g��]�|��/|��َ`�ў���\=��g��6���ti�e^:��{����qq�'k��;m�n3и'��:��	�˫���/=99��/R�V�UR\Ov���`v��zMOZUQ�\\on�8�d�� |���p����ןj{lu�S=��)��@͛���#vnC3ȼv{h��=mn��a+���W]g��������Н[�oZ�y9�\kn����,u�m�c�vEsv�����\u�a���a�@��8�ɕL=��]^�۰a蚹i��A~�۾~s�m[<�A��X�G�z�`�l��F�U��Z���:	70�O�{�{[L�I��,w~�����/�@~$N��h^-,����A����Φ&�s���A!�AÈ�Gn�vr+/U]X/�P@�$��#��r�E�7�ʣɽ�0�R�q�౧�hm�H��pQ�Co*k��L�����4|$�w���@S~�MG�a\�v��)a��7�! "k/�,�B0I�wj��t�w�Xd-i*l�Q�NA>�c���%����v,���0������R	���h��/ލW����=�(q��NX�P�
s��y;]�+�$ :rӮ4�9Ɩ�E��E$���$ā�����5��A{��x�
�Gu�OܐΫ�A�?��h
��v�$��@����&�N���W<��X�۔pO�Î��;D���T���@{��N�@!:��_����(�E�����<�;�4D^�I �@�U�BL�͆�2��F����3��h�vX`�#�}DP$S߭fl_��@�EL8�jI�u���p�3�ݯ{m;=��s�s�ƒ�B	'���"��M��'�@3FȬ��z.u�N���h��*m1`$S}4�H&�HO��__�%¯36�"	��Z��Є���m� �Ŕ�$�(3=Ԉ�����"�	9���$B��*��a�$��ui#�Ft�b�ߦZ�� ָ�<~S�Ϳ=�S���^�G)�Z�\ΝH�l����܄�Hg�m6VHw(+0������<�;> ����"�eϽ1h�r��=��#����\��/DIͻ�Q"����	A!�_Q&'�g�R�3�,?==�9N4Sq�A9$��l�D�[hb��f1di�F��AzU,`��s�Z?O����˨w�sh̕>�J�0�@q�W=�s 8�����,ӯ�[�RPʙ��������,�T ֻ���L������uV s��@ �������ݪ�R�@A]k�fK�ʹc��^�ǪDy9ƕ�����'�|"A$aEQACf�jR��L6�9���3�xCi�6r��g��v=֦�:��ɻ �(���.�&�{�И�jE��Ѳ��� �s�yC�`����$q ra�~m�������6��!��p��s{��0mu8�5�{G8�W��2�X��Kנ�Tr�f�֙��7_�߯����k�#\�z��xh�h���a��`i��)�6	 ��G�=�s�*x����&���>A�2kQ?r��q��.	2�4��Q�A�jL_/�p9ro��s��<�Wt3���O�7q�� �ժɼ_VG���A��p��'��d�C��X�򳤫cG�?k�_	3v̝�	�PT��a���&%�,6ܒ9 �M�'����3��xU�u��'� �M2�<��!M�Р~��(V{D�[0TqT(����-��W��/|��]{Ԭ�a�P6fy��26�`�F�]�_[K:̦k;�� Ә��F^�7`��(�vcdD�95�>A o�RtheL��������}(@���y01����&���q�_&I$\TU�_]��P�O)� Q־Zr��U���Y����k[��d�giX7�B�B�̄�-t���f�D��*-��MH%���:��&IARQN[��� ��q��X�C0�C=���j��L�=��[ ���2 ���瘊�A<o�L�$��S�sZL�I�	�{Iy%��@�8�@�cLD��u�k�sͭ��÷Z��G���6�l���c\�� �P�#�g�=��V�?nM�;�fWDV�:iN����Me���e!"j���{�t8�����q����	ێ��B҅��t0�{n,19Gn���"�k�J_�}�\q��¯u�B�p��͢�Җ�_'5b�c����ӷ	��jC��౰k�A
9{�灎���/�=٪1x5�y�L?�ot���
B������+��n��2�����a2`P�R�
��t[^�NqL<}��_6@�Y�Yݕ5�sE�y uͱ/ VW�x��k�����M��<Pnc6|η���J�ޜ��yL�����:�6ء�n��%ԏt'�j��f��et#C��̷-j�LX=�c�\W���g�}�^؆0X�7$�CvIG�Z����嵂��Y�JI���Lp"��<��9Р,BMd��
��7�1@i��0�L�Ū��\�5
��Q]\e;q��Η��/Kn�&ع�]٥�ڰ��H���;�����)���7����tBQC���B̞6����w�4n������w��V�L���p��Oe�4~�t���uR���`�j"b��q��@5�3��%�֓ݭ�w�k����f�v�t�SG�k�^�<���������d���G�c�{�*����"N	�!�>�1+!�4m���
?}M
���+:(Qv�"*&q�<&��L�uN*��'R*㺫F����Ǆ����K�9#-�c�g��Sx�h�^�[}��D���}�q���}�}s+��ȳ�8@�u��4o�dL圻�N��li�)}��ݝZ�)�*FLn�̱q�x/^w�V
�f���w�*�kכ)*b���c����T�E��?5��c�#s_���gZ9������|~^d��퉧	�sX��*b��뱤^=�7�^:���͗7���zy�e�f���Uj&�^��gFz��9��5��m�,��.4�S�$xۤ��n`�gv�O���.�k����^n}����\Vw.C���<u	s�\���{X��e㱷`�r��8*�;��[v�h�grS��1�Tvc���%�6���vzN]�V��]G&��t���܃�b��+�A�9N��y����x1�:v�ۯ<9�3�sΣ�oi�ɗ8�[�O�D����*ε��kOOFջ5g��[��kHh����t<E���s��;f�!^J9�3*bG��$?/��*���}g��4w�zk�hI?SA�T�T��z�b������׆V��C9g��+�6�25NF�0��J��.�J��R_?�^��R>5]K�S9�[f��N��d���Ac���PT�#ht���~�0������^��O�R�8h4a͔�����O a����* ��wCrF���/�eQ��G��}Hy�UxU\��jR�����u�W^��N���<����x��t�f��*v���VB�.�_M���da�M�a��N=P��y�Ǝ����{��ףԅ��X���H2�$#rP�wi�s�O��|(k�(�o��s����X墘n��n8�Y��?
^+MSh�+EWw�:I�>�]OO_yc�Q8�)H@��6�I�,�ݔ��#���uI<9;z{uF�*�x��<Of�ϲ�]����Ý���W0�%pK^�{�~�����b��Qt���G�y���#o�A0K�\�V��{�J�k�K�����e���Έ���O�Sݞu�|��9�C���_-�WQ�LW�r���e�8ܦFaU���'<�\��!
�(��Ԟhl���������2�YzM'��&t�Uđ�NJ�K��O1O{=��qY�/H�LT���JDz��\��
 d��dE	����ߘ�7W�E2�t��k�}Ҵ\�vMuj��J5��i{�b�!�@��vH�ݙ=a�E�����'L!OŸ�p�pP�H�.�6��={8!>=���@���A�CE0��u���?�>�����'�
>5he{ �^@�̏B�d5"Q�,~���o�H�!f`���ȳ���Ym���by�Ʃ욑�Q��,̮}���Da�����At���@�����?����q;}8�<�kWn����&_�3�X�܉y��u�<�\7Yc�2"&�nF�83T #� g���Ά�~�^�̞��F���J�#��F_���,e|6�\G�:��w	���8�p��"''_��dy[&u��C6��sz�r(����;������}״�}��e��}�G�~m_�nAb�۷�Yi�^�\B�C�A���_�l����w����o�C��|�u8�˝��
TȂ�����PԗA�#.zyx���P[�äN�m=�]�CS4��������ZU˷~3���+W*B˒,�?J�s����4���t�5lW��*�ş��X�B�a�b`*2ێ% ���x٫����=[�x,a�#�Ozav��ҡ��x��#�ʧ��@N����N4f�g��8�8~�@%�X=M��rH�q��F�c�"��w���P��1`:W{hY���ފH�(2p��V'P���z3s�.��/E�o��l I��������luy
������[�=+d�h���Z�L�@\r)x�[�ǆۄ��+�܉��#�:��E�˭q�*~��0�8@��ԙ�>h]n4��T�Ǐ�!���1��\A�$JA_a+�mؽ��h����}�i%���+�aF+�A�u�BȬ�� �v�[!���LueV������+Q$�*�1H�#�r�s4n��}�)ȋ f��U9�Z��;�� �SO�X�����^�������NYU�q~�=k|k�!���	8�`��B����֧d�OJ���q�_ft3�Ӓ���Y��#H�Q݂�Zo����5`�
��]v�1��nD|�Ϊ��"��N�k����p (%���#3��Ye��M��2gahVik.��ٴP?ZyH��VG�ؤl���?P����Q*(nG$��{��?���^�Q��Ѫi`�ۼ�v+訛]��}/\�[f��P�g�=\��X���[?<����י���f�1IL����l������.�\�����a�hN��6���Aa�*�"��Y�`����C��g�=��n���z"��]����R=��E��U��:�L�~� �I�QŌ^4!��֨�+Έ�Z�E�2�v��ƥ�0V��tu�L�?Q��W`�C�IR��ў���9�-��L@��Bю*r�Ȉ~�;�����R֑��~�'|�{����lv��Ó/kʲ����W��n�9Hm��!Z����p�M9$T4ᔾТ�ކ��~�x��G�Unw��:����|���z�}��][gFl��0�́&��=x~��������M�I0�
R�;��>�؏�{OT������+����%�|LT�n�j���I���b��-��F�Ӣ�����b^�0����NC���e��Mt)-31=D��p��mL�.�T���t8g1k�Frx����.¦!�7Bhz�(�(1��b�[���X:�i��D�n6�UWL�fc�\�hͺ�/��>�v��A��D'"a���:����O^s�r��ph�k��v㭸�p��WN�'��8v�N�nq2�o`����B��G$�#���X�ry\&��G7�Aԛt��z�Y�d[��&Fn���<OA���i�6�m��dݖ�Wf�&��u������L�ܛT)qx7�&^4�n3�p񶃃YlV��E�4S�=k�=C�X���+�1��f�fw�Dx�g��Iu��Gvr5���@�q������+L7���0�}ת��{�=4���Fn^Y��1F�T�`��������]�TK�鎪\��H�#zl�����3]k�&���뇤A�C����T�=�L����S�gO+ý��e
F�>SOJR���97Bk�� �щ�zF�v�Ҿ[��ټ �����wm������:�,�k'���ε|M����
8D?[�X��
L	��[�^�j�-���'{4aw���wS��m,#54���Q�ip^#�'~�;4�ͪF������l���ޛ���$�D�}�`eDӄ�Jq��V7R-�~^�X~��J��<ԇ=0�tZXG}=W&ޠ+#J&�Wh��Pg��f�t��A��i+��v�m���s�r�D=mg�JԚ�����-��j�W�&��Z��V�����/#�"[�N�W�P�1���?Q���q�� VK�ņ��H����I���+���ؾ~=X�EBSQ��a�%}�la~�8���-��{�8��b4P�33oh)�2r�������Q�d��k��(~�K����7yK����C�0�����K���]���P�T�r��+��Wr��Hj��B0Ew^�>{��U��� 1�SQ!��7N�l�GG�� vV�-s��_U���(�>A��r\r���Vi	�<FR�OV����>ÄJe��+w�8�JBb��X~4{�Ԩ���Z0(zY�*�N�����4������Oz�*�����{��R>��DOa=�c{�a�ٜ�M�i��	8$�V�dT+����㎆��<�g+x�1����>�g뻁�u��E҃�*������kK6k�!{����&�St��'^��ٶM���)��{v�n�m��N��H���I��>7j�Ri��5������[���n����j�"�͡'i|��'V�'���*���4>��9����gD�kOk����Z�HP�i87>q���]gI�`����K:�M�P�:\}g�}Y5�:~�&�	��40���l��ݧ�/�/�[
!p$�q��u��c~�w8�i
L��`�z��|��x�γ���f��g2�[o�+���;x��S.�3:���p��wm�9�N�Ă;�ro�=�o3�p=�Σ`r@ſߪ���4�U}�R�x*�{f�;�S�{N��]��+�B�x�R��C/N>/I�R�{��g��>ә�Ք9�L�6Pʕ �̭�9F���+�h>mt��ە�_�w����`#�Wu�EJCJ���0�nD�mԫR��,,0���X�h�
n��o^�2���i#)�x1)�M�ze�}nr6�1-����.��wZ��l��޾+����<^Q�E*xkwW�3�FP%���)n��׷�S�㽁��d�.k{;]Wvw�9��N8%gj�����	jb�ÇX��t�e���4B0T�(��MОvD���$3si��$0�6�Y%�o��{kM� `�V��o-X�s���g5k����'U�\ƙ�'�þ�6��P���vB�Dօ�YIN}���i���'�Q�mg�ΗR�E[3x�(R�N��z�YG)u죗em��q%ϋ�]�qd\V��k�sxhg}�of�(C�1�*�t��uCNV��9v����E�VCˠŦ��i�Ui���@fQ��Q���̛�Ӗ�BLjy�^"˙T��1ӯ$�rs˘�J�
;:��,���_F+�6m����eû�e#/�S�����7y�1Q��U&�Mgn8oj殔��][����h���옩w�.�f�pD��v$h�!ɚ�ti��AjP4��&6Y^�`����s�c�/qǲ�U��n�N���inI��B(��"��zf���z��cz��݌�����2�^0}��ˌ���eù:~���Vr�D^��#7n~F��ߋ#�2�H����HUJ��>�~�5���q3�$8k��@E��3z�����Q�.6���ff��������\v�q��K�w,N� 0�7 j�ӷFی�K0�f<;����ƺl�`� �3�t�����͂�}]���:��\��`/'�)��u���t�������4����U�y�g,��r(6A��5�I����8�F�z_9co����iP�G}�}�>%Q���
���PvU1��\@��L�	 nd^vtP�
�z������E�#�u� ��
��R�F�4���O�oM�+&K?-m0�������D��`�+	|D�G�[�W�j�����������?OL�
/�ea&3qXӄQ����g��պo�m
�`Y�ʇ���d��Ѐ��Х5��ަ�z�v��Y;����Gs{d�WZ�S�>Q��+NȞ�ۉ�y��E��3{`�ܤ�C((H(�'w��m�F���o�g�yx�쨘�8RsTr���.��w)i�緫�Y~gy49E�d-���e���b��sAD�!����NE�˒5g�lt�g'y+šbJ�%��l[-A�h��c��Eq+p���ࠇ��M�%���Z�Ƽƭ-ڌI!�1�O����=}�7�4*9�9g]E,�DsB�܅]�j��x]���գ�*��,�фͪ["j
�ݼ[0䍄��% ����e�U�����(y�Ca��}u��d�j�z�㕣�W�*�ItEAI��g��{-�1x���x�<W��S�`n8Ԋ��?�����x���b�G|B�3�e�1+�Ƽ��(ac�WWWlH��E�V+�}<��̉����Ao�FnF�W���q�-��`�<-�u�sfb�&��{/��8�8
$���c���"��8����C5U{�;`�\d�!-�࿱�Ԇ��p��<���w��ߓqR�t��C܅�y*�UC� i
���.�?;C�D��3]*���ګ\�����;0��!L-�u.�ir{�g"�U��ڋ2�n'B������g�
8�c�'*;F����{-�JY
I8T�	$�I$�����ɼ��J5����N�]��x�� »�밷;x�m���T� ��u�7n��OF�n��y���ݦ��
E�v$sy�n�c���F���ͷ;e��s7��ױ�������y����:�1�4󝣐�����z{#ݍ�kXO�����:�Z�Yꎯ\��?���۶�sM�(�y�&|����5�ajyz�]�d��f����!��ˋ��rM��Udڏ��\��������;m|�U�^�=WsW��n��J]ư��n~wxV*������D�s}�0V�~a�{g�@�<��,�JNj��$j��=$�ʥK�)�M<��e���a��p�\-v^����2�p����4e]�b��+R�����\���'��w��+��j��x��z�Z)�Z� �RqT��`},hf��Hd���ڦ̼�F.��.�fЮj|��7��]�������[f��kq�0��B��a(S/�/g�$�i�󜟅�v*��(�Nܧ��"L��=���+�Քjv��}Pz�ǔ�u�?N�j�2��@h!����\`2%�FBIȫ�����*�V0�$���������Zl���-O������tϞU_5��݋�����7ңM�<Kl7��x˶�3�m�������e����+8`yf�x]R�@S�I��6ےMt�@�����Y��`��ͷ
���{�'E]U֟��C�Am��|!F�Y��;%�=�>�^@�$2>��:�[#�#�	r^$~�Wח�����=�t7��C�0�E3`�h)������Jl{-=��Bׄ�"����Ċ���g������qM�W���sKS�!���$n�ڌŬv�8�X#��EQ�[�r�����-�g9�Mn��fEe|�����P\L��QP�S�X�Hv��~���c��2>ď����3^�j��vyᗺ�C���P5\�5�Y�w=�L��D�"f'}�����m��$rR��{V��(�8d��WK�O�����JWC��-�Z٧�_Z����/N�b"Ȁ�B�K�$�n>��Yf��=�0z�/q�ӧ�R�P㼅��Wa {*�w�ΐ3��x~�3M�H���zǺic���wj��خ��)q'���ӆ9mv��/Y�v��\�p���U%�.�ڛ�?���6�k
;�i���+�܋�Aw[ƾ�ڳ�0�Fv���2�Q	1f�O\c�,x�;�_h����%'�7R=��d��2)�iP��z a�w�c�t+�ڌ݂��� a�G�^�[���0��n���^8g��=�"��!m�bΑ������Mo��%�,KŊ���-Lq¢��0��Ԯ��m�������:_�)�b�ԵW`���x��Ӳ�D�yY��u,5����\��Դpf&�}�QߜZ��`��Y�A��}z`Q�Co����Q��8�#�$���{gɏY����F�5��?wJ�@Zh�V�}Y}q\��?3�#*���ݵZ~�Ofdz}eg����N7N�����o��5�C2��c�V^)�.�yyѳ�Oֹ<�](x�K�:�>���F����M�'5��ʏ�߷~��nX�w����Y�"◩ճl{D#�,�g�������i:{=�Sљ��54��{�F	s;�����$�����Z�!�t�����	��i�~c�?�g�`���<<�h��I���Ŏ�ȼU޾���aļȩlk��<+��m��t���p���\�E6��ȗ�;,�͒�"W�j�m�����~��#?5�5��H���(����u�O�߰)my�pB��%�O���,�-yi��OÞ��ۋ���ke}L�Q1�V~�~o�w��G��Q���ƣEdP��叙�pV�<���:����W�}>�d'��Ņ���7j0Xu(f:�nuz����^�0�I����Ne��Ϟ����Ћ��Y<�k �%>���LR!}���Da�.wͶ�2�E
N8�aEd*�%���E���u�ޮ?@���_���eأ�;htO`+,Q�n�:u覊�H���0���ĥ�-~�g�����;��n�HD��e{:��u�q)��<�g�lSۆ*k�v6a�R���Fx�)!"�Oig�dn�`'1�M���E�e����-�CD���zC���T�+��6��*�9\ ���AW�OxT�I�֘[26Ym�$x,B0�.���+����GMv0#����+`�0������Y�U7��'����]w��\���H�@�%D�n8���P+v2z9�8���$V/���@e��Dnۼ�x9DpRT��q���H��b�#!2��J����hg����ƣ�X��#f���GjhZ�1	+yP~�~dWut�Y�C���ӻ�����'P�v�����m�(���3܆�e�#���N*�R���_���]������f��p�9[��a�LwK����-6~r�P���K�
7	�U!󓠾�=�'��z^��\M扲૲��N�e鎞?7q�l+�UK[({Q3�VXK>�/2�ݟ,G�'���$�#2:��>i�;�M��v��X�1�PD�ŷ�n�{r�#Ʋ��4t&��ϒv�I�����\�����A�^(Ƽl�]�����죱�vt�kvrjt��k��D�^7M=mQ�$��\L�m����؜݁8^�d�O6�*�Kb�Ktgϝ�ǰ㊋>�vs��f9{��{T��ax�f�t⽝��=v�v���,����r�;��ź�ϵ���l)�e�r�5Ƀ^ۢ6�q�e��������0-�f�L���6{�5����AI~�]}}O#뵤?ver��r�'��lsu�U��ڮ8/in�?콌�Ta�b!8�pV�d�V)����pK	w�qER͹ح"���]Yt�����ퟕ��48l��k����>U�̯-�Z�k�?�8���Î;��!�ز=2�V�GhT~}/�|qE�f7g�:�x?VI�@ggX�$�'����ZT��<C
�̎)j2cm8�a��.x�^����F��W�4vЈB{�ѡV��Le�=���.*�bg���Zo��-ac�0������쀨�.n#���J��j�v��Q���o+3Qn6}}�]SǸ�͉g�������4��d�����.n�]�Fʁ�d�(�n�u{n��&⚇�ZN뛱�#��2Yx��D��p�b6�qD���(���Q}2q�]V�3����P;4F#
R���*T԰Nu����24�]�2��$�/�a��VB&�rIp74�澇K!�]|�
�jYC�5傮*���\�t��>{����J}��< Ol��@�`�ݭ�7�{ض�U;��kzK���P�v�I�Q'�:�p������� cEwz�lψB����Ax�1�ԽZ��f.�m%щ��i59��8.dlVw�q{}�r�nV��j�jc4�*υt��Ɔ���D�px�|?)TC�Sn9�=���k�<-���'�x�q��I�oP�G����+d#d�}0�~<|�\�%I�kj9����K��n0Ѐ�ӂ�˶5��>�¾�8��4,���-:�`�;j��hUWu4�>�����Y�C�����VW�����ߟp���QO*��wk=cl=v\�z$�{g���{����u��3�v�L�[��+��Y�y}����?Y��U��"q\�`��6�{^P������g�D���q���B�P7+��A����
i�B)H|:鍊]�w��x�(����'5���?l<��.�ۺc�3���5:Yx��}ʰ����'ϡ�W�����E��J2�i���DK�W`�jq8�~�q��p�6�Os�S��$E޼�
�ת�S^Ǹ�x��֍dx��p��Sb�ԍ&-�Hf险���6�Q�����,9��1�,��=z�ԫ���sM��qyOT�Md�8�3�Ck��Kq$�rE��ט-�+�#�NWx�����]!�V���/n�Ռ�aa)z;f�O4�^�վ�T2qޮ��U!���ϒ%-�2L2D�f����!ϳ�"�����}��*m\�������ݸj�}�s��J�7�����,�����"ݬ}Z�@���P���ED�!�<�c�*��_E��t6�a��:������,u�@��R�"8��k�T1+'�O��s��8�B��f�eR6�
u[���>�;�M��采+���������q�cG�y3[*g����p&P�O��Sc���Pf`ü31U��r>��l���Nqȱ�@��R�o(,����/U��#��CE�D?o��#�w���	�(���_[q�yzi�(�|��xtۙD��E#~�st�!��*�B��#28�M��W��6�������ߝ��(\(ZA7�;�Z6T���s�W�x�C���n'��*�����[ZM3r34�!��r/f���(���K�G�m��U7�}�7+٘�Y�'zM�a�=��}�0
ǹ^��I��C!�fIe�0�~z�e����N���.���7��Lb�����f��pB�G�5T���#�[
���*��PAC&$5�d��b�x�\�wh�_2��IָR��L�#1A$���������F��Y��)!�}�PәR���r˧9[s8���usפf�D��/B�ă]�[.H�.8h{�>Y�O��P�B̙^`�+��r�o�����{Ok���FkW�l+����q��q%�|�� �?vEE'�&`��܍H�}�vK��Rw����TDl��y{]�t�l��*k0�����\�6m��0����n�񾧱Y�Æ�Љ���E8Kq֛�"�9�2c,A��1�Y�(�.`��͋c�kQ�9�ak��3v�5W߆e����"쯓���.OƢ((�9����� ��ZvX��ٞ��>�%��;F��]�}B�هM�<���k*
��;a��^�'���S���:�߻V}%ڔ��X�eu�>�X�ԃv'g33H;ܥ��7�k�u��!ń�.�TK�o�u+�B3�:�9B���+��a=Ӗ�T"���Պ񨤺��}�i��r�n��C��{���%>dRZ�P$�n���0�	ťj�GIYe�W������M�jo,C��onj�U5�(ђF�k�0o.'��C����tOL�gM�d�@�P��Q_"�`��po0͌Z�ʫ�#W��βЧ�o��rٚ�sٷ0u����M�@�;&�Y獳]W���4��ރ�̖���D\B�
y@�PA��s[ Ζ��Gk��0R�7�$����!)r<����j�G�������5�v�e��ɘ���p>�ٳ�҃�-��I��pOl�aw�OXA��]	,�JJɘ3#�NXDghY.�.<������Pn$����on�Ϸ�f79mtMز��h�[��Sx���B����Ujʱ�p2����>��Ѻ��kufyTW�A��#U-��!F��Y��ږ[)�&�\�hb��*vg[+p��*�v�$})��A�a3�I1�vi�����h��<��z����a2�(�VwC�khY׻.�b���N��rγ�+R����\3��*M�ou慝Ȟ��������^*�譎����l�* #N�Z�:N��E8of"����k7R����{��(��(��p%��%���$�v�zn.^^�yp��%t�˸��w�����?�fڛ�*ʵK�����S,uu����UUUUUUUUUUUUU�]�N�%���v�6^5ζ���f�8��:�Fk������muׇ���!�6���w'<Y�1�]� ��5�ktU��6t����x���X��ͥ��skq�Jvv���r:6�	�[;���u�óAr���9��6ݸ�F^��ָ_d�gٗC���n�y�z�s����5eQ*�3�&�i�u!kv8�e�I��n��+���[X׵��)��<��'c�=�[��ͧ��ye5��)�f�[u���vj;:�*��bVְk��řݹ�S��tps��nkr�1�p����>i��'\u��6⎞ۭ�Cz�!�p۹�瓕�ݍ��������y�<5�F�l�ō���׈���s�<�vC��zM�qv�t��C�{omRv�΂�:m˸.�1 u�}��;����xzr�>Pn�u��ㅵ�����c��m�s�%�>{1��<��;m;!ϘL�5����C�t�I�0�o]v�ʚ;[��'}���1N88���yxq��q^Җ��z4�d�:�tqG���w��H\m�]kp����p�V�r�����A�wln���&�+�:޲�f�n4�D��:����^���9��gb��\w�\�vh�t��ckDg���Un�&�1���iғ N�i���q&K����v��^mǇFq���=��%�����ޏ ��.���1�y^�3�68-�u�=�3�m�+,ϮT7S�u�u�n���]�3x���s��<���.xK�!scO)��F��K��8z��Y��x��m��y��v3�g��ьn��8e-۳8����ݒez�8ź:�j׎=��
�����-�𯮝u����7	�(��j��x�����9��`�}s��U��a�7X�+�W%�p-�M;@HC�g�(�]:��5�,J��J�7@����p)���4���>-s���ֲ���hA�z����dy�4�qsyf
�٪�Y��pt�S�[n���шŊ���#F3��D�l������v��8�ht��Z��VIdأ�r'h��c�sn�ŲtZ[�qm�ێ��!\x�$�ܳ^xm�FWL�퓋]�����%ƈHq��V�덷�d˶��sv�^%S�m\Y7
<ultb�*t�v�lu�]ȤaV��ێs���J�^}��������z���k�1�����b���a��5�9�^{f:]�Z�n͸�eǤ����I��"ɥ�+!�.�rΙ����;�b�EZ���RR[��z6�iC��A���L�p����pԓ���"e&�86mO�����q���=d�}��dƴ�t�i�`U�(h2t���춎���6�Q�)���#fr��9�@�"�%�a�Xɺ���{��W�Y���}:��1kz��'��N�2�[)=�k��W��%���g}J@���RJv�̜1��l3m���:�j�M��4VB��":����r���ZkGe���[��{�`���f�,��|�l�8��a�,��.�Ǜq�D3%ej#,5�/y^5�����g=�ˮ�u�G�e�.�����e�U��3!)$ς0B��e7�c"Lk���S4k���,<LU�	0��6�ȿ�N)$'�ю�yn�5�)�nno��P�B��l��}��,�u��_DC�0�h��!ӹ��ƙ�{�פM�,6͆Tȓ���ԋ�0;^�����f>D��vU�yt܏0O� �s�Gu�j٦ӽ��Y6IZlY��)`�*�Q��o�v^UaHomac/Xʻ��C}�m��绷-�;��-,mS�cD�N���zM&��,"<G<Yr���L�[wZS3Kb�%�\���ź*��	�r�8�VY"���Z�#"Y����*8Mͬ�����7܃��]���w��)BB2X()��Ծ׷���}����"�}�����)���`���wc��u���g�����/��� ֎_5r�O0_G�EG��{
(��E1�ikU�41�9�
�{�Ø�[�8P������._h��ʮ�%+ҏ�m����l��z�!FdX�Ϡi��`�)��v�<������; <�:g�%,c����Q��$]��?��j��J�y}^T+�ߚ�fQ��ˋ��t�\W�>�U�Usz��4�7b��G&�Zl��C�v�O����Ee]{�w��HOhc@{S�ё������W	��^҇�o��P+CM�d�����ї�Gn(�ݳ���,�a��5\j����t�h�ʔ���zD9E�zı2���)=�T$D��
��u=V�f��7�$;������ƕV��RN����`���h��0�vt���gJ	%�`�D�Nˆ��r�|��4�f(+o5PhtQ��ٱ3:�e�C�+Ec�f�Θs�uss9�ٷ`�ٙsg�ْ!
�!m�S^j�������E�l�iܮEظ��v^t�7�������V{�-W�}~���%!N�{���>B8ܟ��>�=����bŌ4:��C��{j�غ����dV�E
"S�(n��OW��2��}��+��r�W>{[��%�i����Y�u��{D�`RAM̺�/uA��;��k?x���k>B�(�ۂ��hC�,�LĨg�mXR�����@�����ZSztY p�/>���S���WPe����oMv.��"q�H���1�l�7����繊���۟S��YW�<�(j�w�`���.{K�ܻ�����E��R��t!|���G�Y�X��;K��꼛bv�,�u`��&�X�o�h�9��I���I�u�j�]3�欁�z���E�	��^ML9�w�˽ߝeA�ŃG�@���*�F��5um�mRR�ۮ������}gǱ@l�������QD��Ў@�!\������G�K�]�Y�t	c�������9��%g��H>齴6v�~~�<�@�_:�	C���pu�X��P�F9��Z��,���:o\��W'�n�f��y�ӡz.31]��l�X�x�u%�yC��b^��D�o|�{5���
�<�?.��r{�գ^|��AxL�b�� }�����-��o�=༞U���b� ����X�:��������`0�Ox��M���W����,�Ngi��8�PF�H��4�6<�(�Nܢ��N�!�׼=��݀�G�o.tC��k�^v�y}N�D�>�6��__�-�IA�&}�{���8J��6��g��.�S/��#{�RC�����^�P�Ʈhۻ�k���Q�z�]�0X�%�s˨��B�*3B8peUnGs멡���a��W�~洏D��hn������,�>�5d]���`¨@�3���l���l+�f�QuAl�c�ݡ��r�A��z���\W70���̳��z��Mô����?G��0���=�[o\HI$�I#���wmW9�h�#5�:&�z�Y��݇��uו��.���!�s��tm�n-���U�ː�@�*��ڡ��u�]tfh��4:y�Fw�;'��,ug�ۧ���67v9��e˱��N1�� �o]8�/�jb�3�ssxNGm�n�B&㳎l[^�1mEGFx�v�خF��u���Q^v�K�⶧G�3�eh�p����<S���ڛ%
�m�qn�4=�I����^��3�X�<��|�����Wk7s�g�oϻ���Qz�`���<����)#�#��C��^�J�!����A�#�����A�
n���w0��-=��԰�mY�}h,�/��M1[N��v�n�m'k�ki��q���j!Bh�D�(�B����Gۃ�T�_�~�EKj�zf��֏{^�X=;�z�	�1u��̺����"�+}�kw>��RW�I"1�H��b��#1�[QW@��{osyX�-Q��`4��ü��U��^���ע���ǪF��0�7L7�1uB��fd��(���	�)��>��W6;4Z�u��NVl΄x�=U-��i�DY[����`.��҈Ŏ�g���$Ԙ�W��@��mǛ��x�uOeBۃ�6�3�D�����r��qX+i���ߏ߯��L7�l���X��`Q�*>���uE�j�w*WH|��'�e��N�����NJ	��Oz�ߋ���xh�|�6b�����n\���fRa���zi��a��z���tf��%���[4H���ے霋D�ȵ1*��U�,=:�:#nI��H�ԋu�wr��<�B~���9����OS��E�	�xf���O�j<bBȍ��)�/n�ۛyPZ��kjab4�>51l��އm���uI��Den{�Qna�P�Y�+��|ZBB�-��\^�3���o�givi��k}���=W��kw��:���?u]q�S�4�b���[N ��"���mM��3y�����#�	�I|�x�����U�t�Ai��w\��󽼪��۠t�'��� �㝬�m������&�B��8��%���h�z�80��ƃ������L��v;'t�z�N���م����<�J27�<�����2!�u`���4I�2������+{=���ס���k���pV�7���zGf�݁V�,��ה2�j�D�꾐��4�n���&鏎5��y癀����a!q8s��W]u��ԕ�
�c���ߓ���´e�n��{M>���q!殈ڟL��Y��+	rRН>VH]�uB@4�,��\a���[n/��Bz Q��~^5/���y�Y�$�w�Z�;���N�Im�d)Ĝ�8�t�=W��3��ݖ���JCs�)�=��gY�dV��W.�9�:�퇥�����lt(r�D�FKR4c�G�R�s�:�h�>��������½�����$]�E��׾�c��]�9T�L����������ÈO��zz,ЧS�p�����k��N6'5K�֞� iE�JJ4`2A{f���U��~�C��ڤ�믬e�f!V�g��}ᤌ�H��y�o}���zQ��i�F��6��G}�W���ǽ��۔i�}Ǽ}��C�W�:�Ղ��/�^�`�X�wޮ�6�ȋ�_0�Ήf&�m���)�O���ۈ[�}�OX�9�zjt�:Q�o-��-R>"E��M�|�^e�)"t�rh����(�#���k���1�jGp�gei��{�Վ�cktV�x?P|�YF�_���v2����o��y}��Y��cPJ"��0��jysm�f�ؔ�ٵq�$6���	��gW!����uG��v!nԲvy�z���=s�7Ɓ\�w��n7 ɍ�Gǆ?T��:&r˾Vs\�r}Pv��T!�O��{���)y㙦��YU�ʹo�jЂ�_.�lak]8�;�z�&��s[��oS#�6���N��Wf0��������:�۷x9�K�׷%���K����	}�W��8��[
*�6��#��7���+S�}I�G�f�i����n��9���!�8���ލ�ֽE3����5:�?�N��+���5��k���<<��C�Q,7�.�t�b���*�+�3n����{�.��OZ�]�c��*s.>Cldl��)V��]N�(����!�E7�l����c�=Ao�Ԋ�Q�a^>yx�fҪ��9rq�qhd>Q'>��ὂ�n_��f]�����!6a-$������>�*_���V�����2�����|���wwI�}��偺�Ζ�iй�A�fr�G�c楤�&u
�dZK�C̑���[�/�n?���xJ^�Mnx��iCL�j����Y�s׮�J��R� ��Ȓ�$�I�����^J����{x�/W$C��Qt�׭�X��p�peٮ����.KO:�s��K�n�]<;�wI��{��,s�wnc��.�eqێ4�����8��G����ڻ7^�kl�q�#m����^4�7gn�U������ڄ�O0Jv}4˳�aۍ�O7���x瘧r��n������s�O;��� �C]�:^nj�n���F���:j����Dj�^�U������hg�_���o���kz#ș��V��lt�4����S܎��1tT���M=��R�mIR̶�rbl�%� 0�/�w�;�ot>�~�8��8+���"���,ʑ��Xy������?L`pX�#x�r�=��H��iG6a�Y�����øӮ��޲(NO�����fv8(���;ە���}����B9z6��4��[3�d��fD���yeѾ��/y=4a�-L;�(ro?Yb

�U���a��~�,�2%!1�"rM���z�¶������*
^�fe���m����S�{���4OL��즱_"�߅nlm5=��o|�)n��l9{��,��_l��Ƃ�qi���6͞ ���K�#�}ge۔��]�Mnf�{\�=�<�<z"��{	��L�����˸����k����Y�Li�d� h0"��w���N��B˯Z��Px)���k��%�=�^ܔ�7����9b63�e;�T�1̱hT����o�wI<J��vM	#�������^|F��9�l����*^_N �:A��n��fj�XއEGG6���;��i�P��a.Eb�W�k�OL�_a�+��z�ج���1o��z�ќ��g
��U�p��YHw�0@���������U���A|�oc��w�㳶����'R4Y�6}�&8)�2w\.���I^Y����f��&��o�K�9�ڒI�3s`�w��T�r�Jg���1NV��	�w�"0���>��*#!�׹��������Z��Ɲv�b!�Zy����N�Ahă͍�GG3�i-���tb��:8�wwjxoK���%z�9��`���W;nYyX��מ�ۗ�yW1�o�kʾ�XE���"�,���8b*�Xع.&���"6+��&C�;�qv��ܼn�7"����gS�}7�t���)���eh�k�s�!-7�7e���n�V	2�;$���48��Uk����tZ�FFj��u%m:ޱ��A����{�;�yn)&`�Ƚ�o֊ܺ�w������E��K�0�>�x.	tgNq�h#~�����0�ϡ����]�`��p�N.���6�5��c4V���GC�j��d��]H*_�c�.@u���uP:���
��/�U�z��`a�{��!��Z�6¼�j��rA�+��Kْ8,i�W�譣�i귍��}+�4�jW7+T�9ݪGj��i���iG7lp�^�+a�ŜX�0� ���[ܑ���ekT*����b����+v�(�.����s N0�tV���.�A�y��ie01Ȑ��M��-unK�lX����Fe���or���W�ȇ�h{�6��.=z��o*�ˈ��&f�*IN�q��z
�!��9[����_^m-4�f�:9cc�7���o��&c�\��!���^)`�W']��Yk
�Hza�좞��-�)��N(뵩S�2�M�9���iÇ]�:�/��56s��P���ouR�9�0M<)e��2�r�=v�,��M��,�ԺW+�W�DB�C�Ķop\��.f�v[Ca�V�aW�sm�e���T�S@\5th���E�!T&�#Y��2�^�޳�kۤ#�r��Zq.8;kk�9�G�gvs�b��/�e�޷�q�Ə�4園�e>�ٷ|m�Ma�_>ԵR�H7���5�����O��V�)悢�<�P+�v�T/�0��Z�7�3i��lVL��Xt�fz� 2�|fUv��k�/-����)B1A��l����9�o�c��=l����e�a��t�Rg�γ�q^ٻ�9�N�r��|=��}��Gb���G>�G2o�#��9V��bXW�X���V�B���|v�)λ�9��W)��/�`��kT�m�E��wգ��hЁ�C��T����7Y��mà�7���az{C��5�r��2TN6D��$i'|0���;�멹j�)l��c1<��w9��${�q�=�;JWw�;��0�]X�$�	Q.EckS��t��Z�;�n�"Ϫ\�j^uLa����]�����9n7{j�W��[3=Xya#ѹ>���n=��_�⩜q�j�u�%�^ty{׀��U�ʛщ:.��r����
��fl�-%:��iF�pg�0d�`���������V��w���ॎ7�v]���/arMU��U��ٙ�O9&��\���ۇ/u�O;� ��F���}��OE��pc�i�-�[��W;j^@x9�
��
7ﳵ�f�<"T�������#Qȍ��D{�bܜsUQ͗��܏:c�r˅7����_0s�y�1J[�|��D��4}���۰`�ZVP(�&���Kl!�x��i=9�ZMW]vy5�G:�K�757M��f5$����[�~̮y�Gz�K�Yp�i�Wj �r�K�>�u�^���u�}��YR����)�7*�7d�_]+���h�/js�o\+�}j�;��v�&��Z�)L�	���~r�SZ{ �\�qF�m2��7��X�ӻY�z�n�Vz�?m�.C�o�_a�6�)���g}}���XGu�"ǒB"��8㭹S/v��G��Jy��y�r$4=�;�!��~m���m���3:�Q�#��b{�ķI��p�n<�R���v�,a����J{W�%��^[\.��������4��G�&n�}���:	�x�>�w>��������l�)Ec�־6�]�u"�غ�zg<�p�۴��f..��!h�N:H�ydN�#�PR�UU'�\�	W����l�8�;����U�y��E�{D��{v䎺+��s��q⠱�ݒ<u��X��ѝv�	xT8��h�����&�<������tہi�C��wl2!rFemΛ�Ѯ/HIn�eN:��m���n.*6#S�֜��g+%z=׫�^3��]���ѝŞ#��+[v��R�w6 ���Y��u+�Dpn*�&�c��ݺ�n�n׈K��]����v�q� ��
#M�$�p�}S޼��*YAOo��AS~�'�R��&o��4VF�ۻ����u��ϳ	!s>���E�$�X�SЫ�꾘4���~��]/sbj�]]G]��}.��z�qΎ^�2�|Vv��W�.y�jS	(1"eI�ڻݰ�����o��)Z�̷�.� ��-ލL+�1\��{��ڹ����yޙU���إ��7#S�p8cp�2X��=y���vg�q�f�����Y�Q����X���؍+��wTi�'v�<������ǯ4jT��S�rou�eS3�����%x�^7陝�!��Ty�)k��Xf{���۽�y,Z��żM�&����	_(pM��/<LiGp6�=XN�D�p�Z�iX�l�E�!���F��e�{j�yN�����&W&|$��y�^G�W��'��tx-�o�����wn_��p��'Kw7�z�ˋC��A�q�u*e�-�;oIGi�{ϸ- �����MKAfʌt�X"��������eL�|@�+�ʵ���ׁ~�5k��=fAl9|p�>Fu���s�5��`�o�5`��Ʃ��Z��~���+�CIUQ����(����n��v�{7L^��7����a����%���ՅۜE�����<uĄ̒"�L���{@2�m�˩�Ô�s���r���0�=��p�+�ɹ�k���K��[]��.�H�y-�1�IJ
��Ӭ��,.�د\Y���nK��9RR���f|I����8�܊�:jޱo�a<�ZRQ��`���d�v՝p��6v2]��Q��^T�m�;U�������$��9
�E�}U�z��o�w7���Ι�F)�]���ܳϻ�<����i�k��VJ����PH�9�n��tVWMC���ony��Z�6�ݫ_Ǹ��J��ռ_�2�}X�6�JI�L@����1:C�ݴ�.Ǖ9ײ��͑y�N ���B�k*3o�b{z��2��V�Ɂ��!����9wJ�R�v��1Fx�t1'�xYv4d[z* r�]�YW���{\���.�k�y\e��
��ڽe�dȻ��c�=�nJ���f-�������D_��o�ow=���X*����E�N~�O8��2��}��J*F$qW�m������[���4��8m�۝��z���6�-B���?R�&��lpE��̫��OF���!-����"�Rk�d#v��.���ג�2jQ�f�זy�]rD���ǯ�զr�����ux�ҵ��]�xu���^��9����l�:�3z���`舡m9$��{��Qgf*�s�H������}�1�����\)Hy(-���`Wݜ:��(�V�!vFQ��P�D���Y��2�[�}�E���R��7k��Tg�Hf�5��+g|�������U������󩗐'e�q$�;:�<�J�r0�y���"��O[��w���4�#�g32rywL������`��s�7H��ki�����6��՛0e%O����N�1vK�zY6/u=e��,��
̥�J��-�"۪&��{�gVK�5Զ�j	F8T-�u����*�U���K8�y�MY�﬉����d1!�k���o@-�ә��F�P��#����v��Ϯ���m�v����sՒ�A���(c	?�І�Q��qɛ�?a�֜�0����9ł�n�]O,��Zb\�΍[�e�M��6�,(F
+>�"�r8ⱏٕ��n���Y�����6�p�D�Iߤ/�]{�5����U��֕'�Cܦ�Ӟ��D�9jH��0Bd&�I1��gX��v�.'�jU/(����L�OZ�W]�og:�ijua��w��
Gt�3���!ͭ��<	�ܞ�bnl�u
�.��v��YșxƊ�әku�uS6%k�?8�
�<k�nU;s�G�rd�NP0�q���0�]߻%٣dB�9v�����ƤPۗl������_��,�z�R��/k��T�w֦d|_�=\��چ-�n�j#A�ª��yjwXO��~�����3�͢uDY�8G�
ڽν�IL^�p|٭�[�2=��L'd���l9$�H1,�lܽ�K*]u�\���Q���p]��[v�n8&��F���`0�Wp��ןv�i��T�;�u� ͛��
�����@��p�y𡤔6��zwdö��G�ݍ��O���ܜj������{-���zv	�ί��w���Qc��	�=&�7�q�S��yݵ��8�gr3˺���T��7�n�v�8��gY�������×�n��xz�]%nK��ۋ��Z�\K���E��ƈЭ�������g�Mu��9����0���әr��6V_ZS�6�F��Xh��b�т����g5Q����SK������ev��L��U[�g�qy���Vuom�����A/9C�٢�#I�6�87y߷=P����Z�:��}��T�j?gwK�(p����/��P��-�K�:�z�}4+���@�
9+b�%�}�sv�����Jg�9gK�^*���5a뤴��ɣ�uo���s��R^��}#��L��4�c��n6QʿT��©�`e���^Ct��<���T^ygұ��YX&Į�_Z�W��Ei�iB��!6���A̙��M�F3������$��-kn��6$���Y�,zz������t_��j�*������f��F����^�j{�?\��`fH�nH���d#~�ڂ�#�7_{�����z��K/���Wox�g(Xb�S�X7�(�Z�J'��{[j_M��9Ǆ��=5�B�%��p�<����+�u��I�)�z��Lo]�f߷�i��M<t����(���*FڒIxcgQ�߽��)����|-̓i{ۻR!��m@��V���U�'���Z:Y��U�ĤFF�j7 �{�7U������ʻ�|}e�+����y%c����e�3r�&�����)�A)�'R	 �v-��Nw���B�d�G7�#xcZ[�egy�Q\�*G8�	o;�]�,@xG갍w�ţR&�E9m�h��$;E{t��øX���<�OnV�>^%CD��N	�l�Q@�m������b[�i`��V����ʒ���nw�"�v!ҁn1(���7"�'*�S���4����n9��y�����K�p��z �K3���w���5S��엱�o���Jh�vٹG3����!ʅ����z�������P�U�^W���6o�^�1qU��̮�Ք��Ҳ��ƃ���mM;G�~i�>Ꞙ6������[��e�2��#�f��9�=~n�7ME'��؁C>)��NC����O{}!{iԗ�Y�1��T���n������M��v�*�6�w���)�x�Ģ�
�L�d������d�����/O�F�~��~�H�~[٧ЌZ#���n�=�Nw��8��\-��pWeI�)l�2��
x�6�g�e�rmuݽ�q��^���g�j��$	�&�D�p�{iuY��Ć��9{n��&W#�ǘ9-��������]�~;v��p<���9	*(1��5�B����0O��x���q��9z���חW��ȫ<q��^{�`��b���W=<��KFTL�30����1�����qg'9�M!<���;�Ʒ�#R��ۤe���9/�cc�	2F(�͓*n��x�W��z��d~u��ʝHa��NA�f�sY��.�-�|�����Fh�Ҧ��c�5�����Cp�W��_S��u�
1:ZqL�3t��fM�a������
�������y��s*ŜZ>JED@�������e
�-S��R�Ԇ˯yg�T��գ�h&�Eg����s2&�{�n�i�ԩ�Ѩ�P�b�Ą���y�����g��WgY74N�c��tA΅�n��P��H��g��e�M�-݆���s��>�{Omo�^L9���T�~�!�Ŷ�@�QF��V-�����X0��"�wq�`|�48Qm5o�ѕ)����	Q�N��	� 5)�L2�5#L%$�����Wԅ��
���*9����W�t�:l�8筍�StZc8�ud�e�Q��C������Ӟ�v���U���M�h��J�@�
��֪��]O`|6�v��=�p-���H7{��k�+�K{��*<�S.�n��&��d{VrR�,�3���ڼ	/�s��X��[h>����V��J ͘�$�AF�lhvs�pE�Jů��Qj�4{����f��ײ���v�j�-�Gyξ$��z��$:�nY��Wʬ�pL�O=3Tʖ�74rVkp;�ne>�]]tuֽ��w�F�B�J�7^m B+˷s"��g]��qI��f�qY�~�f`����vE��z��K]8���/�U����Ca?���þ�i���-�Hl�f��lۭ�� �vA�:Ӽp�W�N�P��Ԙ�9�����yO�{�F{^nE*��j��+�Wv������3����!u�b��[�R������ʌ
��l5f��,6�u���(R���fd���d��}Z��Ĝ�:V��r�wQ74v�ō;��?M�l?��ӵ^<��1,mY6Q4N`7��%w���?e�Z���ه|^E/)�s��n���6�T{f�\wԅ�-�+n�)�S��P�&7&M���[�N�G����+j�\�$��~��a�n0�6������q����2�T�Y��.v1'`�͜E�`�3��ʸ(�E��ڏ6���G�Z_��oN��T���c���Q���[�����W%�󦄪Wkx6�;L�-Ǔr�ǭk�Cs�2�v.3:���9����=XG9}���Kw;�&M�+�6�.��cb�Vl�{��	�aP�Ni�f�D@�g]�-s:%���6J-K�t��U�hD�A��&]>����&k��;ñ��bc�/F5�-P�~��^5Ȓ��L�##nJ����U��S3Rr�+UlGi��������������NW�U��;����>h��/k�����ۙ�Qp����/k�0�t�&ے�Om�;UҾwh���ड़WT;t��ѳ�/e�{G'����N�sI���kt廣8�;7lm���S�v�ܛ&�x��.s�#\��:��m̸�5��ʂ/Vg��Ƚ��뛰m�5cd9]�Jk@c���-������I=���a�c������ݽ���C=�mYT���H�{ct� Sfk�`����rd����;�]k<��j�4Z�m�v�cr�����婆��;�ʝ���b�,ɒ�\�@��[���'m˭ۮ7 GE]�����s�ƫx�n���&�f�Y�f�Fx��6���{7n.�m��{u�n'\�gllnmq�oC�pS��5���p[b�R{Vn�'Fu�ݺ�ۋ�/cK�AWV�c-���]�,�9딏mU/5�3b���r\��c�r�6�K��g��^�O�gT6�e�۶(3��A�\���ے��\�ܬh�Uk�=�4�ט���΃�xV���\)%�	���xxy	x��s�G�Y���� )�D�;�(7k�lyzm��vn�;�� �ۥ6����NǶcB��k�����;w70����,uï���ӧ���v�U�S�^�<�9"ñ��n(۩�b1�p�tN��Z^�7�U����)�VeyG݂��q{wG:;rĜ���������x5�U�1��vێ���X�nս�S�Y�m������xw/CM�{u�;v����o���z��	��;$�c����{7;p�I��c�����f98ѷ����͚#�.�����x����n;��;̽m�w�\�tY6��̼��Y����:e�W1�����y�(۴[�-պ9�Mn}�aN�����H��c�������M���=ONzM����l�e�q��7F�rz�y�]gd�Ĥ7k��Z�]��{9nc�)���h�h�.�/�����]yv�	-*Ҽ�U:�"�����3��f�w*cRka�>X�sf�l�%,Yɮ��	�1v�w�h�v}�ݟ=��]��;��,���<����0c���N
s����g'b���cgY��ף��ړ�9є�:痕�h%�2��۫Wg�jwa��Eu�U��9��b{���x�UT�.-�q�qwM�/��n�HW�4��Y8�c�y�Y{��6��u��[=#�:V0۷�u����d�hW[������`���$�a�Qk�݅��%��)ȶ}�q�s�߉ܕ8�[Է�>�2�v{�����ΰ�^m�:]�f�H>�I�I�2<�:��|��Lr�ѷ͇5!���&����L	co��~Y}WY����ް�m;�w�el��I&��%������
}h�?#�l���H��ٔw�������o�;��4��w����
4�NĎ/h5w3hS��c[!��_y��4 �r�fg<�e?X�5�1k��y�Ї��UI]�D��R�[v|.�JL����U��dy�5�y�k7�:�p&b�ݗ�u�����v�(�����{�;s:ϯ�yA*!��#zX��.l73���dΝU�V��8��k�����<i�g[l��;n�S?��˜��r�>��;E}Z)�5���:kR��e{gm�6�bo�^�(Gi �|�1�ÒJƲd��y�f8]s:���7W'L\+����(�~��7G
�� �Dgpk7oV,7r��U���Řq�G�$d��YHR�l�|�p��u*�dI�u�Ec��N�T����G�S���[��^�q��-81̳�̿z�^�0^��T�'Xi�5HFV
x(�ynol�p���zn�س)ۚ=�qH�,8#*I�����m�ޕoմ��N�iyDE�-�R��*I[RvM5�}���k�%S_gS�7�HbmA�mt��y�..wu���Sy�9;nNj\�I�%�뱖u�5��{�r(c����G�C��iqחi���qÙ��zPu��ҹ*1��.�3�dw_��}����n���N�ޡ�w�0W�zH�u�˵�k��Ղ�a"�Ƀn
.F�޹��G,Wx����7>`�1@\��d�>�{��n1�R$7��7��`�=(��ޙ�v��.��.�f]��%��[���M�E7
%!n,���.F�׃qح������8H/̫9�<��WvT��z�7&]�sa$ƚ:�vr����'��Y�Ѫ�޼�����N]��U�d4O�7����,���{Z���~�I�j����q9ǁ�ǫ�pHw�g{r����齸�l�\�r���g��S(�U7ω�^�}s>�>��Ԉ.}2(��Lۋq��咫.�+w�����=�o��"�{.V��o������m�:ۖ�óm��MH�W25�[Q�ظ�^n��/n��6�ۺvڱ��rOc�\-�K4�q��䃽z2y�f�^άjԇ���Χ]I��&�zl����G����{[�D�7�\�� ���DD'#J'��h_q޸���7�Xޱ;/��5��U��6gyפN`x����s���(�E��p�fՂ��b5 0��V<m�ݯuK�L�����S)U�[[���E�U7��a�a�Ciz���ofA�V5�?ҙ4�t�rI<��5�𳊂c�_�^��2DCo����T���:�:�����<�!�7^~�j�=Qo��f�^�
�����%��ZZ-	�7J�����u,�H��>&��޵գ�W���,�����F����$O��!A��پ�ylЧ�d�Wdu��3e�gk{�<���D���6G�9E3�M,�RhCs{��K�D܄�`�0���$�9�۲ou��^8��j諪5�u��lVs�n���0�y�`�~
&W'$�{��[t�]tQ��4ԣ�q<	9<�I��<��V�.q�H�1H�koMݾ���f3�w��s���U��}0ml�����y�����*z�秭1��вC1D[.I6�Mۨ�?i^~|[ƽ�%���sDX�EJ׽��e�U���"ئu�r ���$ƌ�^�(��8��oy�B���o��٥-��
�v:-�e�<���Y��Z�s6WH�lH)I�V�a�쐽���N�sv�M���pk2���>�c�F�W.F�Ç�R�8����g��E�֍�6��J�Lj|M�7JZ����^�.�֫�g\;�g<�7����{�NL�f"��#�3-f7u�F���Բ$�XwG��k0)檪N�s�ͧML�Ѭ��{xs�C�ۛ�<�\�xˇ�����HM�}��Z��t����ӷH�.GO�ՠV����o]v��㧕z���]��I���[��۝�N4��v�ۣaНk��R��;:���۝���IMǖ�cu�//*qέ��i�텍��k���Z'��g��RTSӟ ��z��Zφ㛧��a�v8L��q�����[��-/m��V��9�	��wm��8�7\�g������s:{�\*}w�ʑ�;+}6�ݸ�)�{{�v����ݲ�{͛�uϪ���y%�!��#FdI(l����S9�'��\ǒ��n�p'ٳ[3�x<V�g����g8nQ������R"$N:��ɍ�RM�nW�zKߡ��d�����h]�$6jzc����7��RӒ����8�d���\l���q�Y1(��5����D���ꫳ��܂L��&�ωێ�\�Cys<��S-^��}]ٰ�pMU�{F�#��8X���љ�:E�YhF�������TP��;�����㧴�L,sj��������-C�:w �1�s� ���ݡ𽄔���WR�Yss�_n�:B�����h����#�d8��8��9����&ק��_����|G���(Dѹn��򚚬��ɾ���u�#�i�&�%���c��ˋ�
[�]�TK��%2���	}^�Y��^Fv;��!��3yIf��S2Ƞu��*�طk��~y�<3�*�U�Q�0��֭!œ1Ր�(m�[����i
f��jz��J���:�}��~Ά�@��&ӑrΣ�9B"j�Z�洼��Ǟ��x�	���\��7ز���{�\Y���&95	0�A�d6�����+�׻)(w1�jꠃP�_Jս�10�d=�O(-��:���߯7i�e\>�ӆ~-�
��RI����َ�/�/b���o��ة؛"��k]k)q~ p>�eMY�n���䘗xW<i���8�iinz�6D��)<��tD�nr�W��3�7�c/P��u��J6��$^�t������F{=���F�,��H�F+t7K�^�٫pP�4s5��h�)m��ʑ�,�B�("&A���ܖ�^1��q��B��ٝ�wY$�|k�fT��A�m�^�~yy���k_1;e���. h5
7C�]�=���js�(�q��A�]=��A)[P��S~*��X�6�BmgB~�#�M�e�56��;��;��wh�o������PKI��Yç�M�7(��M����Zm���a@�RG�-���*��K�����ݡ�����{T	�鐄��=7|�C\�u��E@�ÒD�V�(߰nmKdOG'���Go'>��
�{H��wV�P��l7������ϨU�^:=Hm�2>�2N�TM����]��s�l���W4.uч5��7'd�AD!(�	Ar�4\r%$w7����f�jk"�r��ݢ��^�3��L;S�9Ӱ3:3k�]�.�ʦ.82ZrO��6 Q�k�!��{n�M�97��mD��b��*�`GC�4�\��Qw���A��^;�Q���ܫ+����q4��0ؑɯr�}G�E�7k��:\^����w)xe�{u�k��c�-��
��� LRre��qcr���tj4mosZ�M��n���O�A����N�)�r�t����tF��L�Oi���sn�����ޮ��2�ը��P���]X��$-!c4ö�ٵ+y����v���ݙL~]w}Xv;Q�S���5(��𭱹�֦	��8�!���7�j�� [����6�vj��J���1�7��|exO�}��#�^��M�z�DC8�8[�rй�i졊&�6�[d8�[�n�5B@�F@Ё6be��ޭ�+ݗ1V;���:������צh�»�fe��[�i�N���&[��I�9E�P�7q�C3��}v�2q�#έ�V�o91iˆѹ��gb]O3�.�us�߫�B��,ےA�!�q����W�K���S�٤n��-�Y��=ȏ3���w�8Ƞ�P������F0@��(Ԑ暙��h�yN"��
5{����ɱ��vMC �ߺ���G,6���w�^jn���9{��)�*}p�p�߻+�X�r�s��Z������鞭Ӑ��vI��]<��w�F��x1������dp���UԳ�y.F�&����0VJ��	�z��Y󝜍�R����t��^;bn�վ��Z�8�,4K�IP�vq�v^q��~�������wkW/Z@�)sv��n�on��ӡ.kpy
@tbsz��d⚚4��v��G��]��:�«=n.y����od���`�&�j��v9��ݞ��x<�B�z�8M��,�g�el� M�H��N�����u�FgF����ܣ0{�q&��1�ݬz��cQ�#<�G������#��4'��Mm��\��mI�n7�.���C��v��y;�ܼۤ�menb��`l]��5���U�~xE��*4*+�O���1Fvb���~���)ݞ�wԦӪ�Wu{]�Z�%MFL*I{+z�����N+��/��h9^����n����c\��uhڮ}"��6��]e$x�S�jI�s��u�Y��>Ge����{�A~�ρ�
d����4Y�vCx�D��K�R����n7��m��]�׋he���h��{����{��d�}%{ſ�o3p����;�u��e�\�-��E�m��쐓�Z�o�^�}�6��ƞ-��g:��+��O(��yk��5�7�����7my{cM����-:S0T�b��qv������jy=���q�����a8��H=�p�֟�Mį���ŗ��.�]�i�Y~ώ'G!c�n�gE��uz��=��-E$/���N9��_U�W�\:�F����%]����1'�M׮xlv���w˴!|��XM\��.r�	tm�&Ø;:l�!,m^���3�4Vҝ!C����3�����D[tY�}Q3*��s���Ú�N��/v��]��!"̖��i�#�Z�u����.�[إ�O�z�ø����ʓ�y�p�w\���P�1VJ�@�-��I5�lBwc3��[�Z����O>�y�5D�����:�:L��;�UW�}�}�hz��"*E#n+���{�D��Rg�XƄ�M���7�b����OD�{�}��i:I�[n�[*�6���Ǿn3[�`E5��s�Ʈ3l����ێw��<��#�1]�d���8���P)�]ǥ��aZ�7��:��ኚ��ĈR�4$٦HfP������d�x��ȗĊ4�^�X�n��j��E�c΃�eY};�`3&�R�g.�����a��6YC٢r�!���꺽"o�ّ�aNI"�!zoF�s�Ţ��3�����]|��;���$�6]O]2�)�u��-l�U�aAvΤ�J%���D�0��e�`x���6��R�R�<��6�Same��&�"<��Ja�H]��ݞ�Q��]7�VP�1֮��:��u"�Z���w4R�x7)3@�4��x�q�2wqsV�k�J��/6:�mZ?:���e��y7;!|�mv��[���r�H;gK�3�^�Q�)B6�bŏ.�!-��NXs���L�poA�!Z^,ƺ��r��{��n�v��ţ��l��o2�L��&��EdV�i�aYl�)��fܡ�1Z�v�e��d+��M.�xp�;h�p�f��␉'_˫�.����\�W�;�|S�I�qn5;.�]j���1J8r�D��=�n9Xi�FprqNPų�ӱi��j%�[�nmd%cNR�}u���Gy������\E����Q'S*b�7���z^�[����U��tc�k)2��^o�v:���N^�կ�t�\���hI����"�'x�u�7fN�z�
͢n��1�7T��Ť���4.�7Y�lx�$]��=yt/fmm7� �Ys�L�k^#u	�C��;��4��-���UJbv%Ӽ�?i9�-e6���n7%�Mi9j2��r�wrY�z��ȕ��1�;���{���ӮZ��K"�mME1nf�wA05י{W����A�i�]������ �+r�c��
9N�Y�{3u��v��n���)���xܢu�n�]N�;k�e^^�u\�V���Y��{���������|�y�A�%�7��>�CD	(&�rA�nߎЙ�Q:��Θ���;��K �V��t�;ҳiht�g'�;�ଙו�\K�Ϥ��*��:~�J�s�b�����ݦ�l]�fE(�M��Ƿ�(��3���6ƈ�@�0�H$]a�-{
�Vvzܥ�Z�m)���OC�Yd!LHZ�3 m�y;�^��힧����8TpjC6�
��%���I�t~��[�:�m/T�B%p"�"u#�jӺs���GB�63��[^+s�eQ�-�=�d^ghrbו���љO���\}b-�1�E�	�G��=�za��us�@��羍��nz!�V�iiU;:��<���]�#��7���hq�Z\�1B�a��w�T=ּ���7/��B'��ι:&����y0�l	:�T=l���D
�!��x��;]E�a���¥�/ʐn��&������pMw�7�g�|`�u�V
wX�.��zݼ�,���DMC����w�p���I�UV����S�$���ND䨵lާN�zxh�K�1ږz�/_�QQ~}��n5��~�^l�^��E��9�kXya$Ӏ��D ѐ�~[.5�v�۬��F]�H����u��ļq��88oD�C�ӎ>�w���b�t3�s�4��x�[���c���@EQ�v]s�*fM���J�X�H=�� �n]]�֜�h�{ڻqY�+6�*�ì�4�![h����-vr�w�ݢx���*���w��^Ǹ"1���`���8/�C��f��gz�}���ކ�n�'�Y޵6>�=�k'�vv}5�jV���ڐ�7����W��e.�� dӜt˃H2nmp��ZsS�at�tS�N�DNS�|���vnx�DC�"AI&ἕ�;F;����������渐:����%�b�A���5���� ��p��\���p������ii��6D���X"q^MTK�!�'���ŝPR��Ý�9Z�i��z~�\��G����f�%��*����Tvt&q�tq�wv�z��u�M�q��-���\=��u�{�L&�.6!��L1�}���iz���=d��m���5]t��[�Yb�-tu��z��kMٰ���v�3���X{r����g&���e�^M�v����ryO�ٺN�"�qr�Guj��έ��s�sˮ��=یe�n�[������l/Z��-�ۮ��������Z���ۣhN��������qPѴ��6:#IӺ�J��a�=��z�4nDa�OEw%�[��K���u���Ta�N�[Ƨ�o6�\��G*Bʑ&\��RnM��Uެ��]X�(���S^�j��({����7��M:e�����wh�d���GBQB2[���)�t��)f�������2�$s�8���ث'+ܢ��>�<�a�4�28�V��o&�����@ۮV�m�}�!�CN�����n�T훇q-���^~�p8�S�M� �"h��L�zEL])��
��h��em?u#����SϾ�c{��+L��W�w�΁�_�~���`�rn1�Vku�*��0s�wj�	�yX�/1�tk�F�}���'����տ�[s6�ݗbaaF>����?��^f8!��F���+G�s��x��I"iș�4���{���6�V�_\�!�ez1��KÛ�C=�f�����+C4|ڠ��o8[���6淚�Ss�+B��tt�i��C�l�^��1��B�}4���sn��_{��[�9�u?K�,zn�u��{��1o{N��KC��&*N�rN>�y<�f~�]\��y�a~O��4�}{���-���G��VB��K�q�[Q8����z v��Zc&<��[���z��3̌�F*ü_���/���k{�,t���5�bgP�
M�* �.'re[���k�wW���k�	��x�o{�Q����L�=���P�Fl�EN���cAT\%��<;؜�-W6�ml���mَ���<��&�H�:���������Ԉ�aG�o���w]1�/"�ݣe���N�����k��[y�K��λ�O�]񑒡$82�wB�V?7��/p�>y)@B�Ն��^>�tY��z��W�>ٯ�\ݙ1[T�[��ĲY��p�$H�T&c�Q�7,>��|�s�G�u�l^�TG� �&�8ﾶWQ���E���Bd;i���.��cV�f����M�a���j�A�"�1��{����-�i��]�؜ŵ�~_��@�������lIqI$��/�3�%S�"=�﶐�d�n:jtl_<�Ӻ�i
e�%� {�*�ʦL?xߨ��ua�(L7`�� �c�q۱����RI@�[A�ؘ��u�����6��?:��Y��*D3<�	�w����]�L�]�����9�&�l�˱�Ղ�Z^][HI���Q�võNI���[���I^�+zyݳaUwl�c��΁:�{�!ݽ�{Z���E�d_A78�hü�c���$D�aA�p�y�	���|U����,pp5y����Bΐ���ٕ57ޔ8�j��4�Ut;�8)pJH�&ۓU��Wq��6�v�~�~3X��Jk9�4�r�m=}�/a��_!I [K���a�zk��ou�v=��7�S6�3g���3�6��E�Cw�m�38�\���9ޢ�����]���5��ʸ1�i�=�-�������:�G�\�'w���������C��-ۓ����`/e�]t��Ì)Q	.&�1DT�X�9��:���K���PX�s��^����[[���t�^kw�!ب�=[�qB�V�(ԍ���$NƹfLmM�l���l��\����î-����r�!>#�	���o��]�cU>���[T<�8�c]͝�ɞ�fs�.�M��8�e�C��'�_`a��G��B�V�����^p܊��w`����s���\!���u�U�Ӯ��Z�o>�ݬ<}d1���Zbp1$,��p��Dz뷟�lmzlח���J�'Uجg���Uh��˨��G�W?9�'}j��j'�L�~I�N�nM�ՕR{N�..̊)�z��/��]]/��)�y�Τ��B��sO=��iľ����b7a�Zv+({�Pp����$����X:�E�&u�M���'�8`�"�hBk!oSԪ�_[��J�0�)o�h
��Ovj'ީ���
ݟ
^�ӛ%QX��F�Hׂ��rn��T��Y��p��ZĿ_��mVڇe��� F�yl���:WZ�����;Kҍ�ϵɱ\�9���f�8]�-�:޹9䁋��;����u��9�-�lܼlf7d(۟s�n�cI$��O4=�y�v�v�z�w�&8�Rc�N£s۫����`��s�n��|��l;p�m���c���OZ8,#8ݹA�3�=`�E�&�\a��ۻj�k��خ1U:��Q�����f�˳�R��3Ŵ���4k�����{Y&�K������6�"�2҄��rM��B���!?�~9R��+x�x=��x�:��#����U3����˺˱[�����C%3e��p�ۦ��yl�~|	|�N��,۽*橳wu_J�b�;��x�L��O�N{]+f�W�g�@�r��]�yسja����S�+�����(�;����y�k}T�y�Ka����.�>@�q����T��cYiy��y=f�a�d�e�j�;����4�<x��uy*�d쮳(��8��Dc��Ԃ�2lu��.�B�{˔5��6*�;!��yn�UA�{�v��0����p�[��F�K�z�N-
&�M�[h��B��c��ѹM=q3�t�u�Y�6�9���@�.�f8J�I"�&$&'��w�������ڟm��^����%"�n:�fm�|s��Vz_������&���IAfD�"�(3�i=�b���{����t ц_4t�au�ܽ��F�X�������9.�*ڍ82��sfYɿq*��#��O7A�v�om�U�ׂ�������Zx�o��\�\^����B�6�����<*k���V����IY��HLDq��v�n����L1�jklC�/x��!����TzȓUE�&�/��>u�<Q�*-���8E$
m�Х�}�W��R�\�ת|�[�w�������d; ��}�&����v�X.��"�����ơB S�|+�w���vgQ�aR��h��Jo|�Ͳ '��o�/�ɀ����E�M��J�3��P|�l3vw���c�;�3ۍ�-��V��s5\i;PЍ(�)0b�)v{�����xz��q7�)�LTDOr��Rv�6%�Re:����c/��.XkĄH��&(�sv��!����vI;����_z��s��4����v+���8U��� �{oM{�Gg[�H|�B������evW,Y"���u2�3"���Z�
��>�㜂�e��њ���ѝp;�lU�%u���Aר�lb�Ej�qq�Mu���̶r��m@D6¹������%��;LB��1���ۅ��߇��`;$�*�yt��?o_Z���q�zR�tm���<�zs��~��[{e���M�IƤ�=��ɪ���YƷV&�<�����զ-�>�\�u������+��wee�E綐�:Ǭ=0�j	�r�T@�pu�h�\�=�o��x��7#����\=�O��j' ��H�A�$U���v4��=9�i��;yM�b��Znm�d�^�3>ة�T	e	�d�d����9��KO�P��&�q֯�ק��y��6�%��*G4�M9���0*Y����8�8�P����rAq�v��엧s�6�PZ�2�nN���ҥ���3�?P���]&��:��MӬ��Ϋ���dw�6��"�f"H�(L�{��Q��9٭�6
�{{���ȫȜ=o�D�h�FM���:鉔�άI���dۺ6p�iܳS�W��х\��t��2��8�2��JǑ�V�yhFv��nr�5=��@
�9ͶT~���O��x"o�L�#&8��
�#��]�,��UZZ_7�֧�����Z57���	��4-��[x)	z{OW��|.��T �KeP&�1�S���\�$�Ӻ�-&��7mZ��-ص�WgfQ����{��f�fv�j�n���4�+���]���c�5F��q�֎�����c�8diFLN-�l��>��c���g��h�~`�F�Hn^��r+�P5<N=���}~��}di~9��x��%$��	$�� ��Yu�2�Ng�*mqg��mC26�g�o:GZ��-�9�[b֪�[�11$�-�Eȶ�fAc0���]��X��<�w���j^GK��d���E�9�e���9�s-T��N�3�j�,||�1��("7y����j���>��=�ޗ���ٰu�ڡP̠�x�^�X+�U6�������%�ď�װ�u�{P;�2\U���겠]x���g��c^"��qBHP�X����$b+0�bnnV؏k�uE�t:-M�W;��aor�,�������,��=�M1��#����kB[Im'&�����+����K%��1ǲ���#x�"������R��.l���
�1eS���qMɈ}�(X&�Iu�V(���x
�tRҧX��#hV��]V��' ��VѧiP��('�?���o0R�}\�#yי��2�еiM����-�)�ӝ�%�h݉.*E6oRν�J�D.j���8���U�,�!�Rb)�P�I�2��]�v���ܨ8�RGٳ(oNK�Ƚ�7%^��m�튰��=xE�A�Tz����T2v�=�^�n�g���E%B	ʕ�%�w7H��ր�P�����N���峒�(��z]^/��/:�a��yOr�Ԥ��0Zk����kY�=�IE��m)2y�P��WJKY�n2a[�cjT��&n�c2�6�����ei{0�x�jm�N�{����W���x�']J�@
r��8����z�c93feN�$��;ɲ� �'R�E�}x�7�u�>]wfIN�R#)Z
��FN2�s�Ug��J�t��\ů�̥�:�H_E���LZ��C/�2*�V��ȏ�H~o�vP�}gp �^f��o:�Z�dᱧ�E��\Z�A3�V˗����r��fm��ݾ쌰�MOv�7X�BEZ���5V��:݅P��4jP�ػ�y��[Vϝ�&���2��UJd�
��UF5UUUUUUUUUUUUW!:C�����nQ�zx`��usne�]�]6�&���U���t�M��OH�{Z
�6�X9��88�%����9��8�}��^����*D�v7;q&�3��^ۛ/�������#ۙ�3v�����c.c+�q������cv��.C8^�N�'e�l����(7�h�}r����Kk�٭��y�*��V�v�nE6�{�v�����s��\���h��v���cs�f�xG=Z����=���q�S�wW\�4�R�������E��I���g�t/O��R�]yDwY�q�(hn�������v����.N���z����H;h�B��;r �����̍���]\v{<�W��%�\��Z���=�g/V!�xn��1Q����t�^wE�k�lu��f�;�ot!h6v�r�V'���wlfr�ԥ��\�\�����}������G8�5]���v�ۉ���u��U��:6��q��ZSu�g��t����m����X���3�h'�s�c�u���oC�Z�w�ͮ{. ���<�yj��WM� ��nՒ(�qWf{�v8�^9C�����{�z9�ζ;gl��
Ä�'����Բ.�c��k��ݭ�r�&���s�n�ms�Vz�>+l���:`�6�\v�7[r��uڔ�؛v�=��v����<vJt�:^�tD!����ɸ-r=z� ���2�3�t����vw\���弆��:��<��`�9W�'7k��n�f�g�3�C�gc�s��Y��t���c�+����}��<<��of��_a�{\��V�m/!��=dC�����]��\�k\�<��Gu�%�s^.�j��M���ݬ.Wa��lfչ=���]�ͷG�O���k�l�ݴ!��v�>��G�h�@+=99��kn���n�rv�I۵�$�9'm��A&��<\��ݜ�t���ۜ�az�ۭ���U�!��)��]ms��˫4��a.�ע�xB�׷:	��UP�vU�p&��/<I�;��;�����ՖTu�ͺ3��a3��u\�P����[]���}�&��7�]�:�A�z��s�:�}2і��xsŧ��l�j:VΙx�qY��z��r�u��v�"N�V��������flܐ�a���u�۴/G�kw#׬�{q���'خw]OB��-�ݨ�r��答p�h�4�Ѥ.��w<ŵ��Ӹ�z���'z�T���d!z�θI͘��慙J [�D�O�?L,��ú���fc�g3�jQ)���b�������i>Pp������ю;������k���h!�ļ���,d�	�i;�U����ӻ���o&��~�Z֥m��9#)��M�8�mS�:�����𲊫��>+�df��f7=��=X�0m���B	*E�QD���ڱ�R�pD%�n��M䳣��d깻�t�`�ܽ@����KԽ��w��Sj��Xa���
7Ns2*=ҹeKn��E�q�`�-��5�Z���6����:(�B
����9��L{���aշ�v� BBT�G��''8���	s�h���Nx��9�o^8jN��X\�'�R�������_���m��W/��N�i]�HΈ���ہP�#�{���=z�+9��I6c�a��bl�'_�In����X��H�]ݼ��Ӷ��0C���R�q�4WkV;�b]4�S��g.gZ��"��c4[�y�v��-mνk���mн��ݹS;�����k%\�_J�p:�u׀���n�<o���_��Ip4����I+���Y���!��92�/�Q�X�e�)�g2�úٮkpN�F��]:��f3e���/m�F��번u)�nd��u��6:.��ˈ O�@�.���V�a�1˚ͻA�����j� ��0�?o����M7��!�7�=�xه��H�^��5z��s�����cH���2�]�Y)s{K���S���=��;kvi?IA�ds��7��[羳��G�-��Ŏ4��hl��FHmt�<�[��8��z�k��nKd�S;utI��
d?��ڂ���-�nw���0�v��zUץ�ݑ<�!�`ًB����V)��C/�x�x��m� i)�N���Y�~��8d2|��($1203��E��a�S��_n+so'�ڋ"��h������~��?W���^��ȣ�8���W���uʲ�q����d�dׅ�լ�բ�K�(̌��)7F�8F�VtS�>�Z�1�����߱���l����� �:��/�-5a�[���ǃ�J�0& Pf]�zq�p�8�Ֆ�ݩX�Ti_X�m������p��	b��s�W�G�3������#O�?=�GJ2H�A����4�j�oϭ����ԉh����q`��f�Փ��@n�6x��B��vj �*�"^�>������͚6������L��Ւ����`�YUE��gEW�\"��}�zt_��#�s�؉��d�y��}�B8HQ���4;\l��7uGz�E0Che�G��Zh����]´�I͔�sд<9zBp��t�u6t<�.qwh��Ϲ�.su�C ���	���%#�8~�8�lU�=ό�|j�Z����Y����O�R�(?_]�[6�#x6�2z�D@�]x�b�~�5����}��	�q�jAw"�ϵ3dI��z_����J�VKE��>u�*��(�$�/�ǯp�CW�聥�9O�xk9F^\d�����@��I2~}g�\�_�q��4��>H�(�~���:~Vl�9ᣄA_��a�����OƢ�.c<~v���'��Y�E����꼘.�'�s�~���iakM��hƢ&E}��#{{T�C/FD��hi�Nn>�g�[�A��E�f���zi��*�7\)�q��@�/�۔��e�{�10]�N����K��ڛ��3y�;�����6��'��ՠT�9�*�9;x�wJ���C��5���3{�/��߫�l��$�(b���ib��E��!4��%mW���^Li�%9ş@���k�Gz~��������H�d\���|j�a���������~�oz��ǺK��DӚs�(�r��v6��]u�j��.��c&�nԜ�v�s�QmB|�q���'��b՞#�&t�^��t4��mnPÚ�mWy͋'����V�&	4;��V+&㏷��Fn�y������}~�+ZxM<�ӑ��91�������*J��Hob�<xx���,�/H�=�pTttϹ�/�6�����	6JZB7��o���Ѕ����s��@��nM���g��Ǫ4A������� �#M��1��������z"���X�<Q'�8�!"Ͻ����77~�g��"��4�txђ7��h@����ݞ7����Ց�h�x`�?���H)G2E���&�4�����ٟG�T$L��G�7�"N�B�"���B�ƐmL&B9����hf."��C�"����7� �|-B���a�7[d����
D�f�N��Q�'e
#O�W�A��{�I�����7���:E��",��D�N�P��8B��=7�*Mid{�(���&�EZ�w�~�����qi�b���L�r��o3�q�٥�Z�2�iW&��w�)�0��O����t|�Wx��T��U����9{P�`���ӛUc�ް�8.�:�[lm�t�uv�M]7=��{�qQ�몀B�.�V=nx��^�h����i�JNG��H���ۇ:L,EsѬj�_3=�k�0�n�癙p+v۽�7-�<�=� pm�OUӆ�{�����Z��Z�wSVԝ��l��Y���n��v�S	^͋z:�.��I����h��6匑1�y���e���댵ۘG\mD�p�s'Æ.�\�UU|�/�P�`��~}�4]/Υ�qa��^��2ɸq��<pd!ޫ�b3�����T�!�C:x����u�R�}�#�������"�gѨ�d�)ɯ����JYX�����jD��K��,��U�~B�W7�D�V.��Y�}�V'�Y��3�O�wƶr!�yfɘ�����7�.?.���0������������8���\:\�>��Pv%�v��a"5z����u
5��3�dI���͂E��Q��8���߫�ɔ-	�S5S@��<�4�V~VO����S���~ȡ�a�T/�ㄇ�>.7�����]x.)�잊�6�3y�5$_�z*͞"!|��8����4�p8p�$L��:�����$yw�h��cU�UW��wD״1��CO�6�S?`hO;�5k��?2]�}�~���� ���,0[պ8�����Mͧt=:6d	�����zy���k6�a7���ڱ�����s,�6ښ�������f	ӫ�����ЬG��p��b���0����!�N�s�@�ٱ�-|����G�Q ��)�^1q�	��b�ǅ�M��F-&ׂ-�$}*$�#3�Hx�d4#�Z��7O�!��Dѵ�x���G�4����"��(������{D��Z�"`_G&1�]�s���5����jאM���SM>��f�yq{�7ޏ���y|� �ͪ�(L�F���}�R,�9�մ�?ּ2$w��������Z�W�#؂:/�G�G�;��'�j��C_a�]��/�hQ
�_��蜕�HÓ�/�����<r��&�s���6���?{��W��211ȤT;�3DKGf��ҫ�V��7=2��4d��E��^b����E�$�B'=�/�E���G��T=A���5GOݧ�#?$G�P���p��J4܂��r,��"nLg���《:k�#�1���=|�G���c-W�hQ����߱X�p�DB�:}�j��m
�+֣O��Y��A��S �bbA��N��m�'.�;�C�R����z�ޏH3�c[��F���\8=��D�����ET�y��Oj҈�t2h��zh3�����s��b�ު�����G#�>�����~��H�LaG�K�R��`�N7n*t�V~�GG�Yߩ����f|����"�{)��}��qJrSש7HW�z��G�C?Y�y^�L�}���!��"��px�a��*TR:����.�+k��W[xG�l�=�g�AV���������8�+�)�9�̾�Ev�%/n�f�j�F�z� $�P���NQr�"�]�>޵ݹ��]ˮG>��*��.Y{���J?���2A��`�Er3~Y��5	|(Pdf��}� ��$L	J2b&M�ŵE�v�>��|�8<��a��N�$o!`᧱^�u��J�.J�6��}�١��PCH3��}�
^�|zm�Bψ��YgO�#|~	D(*DB�&&%X|��!����=������@���΍����?Y'����Z���9�2)�O�ڽ��+O���dY�)�_��`��f]9{B]�Io X��O΢!l\�pd��7\�nA7pzcr��݈���"�2�n7a�������!����ٰʤ'��}gQ9����(a������*���4�ݷm�o���|���W<�2Q���Z~��I~h����l��.I,h8Y�i�D=���M��`��jE�dP(6D�˸P��o�#���X
,�ú�6h����d��&~ȎmMTcŬ�0�@�p�k\@��F�^�w߮����'�z�5��"�I�'��/�_:�#ݹ�/rUv��8^/��4)�"��3E��Nw>w��F��َs:F��='�QN|�jF��Ac���<:X�νe����t{F>��?n4c�����A����~V2�|���5BT��\�G/��ؓn�w�.{�ь#��,L�^�c�x#��Ѷ
�nU�ƕ<�.��)��8-�(�xJ7���y:�l?�#�� ��|����F�9+��F�#H8�$D⯳ɚ?o*��o�ȡ��If=��Rv���f�ƽ���m_רQt�;hO�z����2ܱv���9,�W*��ε�򛂷���z$K*ĆB�����"�����.6�Wn�rl!�cNֶ��:�O����Wh�j�T�U|�˱|	�R&��}][i���,�޿E	���	�8��^����\cD�!.��Q}��H!�#>��Qu�x��CD��M�Q^����bO�nHk��۸X�4����f�Z;�4�g����z}°��E�d�]���=�&pz���(����~8Y	A�98�SQm�����N��J�G����(AR,xƬ��K8P+�^�7�"O�5ȳ�C2=�A{���B^��1��u�IY��(�	~W�����7���oa/ǂ*&�6��[ʝ?R�FBj��<���^驪�فdC4��f�W���B��+������t��C���~�g/������4<x�hH,сk���ԉِJr0�p����uar���L�\�����SQ��t�e>޲��.�p�J�)�|p�JP'5��´��$F�0x�/E�ߵ���
�����c��>�q?Ə�*��Y���-I���tj��ì��
��ջ��0u��G^��K��1��{QV�cV@�$m�0R��UUUgv����m�,�ݪ�Wj�ż�Yy<�v{{9�ўێn7]U��T׍���a��u�f7[���k���k���Y�y�N�[��h}�c.;r��x^���Վ�vG���kv��v5�`Nu�y������I�kq��u[�[�M���l+��{O>��|^��W;�m��[a72.ǻY�n�6�\�u����9�֧���H͵v뭱���6g�U�Y͓�������mt��v�|�et��H�4�.6܃���P/5h _�!����ծk��+(���nG'�g-(_s���f���Q	^�G��\O$gS�G����͕�M��e�Nq�˵��ɘz*e7q�������m#ο?����[:�>�Ͼ��#os��]"Ν#*s���='�"ݹ��8�;�����:p���5`N��B���9��ߴ��J n7��,i�g�{����5��/��D�~�t����P�=�~��^�����ء�������z|�W�3�?��쬶��q�?�R������<B�D�/���B^�?��,�C�[KI�������#J<C���������f���{�7�Pb�a�|��&���#�!�q�f����2d#*J�SO0��$>���ŧ�����������ԉ����B���#$��,�p]zh]l28��D�L�E?��㗳熑j3��8�m����b۞�M�L\�k�`��pvlcjָ=\�ۚ-�w8+S۞" ���SlX5�W�v�>�g,�Z����Y���P�d"(�f�Np<{��/�����}�2�:-!��<\��d�K���R��)ܑ��p_�"�����k����I���X��fZj�d'!���]���n�#�fu��9d�a�+ي�j7�:�K�����P	Ӟ@��T��C�b"q;Ko��|E��"�B^{ʄ�Ν(�KbgR�3ƴ�A���ǯ_f��	��������Җ�dNF�rC�O�������ns�>4d�}JRS��b;�C8w֝x�u�/��R;s|(7q�P��aW��~���q�<���k�����Q�n�W�g�'����5�`�xY�d]'��hw/b�5��3ʽ�o�#)E�"}��B�`a���R}[���ޣ�s��k�dZ����'��Y�C���q��q�c�M�Dx���6�f{�}gV���Eq����E=,*sSB}��BT�d�P�{�P�=Y(2F��3^44�T��8Af�?du?��]X��������Bm�hǋ�1�p�2�����77����玈�9��L���i�'\l_�����-i٥(��v��m�|�B���Y�z}(vFq�����/۔�7`ĩG�)�y�
@��_�D-(�9RIc�BH����{�g��PqG���g�S4+�h3��>����L�?2"�>�ױP�_L���˝��L�2+�"KҊTM�����f��K�}S��:��͘j�Z5�1XI�!�w�M�T%�ߊ/q7��@cX���'m�C�p�EZ��N�ͮX�1�@��]g`,��n�4ۇ���u��%7T��F�`�7�즠<m���F�6+D�D;)ӍlQOb�@�GBˠ���j�r`���f%��6J*0��̖���3~����dΥ��0U5w�T�D4凵d-z�۠��Y�0�Ǖj��Q��׆�B��s'��`݌�p�ѝ5���I-œ�:\�xm�����ї��^��܁R')�y)jo�}��*���t'�CQZ�cRZ��7�ݖ�~�b�[�VCwS[&�d̍Q����`�5���z�3aӹ,��v���u���A�C���U�S�a�SsV�W�O���Y���2a��&�pS0�����IB�e=ڼaY2�1�{"���'mޚ�V�4ڲ&�jd8���"c�j��%a`�A��wJ.&�&���&�J�z����i��cE�(aJ���4�&R;�>8��E{ޔ(��%�����)�9U��Tt�y.��K���v̗�v(�j�^u�NU�ۙ�COi�x��r;����y��v�.���U�Pm�\��mnU�8��8�B�"�+�`i��&�������F��`���ʛ��Z���HZl�dRSn뚾�O6��^y6��{�m��p��Op`��Ԯ�*^OR>�F	uZ�q��xg���Ҫ�������Z�Y�{h^��1`ԕ��y�o�����ԯSۻ��2����F�*+�3���n�j�n����YQ��In����&ӱzn����x���r?E��$���܃#H��adu��#�Y�.4L%H�x�����LW�%�A#c�پ#QhY�>�B�b��8ɛZE���Oy�,|��p��1S�SG��%ec���:E!|����c5J�STܪSR��W���ɂ�>�}V�Y��l�W��9O�@t��W���n�2p�=;�*����L�y��lW�h���LCu-x�Q����m���d��0��븮�nj:vM]�C���c�k�3V�F����u	 !�q����̌?B7�w�d�9�6�/�w��b��tH"���y
�N���Ֆ�.1�F�GY_V��i~Q��2.�"��NB�))%J*2܂ǎ����i�j���<vg.�b�=C����z-ٻ$��I8�ꖄ83j��Q����ja[����eD�><̇y����˽8~�t�?�H�N$!���a�+4��f��Vk��o5�?V
��������G�N�Wz=A?���'�8�r
�0�@���J�3�}W��<kK2�J;�>�פˀ� �GN��g�F�=��?�~:/��W_ib�q�����U�ђQ���jH�>�c��Oϐ�!{>q���Le�"�r���Y�n�K�1��0�Yf�����>�:
��%�Iիr��:XR���J�tz�:��2.F�Ad�"x�
U*?UYvK��p�����|~�j��/�$�y�g���RG0h���6.�TDx�L�@~��p��I{���� �)04�jȥw��L}^D3��+m�u�z��i�0��!�[M2�뭰��N�upttv�swO�[�u3O爩��%�we�����e��Z�=���бT��"����tт+ޟM����U��1���
K�#�9������$�}N�)�^�())0��"f%PdQ�0�";��&��X��q[͞H���������s�H�N;|�ЩL�մ�#=��Z 䗜.���H�Y{>;���!h���`��0*f��!34��
���~�\=���`�J�W�I���_iDf:[���E�x�F�Q�M�g8FpN�.���<F����Fc�qI{���9"q�tq%8ۺ�%�=Y��Tol�ϰѣ�rp�hW�����~�g����;�CRDYZ���s� ��������0���ǈ䰋���FI�An��F|��f�m`��9�k�}�{��GP��!z�׷���0��F�کÞ��Cܴ��fD���;5di ��L�t�Dk}ٽ�J�BK+�[!J��ɳ��=xhvd��Ջ�*���8M�Ӽ�ݫ�'ؕ����ZhL�*W���+���D�A6$��ĒI$=�bO���[b�vݡ�S���z�u�@]���ݸ��k#�K�ݮj78��뛭�G�ӥ�:W��+[*�c��`���KYzEݺ�'B���]m]�ۭ�p�]<=�4o.��ܮ8��q�;sƿ��s���τ�LdSN�#��ஜ���7.�x�\%�Ѻ)�<v#nͱ�6Ic����w3p��u)u��G;�ٛp��;��pb��}���&��ȶNŹs�3mX�r�9Gt��x��u��v�;b3[K��D��%_��J�Z�5�����Az��@�l�&~��~�1b]߇�f�NE�d\���<D4�{�A�#EjT����Ĳ����E�0B 1!R����"�������<C���;���� ��*_G{E���z�qN	w�+�x����UT�<c=k&�ݨ)_Fw��G�!D��*0Ԓ���Wm��<�~���V��A�͑�Ȏ�� ���w�ƒc�\�m�3���1C��4�'��y��x�5
0�#���J8W�C9��N.PŠ�n�+��!���{O���Oof0�~��U�bf��I��ޛ��E��6}��	z{�Ϣ�[<�D�R8ɓ��~�)Y&)�(�)��\8-"m������G�i��e�t��t��;�v�Rq�����,0�����&�_G�~,�O� 0h���(�=��O�V![�
�j�.�2j�@uݛ�%�O��f �o�N�f6T�uu%ly�t7Ny�ލ.�����zض��j֙O��Ƹ�G�����
"������yX,�tJa��[Ӵ;E�L{3i�y��-�W���à��9jԊƏ$D��� �wo�����H��foh�WK�0��_�%iI����7���r��;�ǆW9��h������Nm���q�V�H��Qr)�`���
�ۅ� n��	�o
��'"��/�;���E���8�EhDF,"�I��@R8�M��ă���}�H����t�L�$ZH��k�ߌX������_�d�eU�`�!����y5HC@�$]��ME���X~�8d��˒'#�TF������]o~��� ��࿼t:F�f��~������er�(Ta��Q3�B��'���m�)�͋�E�=�u]�#[��p�QB�����}�<H����a�e	I>��S~��^����Y�ؑ��0N,O����9b�KC۱V�=y�d��Q�O)��,���9U��<.�2�6� `�T����ޚ^$�Ɏ2:�5-��b��φѝ�у�r����wET�ux_Â�����d�����XtْN��f���y{�`�z>dW/�L��i�60o��OZ���8A�4����zC�χ��_f�=S-��I�s�0/�m}ꬂ�	�\U
ç��>���hdNN��-&j��@�֑�HS��M�GM�g���*B��͊�5��v�Ͼ�����8ݑ�]���a	D�J���9*!u�d+�F��̐l���W�\M*�\|�UUq1�u�i{�7����%SY1�>l�d�o��OV^�\a;Gqɜ�ںp�sS9<���}���Ŵ�(h�4zom5I�_��Ya��Y����Ӎ�'�'�j����i�-}ͺ����>Hf(M�_q����yB�T�k��;�4G�lW�j���`֨"ҐS�y�("4(�"w�X�9P֊��a�F��������4��Iea�2?rL�D�(F�I"�J��*L:L�0`{����5����5+lW��>��v��`��lA_��A@�^��RnН(h�����y�_��]�Ս��̓2�<��m}�E��;��Z��W����u`3n��!@LyH��
ry�u��܇l��`�Ԇ�V���7欏�`'���p�x4�T��AO�tH���y��K����T�{UY�/#��塓t�A�"s<�.�dI�b������i�h�
1�Ð����?Qr���������~�'���+yq�_���T�>�}����-6i ]T�?}���ӧ�k��m��_u�B�ȭ��rV,c�{��4Sq2�i��Tp���o��dB�?��g=hQ�(8�@���U�hH�B�(t }&�f��~>&��
�]B��(q�!ڣ�jw�
��R �N�E�8%�����a�%Y�0�V���p27{=�0x��,!b�ˁV��:���J#J��]�c���hm`l�>� ����WR-^���DM?��Y���X�Eo�@obډ���fz�u�ZZݬ�����9^NN�
o����F�������ZE��im�?A���7��AV��Ĝ#�ࡥxL3d&�����)��$w�����0 ���{
��a��
_O���F�>�xm�H������H�����;�y�fG��� �w!�7v�6�ۮu��9���om��'+F�P���q�C	�e)��p�|�R��[�_6��2ȳ�q ��Rz߲*�5n~�z�_܂;1�Vo��${[�}3"�P�����n�"�^����� "$OD/�,�I���La��X�4X)4N�$w���ŧ�/p�M�)<lв�	X�s~/�p�klVE�}�Z5}~CH}w�H��曓gHw]��O�.�e��g��G��#QI�✁�NIC@�% u@jM�1g��'���|�e߷*ˌ��<�K=3 Y���}>�u@�K�_V!����^H�;L�������;꼛��Z��������a��$�&�R*�N�
��k3����S�=h9w�j�i�&:���2=W��2���Q���};<�y��ў�ώbwo�P�sq]�"=K�R����	&|Xp��.8�d����W�T�����Y�a"�r�4�����h~
�o���:_���~-,>?lC���j�D�#���8�o��s�J�'=J!Q*J4��a���M��9��Ğξ�i�djo\lw:�1у�E9�5Xo��%.�W}��d��p�DLͽKf5�4�4�]TȠ*��������c��n�p��<v���j3v�5�^��\�`ʼ�[`�x�T�Wf�J�ܦ3�7`"�,s���0m�"�8;74�c�`ꇳ���jt�F����!���ڋG$�Dl���<������;t��7��|v�c���n8�T���'��Q�Ҍ�ݥ��Fn;g�Q2�/�J�P���먕�ZM��:�'G[��Y��5v}s�n�`��k��׌U�طn�6��x)�;�<Vy�2����nhR�>?{��)���"�������jE>U?i�������a)�+HB_���>����ut+C5�aX�5Y,������M^��X0���~�Ǣl9����qɘ�63�"r�i���ɭ�r8��dߛ�U+|Es�G�u܋�Vl�ӊ�k���z���ڧ�XUk�LD�j #����b�M��9$��k�jb��c��L�M�1
fG$������П�������>TX(��D�Gu��ZD�.<�`��7�UY��ˀ�����7�"�L? ��L�ߋ�i�X������������URn��������w81����}�\_MT;�`������$	5��-���ǆ�dQ�A�>��\n}W��v{�y����@�E3�F�=ί_�+�G�ى��po����B�������\ض� a.>��3�k�}�r�|��Ą|jW�� �����- E�4�D{���t<|	�C�H:�����u�o�B�
����'(%�}�^�v�u=��p�t��᳘�l��((�n6"	��C����*"~K��h^]�f��H��j
�o�P�yV�bP�B�1v}���tGOk�B
�H��D��qn�gW ��! ��}��ND'N�IUFtB��mcʉ6Q��MX,���H�b�zī��m���vJNK�<�\�զ�Լc	�I���9-̷y�,Ҽӡ��nM�x�5r��p��X����`���g���,���ܴ�)qS(O?R��t�A�"<�K�roroD{dH�Gg�����b��G�>?:��uJ��@�)�
N��?e�_�Q$r�R&f���1���FA@ٳ�O��_vuP$�w��z#�UΞ�<H'Hw�ʘ2p�6���MdA'�=��f!�=J�U�N7�p�X�$�I9a�8~{%}���)�`vH�����h{���>W��;��r(X3��<�@�Y�W��>>��T�������G�[�� ���.�IPV�� ��#Q��m)Y>B�*i�9��X%n|�a���P�/n��T��zzIl��ڡ�0�Foe��&'��٪*D����D�;�xn�"�"�܊�&O=Ib�5%�!��~����v�����{;��Z^��Gm�Yu��Q�WZ��u���(njz�Xj~�[o�d��O�ߧ�֍KA��Z$�������d;�U91Kʂ�sދ�{����ެ��{�g1�]���8�����?8ʅ�d`�$�bUhP7(i�����L������Yx`�G�s_r@����X�Z��0��RJ�9���Nb)[E� �"}ލ��?���QکkҨp�̈i�����
B~��	�\�� �M�Jv���>�Y����*��s�U�����=�zo���6c��̬�jumq\l` fM�dxug_fII���^mZڲu�P�����Q�ö�|d:��9C+dn¼u}�C���ޫ堓�CdSA$�"@��1~�ERIi{#��{����Dp��.)X�Ć��,�3_����L{�YGV��^Y'
2QawV�!+0gِ�k�3��Y2Q���I^��~ɇ�J�i�ߢ��9 ChG$w}��n��P<�J�D�	D���������O�"��V-�F$/ǣ�/}���9Y|�";/���(F�:a��~�ZTGO�7&I#�'gۓu�o�/��{�Q�����~�:�w�ѝv��Rw�n�����5ԏa �"�W:��y�t��y�&�Q�W̩ph��Ң'�z2Yw���t���B�d�9}���6��~��}�kŋ�#�|�!gի�/�B1�|+�Y��tQ,�������J$EF'R�O����cd�����{�Ƞ�U�ҸN�Qz"� Q�=�̊X(̏J�Y#~��ر|�1S`����Y �<�`�3m��ԁ �'h�?�)%$!H�I7�Drymx�d�-��ٿ���[>���	��U�i�:�w�!A�}��qlO���g	�Z�k����/N�$�d]�V�mN?�+�!|��9a&U/�v���3�Z�<B'[�b��mt�`X�~��f��P�q����-��o������䁐���P1܇eY�&U�^t���ć�[�
K�����[��Oj��M=ʪ�{,�-'��q!	i��SM�2��yy^vy\Z(��.���s�8�Òi��SSOkfvgFt��@�(�:���AewF���Ӟ���7�T)���|`r�	.��.�:C�9��9/��a+������4y��E8x��ݽ᝾�V�����<��ě�\Q ���;��םS�ؕ�W3bې���4s�ue_G2`F�������+��$����W����U�]� ƍq�ZS�B{=jřn���Dl��.q�.�u��#���#s~�z�<I�}Wζ��{���LA���h�'�&�IH�QX��paj�'�"� �"<��m�x��42~{�"vot		��J�Dy��%=����}��-�0	�S�}�� ш�4`�5�f	�g��m�#R�k���[�lߗ�_��ٽ�_F �=��4�R�B%��$�$VX 蘭�ߖ{e;X Z���a�+�O��h�{��x+��R6f���h����x4�;Ϲ6�G�.���A��rӎ��¢D��}����A{v�
���֘G��~%�A�IN(Sp]��)���#�
o}�EE�)&�@��g�����;<;m8�L�߷r� �����9�p�U�y�\�<�Rp���9/W�z8^k ��o+��҉0��?pSJ'���ĸ$I���#���S�lF�ӳ*����vt��|Y�jQ��f�;֟;�g6�d)�F6xh��/}���cZ"D4��I;E}�YZ�� �H>eJA�H2T��R�)ҥ �R�*R�JA�R�mT����%JA�T��)�JA�R�l�H7*T�l"*4T�J����d�Md6ܒHu�~�A@����|��}���o� ���}�H�I_m�hU(�mn�PP�Uq�h�XIk
i��]md�%":�I��"��D�P�
]0��D��  �$���BH�EEJ�H	H�U$T���HUQR%IR��$�D�UE%�"�)
J)J��"�w��k�{ﾽ���ϐG�}���_)5���yye���O��yn�z�ky�mmc�J��s���m���y��ݻw�Ǽ�u�v�������x==�����=}�wm�v�r{5()Q|}H�)B�R�P|���l�|����WW���c`�X-a��q��<u������}��7@
�|��������n� /������R��d��f}�=}�=�v���)U�hI=�>�T��Е<}�x}yGi�=�a� }�}��
]w�p:� ���_s�E�������l�����g}������{�^�v��� ��c��Jp�@��-�QR�"���>����T����QG�}�m}˱�כ�WT��q����� /y�ꈾ�6��&��`t�nq���]:/}���}R��ރ��{�R��7p���Yy������E�r}�tj�P�*���>������H�d};m(g��=�z֚/,�0h�ԟE��t�K�o��#|zo{���}s@����Z {p>}�:��R�]�JO�}��5�: 
/��A�DEI6Ϡ��e4ӣw�Нm٧��m��D�L��������W͟ ������i�|�����ށ݀t}S>Ǿ���;>�4��g���JB�ٝ]�zQ���|_|EK�ׯ-�^�����}�= 
<����v��続�Kͻy�ϒI�M��f�:+�^���;�<��4o}��ʵ����E�|�(<��� �UN�UHQ-�>U
� �D�R��{��t��s��t�>�=���@>{YV����� �ٞ��A��m}�{ϻ���^����}�u�������[���������J=�n�>�UZ������J(T���h�� �*N���}����w�w0[��>�}]�����[�wvQ�aѦ{�������k�a�q��T��}�ﾹ�P	{��}�΀z����=��K�R�ݎ�D�}(�F��T���I(U	B*�������T���W6��;-�������k)yj�m}R�>'����f_ngw����I�·��=s[,u����}��wbyb�����ԕ_}}�{�zѭc�ϛ�i�҇�w�[G�:� �E?&T��hѣ@ �C&�@*�FI*UC a0  �?ɈIT��C@4    ��P
R�� �` LL�F5ObUEb     y(�i24�E2z�=M4������/�/�nI��[�\�v�i����-��z�zhz�_i紩������wwW����$��ww�t����Ӻwtd�I���wt����I:ww2O��/��^wO�����ww������'ww���;�wwt�����?7O�����tI���� t��I�$Ir$��"wbIv;�:$N��N��b���JN�:wS�;�:N�N�%:I�IIӤN��@�'t��N�t�t��S��t�;�t���;�t�I��9'IӺ$���$���wwwt��%'t��I$�N��:I'c����JwN�%$�$���%;��I��'t�N��Ғt�ԒrN�'$�wwtN��ӻ�bwN�N��t��;����D�'N�'wD�$���$��IӤ��:Rt��D��N�Ӻ$��;�wI�:t�N�I�u;�$����'I�$��I�;�:N���$��Iܝ:I�$��NN��w��ӱ;�'D����:rD�%;�&'LIҝ���t�I:��$��$�NIҝ�ҁ���ч5�w_�.�������<�o�������«���$���>��/�M�Qt�ǝ��e�du�������]1G�����<�L�ës���Q�6!z1�i��%����a3Ɉ�=�su�2���k&
 Rn,�jkWg��F�sq6�T+H�e6��gv���G����T�{�2{2J;��G�y]��Ms�_fw�n�O[e;����Cɉ:�<:t�$��$�t�$鬝'ON��Ѳt�y�=���>'�@+�����S!��1�ޖy=�h;#�K`й:���}W�`s�ѽ����f�ʹR�Ujm䱇�(6NUԸ�[9�>};�t�Р�o�=�t��L�J�Hr�E'	�_7�2ȳ�&��������6�ŕa~$�W+%�����Y{k�O��/,�Sv-.<n�]ͼ۱$2�fc��c̓���,͸�c%��y8�Dڨ�:�ko]e؂�%ۏP��GwV3�n����
��7�T�T���n��²&6�\��uڦ(*��)3��b-��gl��'��˹��i����WB�*��%�L��ø�v.Y}�MZ"�r��8UFr�T�S�_�.����q�k�V����T�*�Ԣ�Yzh��-�<��j�!Q8����t��.�@Jf�ҁѓl�^�B �˪��LU��r��F�P�)�
�(�q[*�����v���$f��;h¢R���W�
��l�YhK^8�݈w+s�s�L}���j��ҮS4�I� -��b�]��U��y)[��R����h��Ȝ��M����25˨ո���.��D*�ộM�"����ڨ
�p�E�}I�R��16�TԊ�5��%��qw.쾖N���z3]Z,�����sI�z�߿\)Qlu���@p�f@2�hG�\�}�����ƅf� �0nR���=��E3jk)K���d�Uv�?-��l��2N2:D��Q�"�u6aǨCv�J#Va�%��##F��� ~����d�����ݒ��V�+�5���[bܦeՓ�E��'r���S�4'J�^� ��	H�p_�cw.��:
�u��j�:4��6��7�w����%�q#RTl�,�L�����(fqv,�1t�
�Y*ؽ�$r���J��Q�4#��)6F���</���.���//'n�'�'Mc�;��f��j��A7���\��b�e��)�!��a�^J��X��7"�K�i����U�4XZJN�0�2��&�Dt����e���<Q�jLq�F��*҅�1��wF�Wa/��v0ց!�Yl9���b8�Q� VMǱ^5�	���H��&֗IP{Fg��&;T%d�Y�YQ<��&�&ݙ��j@�w�2b�b�֬e�5�QN%,�3Ru(Vˁ%�̨0�0D�[�C)���5҃F�����6n�Je�N�U75�v��Oi��異�w��}�����1�~���)�����ֆ�z�soiݛ�	��M��ˆ�(���s8�/�L³�c](���๦3�jeG��:�V:���ݚ��wyzi��A����v��A��%����+Nv[�_�;!j�����:��6�ux-M�n�,7�]�=��J�g��20�%��)-et:hZT��5�Ͱ��e
s!�{��ekՐ�Gidv#��s0=����s6�կa��H�.���!,-���Qj�7wb����ƆiW��ei��)�a�1e�u4������T�����!Xr}���_�
�LVՖ`���ƀ�32��w(����L�Gn�]_$�]7�1����,��y��5��?f���&�
�V��ڸ���}
Q�L��[�`*���ʂۙ���[����7wY�� hѣ+i�T1�lHia.M�H ��@ݽ4�E��޷72$��ǀ�i����b�<g L�� �5��ax��l�o6��I���y�F6/wQ�
n+�Sj�P�5Z��-z��mWt�&h�RkA��@]���=��AYx�t� �J�Q������ �,���܁^ ��إ����j���+af�f]=gh�Qn~�i�6#�i,V;5�j�~9z�	@e�̗��shem8�ıZ�Z���H-F�h���D�JΒPmT�����u���#��[[����#�ڈBJ��t˹�)�Au�m2i�.�恳@1F�OSٚ�lj�� ��F���]���^m�#e��	K �p�մ�:F���T�i����h��!U�U��6�t���yo6��B�fn��M���/^�i3wF���q�tnʷT���wv�6��kr�� у��aֺx[��ո�n�ХB�.�'D0)�{-�tUЀ8ԛV �%��2^kz�w���R�ȍL�7)�2J.��۠E*\w�Lw�5��Pk���_��r�T���ē3l�[$+bX�U͕t+ oMSl˟��7g�+fS,��	���%��jb9p1&S�ld����W���!x):���0��ͧw5\Tk.�� '.�լ��L�a��Zo��i���Y�k�^��(�Kq�Lڼ����3�"b~��2>��E����?U{��H�d.!��V��  B̎�]X�������Y�^I*���D|p�
W3.�m��8�a��"�ڷ!7x�~��j�:���hJ�R�hgG>ٔD�-dK��$�M��^�v�α�.�d�آ;��.�w��\QX��c��{o��%�`_g^J�9��:��:�U	�0,�Ǘ�����ձ!Sku%7�0b�U4��w��u�ͣ�1;&oUԴ���yH��,�g�;�ձk�K�����%l�o6U�uzV�Jl��.�fb���L�����:���9�H����.�E�@�J��,&��%ڂ���+��l���eo`���h⼶p>���t#�)ŭ8���E� �Y��^�:S�V�+*���W�gY�ğ��wF�g¨(.l����M'�Ŝv��^	 d��q��s�ۆ��1����:��/�Y�r�i,����*�1�Jku�*�*&B-��g/��g(K�d�2Qk1ٶ�Ԙ�ȝ%gV!������.B)��&���fۡ���b��s2��y.�Q��q]��2Ŗh�l���,"	5��R\]����2lcf�5$R��%Ӻ`9Պ��ya�Nfd��၌E��U�#��t�+�*��u�%wW u�(n�5�٬�B�PG�u�BR��m�Y3ىX05�J�5L��(�M	x�2�$`�ˑF�j�b�tE�S�zC�(�>m���{m]�CRyY�h[��u 
^a��&K��4�5@bN�h�{1;FK�8[TX����@�ܕ;�W7&bhm�4V�Se�$�ouk��7W�ygfX��q�{a�f�!M7M��k��v���v�������F5kR��i/��a�3/|r�Y}��(��!�H:�I\�蘐����*�e3�֚���E��(G@Z�
*�W��dbv2Ū�K�X��`S���a +m�ak;m泯KL�WhL��K��7�yrg�d�;d�(e�P�������yWy�N�Ljԟ�Vʟ���Ƨ^�T��1)���dwp�(�8���Bm(��Ʉ�Wf��� �ܚ�'��Xr��Z\UJl�qX������]e�j	��5� .T��,�R�Qr��̔�j9Yc2�;�����D؍�a��,*�wu����ױ���ȕV5s�jЌ����v�nD����ePt�e/FK MR�VDܭ�um�*fvL�r���L)\++�B�W���W�`}��~J|"�_Qf��`t�@	\��7�(Y*���da/�J��Y��5-�Dt]0T���γF�~)n��#21�DH:C��pP�d�]1�6Trޱx�R*H�\tX��x�Sb��[��Vc���0�C*#���֩u{�i��1m��tm�^˥}Ʒ&g�|K���A_�M��Yu��k�x��3,�V��z�0�+����Z̟���oT�e�Ž�3#�h]��ܬ�%��A5R�Q�y&F����SZ�g�D�w������tJ[t4-@%��Vi�U��Lwįh�]���U�4�>˵m4COs{�|��Kfuh8�ъV�B^H�̕�IyM4����˻̔@L*7t�j+�*��3kV��Ƹ�MGR{WGk��cr�����`ܧ}y\Z �ګl��F��6��JZq��0�n�ǀU��hG��
5�r0�F2���J�e3���]�%H)��b�.�\��x�̈Ʊ�$Q!���-�ܼ�%Ss�Ҍ$�� f\����Է*��Ym�q��`�G2�\32��S.ld�]cW�ME��"���neҜ��T۠Տ*ʆ�vM([)=h�&5�����AC�j�eK���隸�ҺIXC�"�EUd[pؕ��(�	�]��x���c���Ch�������0��J�]M�f�[z����j��kSPC,�{���?a���*Rrls	����d�?Xʺ�c�L�U�Y�*��˨ ���.�"&�����J�[��O�́:�4Drθ��K)�َ��wrm���zD��L[ѮJ�[��5�*�(lIw��:�Զ��D碥Zpj�AM����쌴���]j�{n���2TLg7nHn���o6PghIx
��ّiEm
69d�ٺ!')�`�R�X�W	�aFm7�v�b>��e(TZ?%�`x���z�
wc7lc�5m>�{7���.�/�Qт�p�v��C������CY��2 4��� 7��.��T��)u��&�ʛ���T�p���Y��QǷ!�k!ހ�]�v�%���n�b�!��w�Ù�,w� Y�����~�s,�����V��]��j�l�#p!
"@s����8����ʎ��Z2�N���L�����WVӦ�����V�˖XXl67�l�#yD���(��=sB�k����KmN�k\ރ�p}�-���7���V��F/#�W��~����R��9��;u������nci�n�v*M�,N�}pouFh;<�P4���Z��m��)��]�%6ٻ�atw���j�+�=�pN�-���5CC (������+�oxG[T'_F�E��"��Tԗt+�w�v���ʳ�S���pA�����uj�6�)}�"yNA��ΠĶPs��Qv�uK��6V�7��-]tۿڒsQm���녡�<�̳y#;jfwj� �G���n�����CNT�c|���vd���h��q<�l�6���Q�ާm��J��q�zsi��vV]� �=����B��橪�b:�
-�٫���*%l��H�c(�W�U�f-���lY���*�jI�ظ�]�s��s�6�_co�ww�[*%�L3 F7�W�:9֩{^��C�!�-Rl&�r�s;Yڄp��)� B���ՋW���YtV��(ԭ  �:�H��0
\(h���%�Gv!���L�nm@�/��"�AS��PU������e��^��i��F�Eܖ!0D�f]�s�@*3$���ต��[�W-ɭT��WKhT�l�t��s�[�S�e;3	;q��#���% �J����2���i��L�m��3'A��H��K��j�G\��0���'N��&���Q~ιo^���iL��ֶY�^Y�Լ���i��鳭i�e�Ѳ:>PR�w���S�gZS�e�O#��n8q�%^-�YWi�h+�3�ƌu�إ��s��'�E�}�f���l�A\�E޹�oa��ݴ\�x��{
!*v�̷�p�,��2�׽l��t1���+p�/n��p����\�0��K(��l;n���ד�R�h�z��sv�FDwI]�:v���M,���k1��Vs�[�ƈ��i��.�Ev�-�����U�m*E7�H&�e�o6��h��;ٔ�0ZKw�-�%�������[�F;t�h�t���lUt��R���t�.FK�t�=/J"��yVj>���W	[��͔	DC�:����M�1�6�f	B��%��s(K��y������vTx��V��)LHt��J��Mٳ#;A�2��4*�2����w2�.�n�3�	ng���ɭ虣kW�cю��k.�cۗ�	B=�ky�?����bf���"����v(��S(PY��Ʋ!�	�lv�-�Ւ9zTLX��aM����ˬ4��Cx@əuR�ō�ge�zLAe�^�%R2凊�D%�B��6P͖���7Bٴ����H6id�w�b���9�0N�2�)D���7L��Qٻy���PJ�c�R��8�w(�6FZ�&
�5�v#M��X%�m�q��J���<��7t��a���KX�=����
bl�%��KfC���K�KdYj�8�֌�'�*�7z�0��Æ���[V�hOc���E�ĸ4�6	0���C3��^����Q��jw,嚴XŘ5H�7�ԲGF凙G��L�e�W��]����˭����f���r�E�ya�
��޼��F��(Wu	�����9B~��D?�c��w6:�!f�ܩC8����Z�(�oe�2�0��xu+B�y�-��+
���EԦv���x.U�i�4�X��
n���ҙ#M�P�.7����Fsix�b�RH���'PaYt�dXk2�c��\cM�4�y���X\h�Si�A�gS�a��;��!���W3כjv=�AQ���e]H��� M܆�^C�Փ�a?��c��\TF�@�Kou�^:�!�uwe�݃r��i٠EU�:��r�X�8��9K��8�9�59��mG]At�\x.,�\V�oE�s��ѹy��o�[�;%�p�wѡ��g[�C�>7P��̸�/26r��Φ?��������}�����i���@�* �AU]T@6E@�2%�7.UV�(���UU_���ϊ�����������<x𪪪������������������������������������������������|����U]���;)��U\��UU�Uv�eUU`;Z�����UP�����������ٺ�-@Uv�ŀ
�*������r��U6vŪ�����U]����eUUU P@Uj�� ������a���UUUUUU@bڀ* � ll���\�PM�U3�U]��������UUUPv]����Ü-� AUL�Wlڪ��UPVm����/X-)uj��ٕض�V]5����.�3u��Z	�m"�u9lL.[��n���,
ͮ��(]Ժ�q�nNh��j�	���8$�Ȑ��-�#GM��%5�.l�R=��b+���$!]a��.p�%4�l��fdU�M+��%ٷcf[tЭ�72ZgPp���Y�6!��f���(�R��[�tz��jF��Dw+�S^.P���A�Q1�h�ԥ͢9��&ɀta�e&ۀ�H�s������]h�:��R��1�ah��۳��6�g(2���L�,�9�f�̮�kY��cI�b�宛0�s�{�K�n�p`�Li+5,��]�)��2/J�%u����`���­��E�Q:�Ep`�j1����Itmf�0�`E�\fV9�Hv��ֹ;F��h��m��UR�U%I�ImnD���n�R*m �!���X�ش`�4i"�bF���{;M.��U�L��Zڦ�`���THj״�P�[-!�8���BV�Z1��3EՃ�r\JlU�]����"�HV���I]�$��HK-X܆����6�	�F�*�Q�6���v�L��j9��4M]tA���J�����r3����i(K��n�qbŖe�:��	t���]��S,C;X�j��Ք��&b��(��C��ka)M-+��\�� Z�(۴m�2�j���M�cW��ghjJ�(�b:�����#�.n/ST�35E�6�6��Vdi6�L3[,��c���Cd���V���[4�J&���뢣�b���J����4R�j����+�\�P-�=���6��Ymf�R�rmi�1qYu�끥)r�^Yn���H��0\KM����v��jT�M��k.�e�J�Q�ٓ:��e�Ի�
�F.�X'g.�W\��v֤���J�6<�x��
2�qJ�3M��ani�x�F�#]��B�Ԁmu"뗶b�69�pY3FQ�Cj���kj�SPlG��Q���[	��\���^���vu5	b�ش"��R�P�B �m6�Ĳ�/U���;��%��6. @�.�$Dq����֕J�e(j�3��fS:�\)�*mfm:��,n�]���ZQ��і��Z�	N.�$	MJ�V�c\�572�)�5���h& ���s���ci��J���-��CT����-8�e��ݵ��i��B
�XVTΕt-�7:k(:����&�4֙hRm{ b��a�L�.��2�t*3C8���ns�s�9�AHG�j��F�K3�Amcr�+���R`�
k����+e��:�D�<�e
Lg3A�4i[c���`50�)7d��TH�LmJ��!)uH�ŤE�5�,�h�[K֗T�Rc$j�3����n�Rڡ))�,@pU6�&�W��:5U���D�V]mn.�[�0ӫ`F�uR�CAeXk�����5`��]l�gB�C���:�QX�1ÙM���� v�ƚ�vM��Q�nxʰ���l�RY+1/�/^�%�h�Kir��W���[�����#r�n,�GM��G%�M�т֒�����1c.q��i���J�ь&8�W k�K�܊�Hu $)*]j�`^�+��w/Xi���P��8avhF�5�2:6�d� J��WEX��ԣf�i�\M.��e��.���\�7WX+�-mCe:�uEkl�(#C��t3\�޺��4{��[��F�jr%�a������b�m�]�d#�Z�H[�˳*\��)kƻl$L�6�5����r���-uV��a,�l���K�!#�ı�t&�VٳV�!r�%��lUB������p��n�Y�� �Ԉ1���%�`ږ�ʽ`i�fRM��
Yd��%֙-�P����D-ѳXSJ��4�%i���B4�ŎrK������.�u�J��	x�(P-ۜ�l��+u���\[ y#����j��j7���1�*�gH;j�°�tfY5�4��bl(���8j�]3F�,&"0�]��%5�5���1P���n
�dۅbV�bF3!ysH]�k[1kH�a@�B3[v�Df�fG��ڏb��]�
MhL'mسRK1f�fa�y��`�gZD��^Π̬�TΗ,�,�ʵl1J0
J�,�c���Thi��ƙ�d�t�4�`8��ԱI�E�1�3%��46[�\R<��TFXKqæS=F:`-6�k5´��5��lfU��-���g���bclࢧ�ˀM���)�Y�@�F6l�3
JB�RY�R��M1
�¥I� 	f�b�RL۸�WEf0�6ն��k��@��2��@��Yu��L��d�u�d#��ƄsvB	����ٮ��(s�Mf�z�D��B�B�  @&L�+���`)/f��fmA�B�.&P�:��k�\B]d��k(萊���ڔ��el�u#��kH���
%5]5�<$5%�fb�t-�+��\��Yl�B�B�m��Ra�j��t�NmݫY��G��cYf�C�kq�A:�V���@���TiR�l�%&iRX[a��8�B[����pFֶ9e�D��5�&Ku�,�2ؤ�(�����V�T�͉����e����hQML��-�!���ZF��R�t5�lk�u��mf*�u8P]�2��
��"��a؈��4���&e��.(���]-qJ��:�7C2�DM\��*hZ�ey�0��v�t�ݣ�WPv�BmEк4F,�v�q�e��hv��\J�\�f��K�RUK`��T��P�K�����.�WSK.����E�v����u�Ye�ѕ��3U����(�b�������pJ:¤ k����[�uږюX���n�n\(�z��j-K0��������qt��c)2p�R-׳�(�w!�ű&Iq[sZ�JX-�bF fiv���ز��9�\�.�A$%�Yr�k��f��[�\(&�`�uf��P��
�u!u�MR[]aN	Yk��a�K,f�9��l�J�+����+&�@�����a�v���fU��U�&�6�Bj��Ɲt0�J���v1k��JM\�iE���d�)��\6�m�](��
i�c��f�����]��k�%�hl�1B�(i�5f.!� &���#��	�k(43a��\7Mr�vt��6-�l�#{T�c"h�ۆ��5�{\B����X����v7;�::p3v%S���6�M�W&͸�t5����a���4�:���k�G����\�FL�.+�K�k�XqF�]�$��R	u9й�P�Z�+X���iq��[vk�t ��ʹ����nk�,��T�2�3sZ��SmM,�m\�D�x���h�Ҭְn�^���7;e�X�	������yqp<0w]-��)�K��=�a�Ⱥ��K��鈶�A�Ya��I��M���B���J����v����ҥ�K8�V��$#l\ɒs�@Zf�Z��j���uj#35�b��T2�5GC0.�q�6��fU��,4�K��J�[��G����ʣ`�hK)��B�A��H�6y�.�kXT�he���qV�X%�љ/lB3I��Ґ.�P�JƛA�"��3S[6����1���Q�/\�#dQKԆ5XҤnZ�l�Y���n�̲����ᘅ�Դ,�i�+VeW9a.�.��V�V�lĹ@�n�:�^�gP�żQ�j����X��Xٝ�Mu.*7
����0��l��0r���l��4�f�R�cRc�bn��H6�W���)4\��Bʻl����5��V�2�V]��#k�5����Ą(�v-�eZ�j2䫚�����	�M��#��*��1Q��s���X-���R�4z7Y)f�c+��h[�jf�m��r4n�r�RWX��&t ��j��˶��.�f��v�B�us,�ZE-,�eك۴euʱH��Q)�֜bd�hRi���2��3� j�%�S�a��L+�-tu���`7J����V�^�ژ��T�]��,��f��B�k]�R���H���..�.`l�Zj<��n�&F`�LGE��{fb�l�r\K�i���f2�yb�����$l���8L�p�������Q�e��WT�Ё�6���LM2���`2�4 �giv��`�254l����(WYB����f�B�hb��sq�,�[��F7��,%�R�61��M�L-�n5"ƣL�+����]\�IM����)�����Y��6!c���4R�1-0����ƪ�d�jS\C@��&��Z�� �My��;,�f�l��6�j�B2�+��]��wRաs���6�XEװԧkB0#�����e�@]����e�kv*B�FS+R+.���[ڎ���b�چn�b^���a.��v&�h�Ke۰�h�R�D\mf����*e��nRm+4i��հ��D� ����qմT���n���˕�c�Y�c�+�U��feK�(i���ԫ,�r��=\[3`YbR7F4�]���X�5���9Ě4ZV���A��͘�ٴt�U�BR:��`x����e��4�[��I��hW��n�P�,]Sl1n����q33H;c����te�S�Cv�-%�$s�ʺ@��	��Ł%��88K4@z.HK4��,�4Թ�������M�8�-�a
&K5�,1��%6��n1�� �9x�L�1�7$�*EΣ��MuD����Y��Y��QY�0�����t����N�;�N��_O����w�{��N�������������ߟ����I�$�'����Ϲ�QUUUUUUUUUUU��N���?2I;��ӧt� t�Ӡt�t�;�N�t�$���I;���������U4�o�W��1�����m��o��t=���!���@�.�x.�I�i����m�I.�!N�nH$)>����sK�E��X����܅�lɘ����	�~ꙭJ܃Ʃ�T�r�}���j�ۍ�M�{�AуDrFR�8���XAfĭ�}�}��1�t�����C{}�^{�c�OON'�6�z]ߝG��[�͖���$M
�����#� �4�mNÑV־�bwQ��Mx�Q߮��I��z�mm˩m`�Ұ,�.卫��=��FLj��i@���-�&b���1��s�vboz����V�?7O���I��OյycSA�oGy-�a��o	@�b"�ܳs-��ދ}�Al+�� W���o){�+�>�gI��L�e��iLkq�\������V�0!�Ew)�ڰ�x�ѵ��+7฻Um��u3��vc�r�J+im{
�ĺ�s{�{X�ӟG���>����PE*�8�Y�%6�/[�����;�Z˸k�Xឧt),��m���� ]���1�T�N0e�u��shn`|*�4KڛnT,-1Q�F�ޘ���=�����k��eV*�Z�.Bg6tʓk[��¥��,&K�6�mLX���.�(a�����hJJ�]2\��J�1�M��\u�K&�H�kph�r���l��|!J��vF���4Ĥ�
�6	ɦ�X7K�
Xb���T�ff�h�*�^�ҖʳLia5��K�\l� <�6��1�⃁�G�.eT�Ms)b�-9򑦩�'��y���q�jŲ�_6Q�=����ޭ�XMH�-��o���'�>}��,�s���!�$��������w��\z��aa3;:�NMlgr�����&�P�tL�n��_vt�m78(��<H/~�]��FyY����ޫ���
����18��m����h467�%dR�/�
��7f�9��]�v������>�9�z�'�/��З�nwHw��B!Id�����u�kx,�G�.ן�n�5���mz�g��N��f�޷�����\����Ig[]囐{��o��EM��J�kpf�y���ɒ꘠^P<�`��k�Wd�Ç��]��������z�8m���T�<�V�+@*T�w��+�N3�S~��O�nb`<��z�+�R�J��2nD�r�6�Gw8oHgA�{s��2;�wFL"�@��E�5��Q���9>��?�G�����������0wR��	;��z�k^5����/���O�v�]a��wo�Ev�Z���b�l�v�U���������d��:�	91[�=]d��ǆ�E��86�=�u�٘�.K���\EN4E�q�F��[�e:�vYHމ�d�
Y�e���6�[���ӛ����-u#�]N@ڈ�!��"���*m��bܩ�W�OJt�a��9����Q���B�q�%��s49W�t�)�
�B�=�N�ug��Ay���'�<�;�^^L�s{m<"����?�}ޜ�?&��.B�x;��ܳ� h�ۂ4�:��!�W�����ڐ��ݕ~̊m��s�̈W�z^gm���ږ�	Ɠ�	��j�}��y�w�S��_%f��q��.%�a�D{���Z�����_+3ץ߼���\�!X�s�X���%kT9�]����'[x��6	n"�)Ĕ�l����w�Y�j#	��b�	��=:'�D�i�+��hm�n�V%��s��Y��ݛ��K|;��IVAHP��z{��qd'���ݓ�\���-^V�2�G2�ei.+n&��U5���ԅH���ö��,� 
^N��^Q�e:�<^�*gDņD�VS�S@��=�׶��x������p��z9c:�y��.������T�9K����<e��-��	ۮF���kYÉ�7��0�w�|׺G��g���D�t�X�������)Ty˥Y�������p��ܝ{,^ �*Q��߼d>^jb�N�W�h{�	% AO�;J�΋vn��bK�wMT�T7��?�Ն�h����W_>��i�A�v�oR8*t4z��l�C� ��	~J��a�M�!k��J�s���X��u/޾���~��o���a4�������n��g�D�p�Uj�E�[	t�:Nz*��j��+i�"�jx&�L����hX!�����SsӔ����O}Ͽo&V��o��2#F5D�B��D�[۳���&;�Y���尥h���bM�3 ]f6��၆bTFJ�f�-��C0V�?G=�G�g����sKa���}/7tڳ�^�t���ފV�:�l_ì*F�mX����M��'�� �;׹n�1s&�|t��s���S�_�`�i����������
V��_���9����l��w%�Ϯ�Z��#x��8���e������sn����-]Wy�;�c�b�]1����(Ԓ�n4eϠR�n��_�i͓]��ܱh�BS�Y��u�^�M��0e��^��P��[��p��.�}cjnʳ����=WGرy�=�YOW[>g�:�w�����o���';�iY��{UV�D��-@a�9#�$f�{� �1δN���q+��$�v2�p]u+��v>���r�����Qd�m_��������QgG�5���zػA]��w��gb����{~�uϽ����˻��{tq>�"SHG"�6�������6�eÖ�\]��;L�	�?=�7�݌=���2�V��]�3hg�z{1��Ki�����r֩�,B�qi�����f�ߐy�5�؉ҽ�Z��zg��i����Y5o�yH�no�mg�݇uWHG9���q�q��	�u�mĨ�yd�gz�Sc6�;{6�_o��f�O/k]w=���
��$S�j�d�"��nR���ֻ���k
c.�~��D��5��������g�J�Y�[*�����X{yI�f�����6�^���z$2�kF�����j��̴UM-����rer�'
��|�ǿ^����>j�ECZ�������h�M{w�6U��y,"(ղ ��J�F���]��2ː�2�0�V�k7f�@u�f�h�ؑ]�9���n.��Mh���Z�ؖ��XEcc�.5����"��1f�^��雠u��f�J�\�X�5Y���6�nxjcm�1b���-�*��h�ٹ�قf��Qض�̼f	ap.�.�/)��I��:�r�7�R��0p_s����n�}�#,�۹���Sq�Z."G�zPy�d�P�m��~O���|��d��H+�kx��K.�����F�f��>�ف�xw蒽_�1��$��(2�o�fв��'}:���|2Z�}�>xކ�-���F!��v!s��J4����l<�*�(c�D�p�JI�B$������fkM%���ߠW.wu.��3��qN��]+��ڳy�wa�8F��HZ9�����;����B����l��,y�~�>����5޻dX"�옻=��Q�b:�9pKwǘyav�TlT�reBE�u�=���;D5{^rp�t2�{7���\��U�:����Bu�1���J���5��L4�9gZ'!�*{���yU��Ӿ�	���j�GO_#�:���{q�3~�����n`/I���Gs��32�p,E]uf
�s��s:�)ԛn���J�Ke�p���nl�9�i�
�Y/*�x���P�A����uʡ��Yڀ��=7����jv�m���ʼ����S��rմx��F��ͦݲ�.��gdҙYo$	�m�#��Թ6c�}~9Z4)�k1rN�&��0Y �2��4p�fڎ�Ի4�6j-]H3%�D�e��X�3=���a|��ԡ��rlh�o͋�<+�9�s�EP ]�a^-��L̒jW�l�4�;�C��5]nE~� 8�u_a�#}�w���n�1�o)�om}���%�/:e����e����E��|�.�K+m�G���Ny3���f�_��m&l�݉b�Mx:��+A?�	�T����[iȪ��ݓ'zR��#Z���|<*�C�Z�u��y�sxM�5��t�R_p�.��'J-ء�%�U�=�L�'a3�F��W�ظ��vrϦ��U~-#�Bb�*}Sx�)���k}���bb6���-�����G�,>��J\�����
_!��s3n斺�dP�	�nc��Ĳ�v^Pp�hJ�BHAc�>����w����UK����Y���s�l�"������n~�:M�;`��fh.��D��T���.ƴ�x,R��r�3����{R���+!�#Bms�*��AY�
l�*���1�9R�9�����[�6�+�P�g��r��8���K5wG{X�Q{�j��A��V�(�Z�R����d��ҊQ��s��P%*Ww@���ܫ;�U���e���_Mf�*j<�$���ӻ��m>���;�?FN�i������.�a�yi����4�I�Ӎ�I��׼��������zx������ᢤ=�<�ܝ����ȭ�3��X���]�Ӊ�J�-t�sZ��;�{u��~��~��9fJR�pVa��-�Y4�x>u+�,�$lz������f��K������<�S�K�g�SyZ�̭�F� U�)"�inv���Z*��]�%u�[m�W)Nu&Ql.'�?>|*��x"Iw��n^׸ّW�/�F�<�[`���8��*�R(u�9Co�����X/��~��1�#��en!�^｜�Ry�R�KW�W�Wnu��N"˻+�$+�j5�L5皦���;y/o�t���Mnx�2ۭ�2���@��XM�*�kxjr�s�� *�=uJ�i�66�)��q��J�u����NKڔ�#���4޷={���d�bAR���~+P��M��._B� P,&�r�`|�w��
��<}���$�2�U�d�\�OV� b��(���Q��:�ڻ7e���"�ݮq:�.`v/OBt�)��>�)��=�����[�f�ڇ�fz����w'[]�WS�i2S"n����A���QIcS��~s#�B���%�,"�����Xj2���2���A�y ډ��	��L"���n+$=��*C�w�"�fu����ݞ��tq�.w=�T���r*&HI��V�R�!X����������x���[�ކr
��^���^���L�ٖ�����.���o���*��n�IQ7C�,�:����&|Ew��wܬ{/_��#j��7�{;��1�g��qNV������6r�I�@��S������	'V?NPS~�[�ڛ�~��������05���]�f!y't�i풭۾OT}ySI�QN������o�LU�{a]��JSj�������������b/�K�wb��6E�H/׋m���a����Wl�BlF��%3[����t0uŢR3v�\yB'��-ܱ�3&����qa��1&�sjh`b�[omw]`&q��G.m�.nf�M&���,F�S1.�+�#]R&�ah��4�2��7,��kf���h��F��hR�4ee�0�v.Ak�c����FC+F����,��Զ#�B0Ɇa�d��}��Z����$˹�<�^m�.���o�n�Z�׺�4�Uvn�<�*�'VOMdynEoe����A��A�A��5����R��n��s*�ԛ�- �����&ݜ^k V�'�T.��]
V8����ޙ��<�:��r�E ��k�9�)��nV���bk`���jc���B3�j˘]������nnsf��|�E#�J�$��p�ۏ^8��f��2���TٺEQvn���Jjv����߲�����Zѫ�y"���j�]�*^��c?-�ag�l+!��2�r�{��5*f�I����Vɷ��x�Uʊ��?7�fg�������3pJ��ҭ�6[�odK��P[�IHE
)zM�sS��@������q�㻃Erq��ΏȆ<�fѤ)ߚ��X>�)��gd+�� (>p�i((�.B��;�=�����y�'���"�0���r�}=�|��!		: 'z�l&��{\H-6����ǋN2\�ŹP���8mr�G���ƌy2�v:���a�U'щ�u�8���O��f�ؤso��l�����m0��:����vl�w�j�,|9�<�<٪� C ����L��2X)�dK9��s ��y��m5�n���o�_��]��Wof���h��G*w=��s��w�Ե�M�4e�Ѻ�ɉݬhq��\�·{��G;LH�-��l;�]�����[m�}{�ј���u}x	Y���)3��1K|a3�;�4~��vK�fέ�$8Q����Ƥ����+�)"��]fr|{�\W��k\�
�,�tҗ�l+�j��|$y5-�f��Ų�w?�+���X|��}Ma����,�:�٤�o"z;��6+s�G��F�������t���J�7s�,�����Hr�_C5sTDlU�����ٔ��U��խ�m��j�Y�Z��H6�r!�V>�\$�'=�?T�9��6U�~���K���7O�oecǎ"3�u�g����L��;����;��gD!��1.�/	���R
�gSA��L�DѺ�u�^�02��(�+�Yő�fӋv�+��W�+�CF����6�f:݅Yڨֹ|�ge�Y�X=�mɢ���0��C�];��;�mX]8>4���,��-fU�Qe^�^q��"em;�8�m��sG�{ظw&�í��w�9>ڐB_A[؉��70�άJ���v����ݧp���eUuR�`V�mUP UvʻeTU6ڂ�쥠�Ur�S.��+���m5���L���e�ðAZ0�f2����R])V6��E6BQ!ns+�E��\�u�j�R����ڦ���$-aC#��\��b:/]�R��%�k��6 5%������A�f�P�� ��+�:jl�iM�Z��e�ȕP�LE�3C�mv���U�Npb�6ѫ��%�L����2�`��i0,�37K����kN5������B�
��cM�pP7::�5q��A��&�8mmd���+&e9 �7\^�V��C+E�ݥKs��m�%Z���D�J����M�����&de�A��X���Yf���;`,�7i���l䔶��1wCU����a-��.�b;`��ns��H5V�my��(��C]Ve��e0-K
爖k�J=mu�p6��z�H$��v�3U �+Rjؙƕ�m(*nU�̈́6tB^ZKń�H��
�f���G1�3$p�v�J�5�$r�l�u���)�&x�m�YPԷ0�\��@&���5�
C��]�dRҍ��bY�n��ѽ���L��B���έ�0�#إ�K�d5&B���5X�l�p4��;�x��,څs�ےV�����LaR��W)����+
�2��@�&�GE��%�u��2Tq��mՂ��`۫,c��WP�V��i�;4��lsm��kk�sP��B1�Ҕ@�2��[�Rm��:�,f����ڴА%�p��k���R�x��9�X��W�Xk^��E%��[X�q4f��L�Ga��s���*GL��T�I�7��Qn��{b�=I��ִtM ��my�Ai�ŊTfY+�3��u5�Xl�L�0��ccD�ilЍ���SlݍQ#�h�c�'g��G�[u,�,`�P�6��l����h�2آ���3c��ݭqM���&�	p�������A�V��*c���*�Od����W��i�X)CD�b��.��Q�R6�;
�5�������d`�rҲ�ҍ[4�ו���.�cT֔k���ƴ��eF��Р�l�d���V����{1)I�k�u��X����{=���`��N\��/���/I�ÎA"�@6!�3�r������~0��C���CE�B�x�=�;Ck+��ߜ�'�w3�H{ӽ�i�Ty�M�8���w�d�2wЛl8m�H�񡀏	W�&���P�9�{]�<��˅^�{Z.����'��O���T�h�S�y'G�=�ul�τ\�F�?r��ۜ-6�Լ�a�נ�Hш�o����ە3+���N���1�enS���PF��8��ڇ�j���5�U�bo�rCD���O4f�[���X��h�]�_p�K�8k��߫p��ȼ����]y	�S��5�N����X9>� i|P=������'��̸�V��9�6�~ɮ���}#�RI� (j��t�Ei�<��t/-c�/8�O1tx=�E������,Za0h�&F�lma^[-1uM��e��-A�%'�E"�A9��S|�*�>�F8�M�]6��b�IV�w͓[�xg�L_�x���=:�(.�4�xe�(�L];��~�Xz46��dyn*��/�Cy�s��3rIû��6���6'�Ӧm�`���HH�����Y_+S[�}Sz?�}��kMt��}�2�X+7�,^	��W�{J�~_���%���A�ļg~7�YM6,��I$UX�\�	�6p�9��@w���^^���)f��+}:�s;6�����ډ�P��PQǈs��wTA�V̚e��-�6cs���`��(&�@���[Y6�띲+�m����F�M�}�"w��]A��R
�']�k�Ë����i���*�����e��R����v���;�:��/s�s�Cr�R���,k(.�X=8�8vխ�������x�C�X(^
�t*��F#��{�v뒃�O�� #4h��F�ll����qpܬ��Z���ޞ�w�0���U4�1aJ�Q�s��Z�V��X9D�`Mِ�E�^f�U�
�7bB�2k�u�ɏ���f�N�����Ld���_kߧe����f�$W�� ��6s&:�z<���r&��ں�:;(���ewS����h��]>�%�=:��v/����ɩ��Z�g�P� ���i�<0��E�u�k�H�~w׋�P��C$��o�02]�8�5˶@�m�Yݺzw �Z�0�5�-��K;[�Fl�L����B�ͻ�z�1$�[m��^��8�4{g��Mʥ:~���sǭj�8H�B~�M�B�V���4�"Խ�����.�3omn��=� $BH�*���~/P�N��rַ���}u�b�o�]�3Dfޜ�g
��d�ǣ���h�h~�����{9��{�$�yd�:w��؝�pw����:WK�a ����G�*�ޤ���l;��}�P�����R�&����k���*LA����Ѭ"��*$wy`<z��.+���c�͹]3�#Y���Q7���p��&�}bUō�h��G�,�IHت�ջWIn�����/�����9t�f�p&�P�!�@���&/:�ŭ���IpU��{XJhD��'	`e�g0���h�͵��֬���ҧ!�s'�0v��\�ς��\e1�z�Ձ3�=3K�U���{�x$Kh���uS&ƻ֨�[[N�X�~��K��I����K(�M�U
k:ӿ����+�g�K�u���t�2�|�f�8��9��0�C��~�����Ӥ�W����م�aY�!�l��:���yM����f��v�ƍ��0ٟM��dQ��|�e����g�z������>+�SA��Hd��K�-웍�����E���S�ٙA����|�z�܆+�|@����4	0�9t�,t�
�7:�_^���($��S�9�蛴����V��MXv��
v:�[����v��z�ʾ���[Wi
�UB	h8�+�m�L7ST^`Ko3d؍�ֶ�1l�5m��0qe�`�C;1�+�QZ�2륔�R&�S6�I������0WU�����Ա��*iM@%���uU�� ��7Q���,bW���@b�f��`L���h�цɵt���Z�&�.c�9������.t������p�����1\��JnюWT�f&�h����X�x���D{-1�?Z's�Vt�h�����>S��ҵ��4K��������ݐ�o�`z��������9�����3Ms>ϻ|;K�>��Be|,b�>(�'��ۛ��Լ��ّ��$1p�J�צU:�m�fe14��Hz� ���l�p��3�\��i6B���t)cf��^�gL#��,��[��^��_�W���+�sܯ�^����0>4;ǧ$+Uz��nrJڗ�Xv1�9-��Nv�?f���6:�����~C�'��JL�3o��N��ξ�B�H���>|�wyޅ�D�>�"wْ��k����n*� Gp�i�	��<LV��>�L֪�h�"�y�>�%#8�4�k����YZ�p�~�.8Б����z�oF�����u9���=�õ�=�W�����a��e�?N�P���o�d}���o���M�v���<�����C<jf�����Gd�nX��SC8V���3c�l�`��p��x�m_���{,l�_;���t�WK��PK<|O`�+%7ctF��]��9\�C��X!�ŗ�La�N�����o*��:�n�vJ��t���bͧ��\�Ke�`�c��1�}6Ϸ�o���R�e�Ée����M�"�H����������p^��UQ�EA>F��U���h�["��(��b���N�ki-����q�7T*x%��;��_8����p{`�[���v,T�+X��>�.�<�f�߽����IA騮�y<I׬J����Q4
G�^.�خG�ںՐ��}�d��vE��R�%#�r�$D�q�2�����u�ڏ(Ma����w!d���^����d�Y;�vr�f��r�T��T� ���hP�����;<��VO7+��k������>��w���x��H��N
�@�2�Wwrc7�q��H�:s'�1�
;S��y9�LI�_��[# �qn�GV�H�z�V�e˷�����}H�-i&B��)V�_�%!o��f�Xh���1��W���FE��m}]S��ª:���R9�<���](�s��I�'2^��2��#y�B$&ȀZ�"A�h;Ŝ�]��vp��9bt�؆�"�o�ǭͨ\�ĶK	t��hʎm�$8�-tM�2�m���G��g��ghM1�wln�]g	Bb��v*�w!�UD���J�4�簲\a<b��;�z*�w+��,=��N��2G&&(Ѧ����g�F�-ʍ�uaU��W~Opr�2�p���q�%���i�W�H���pPU�nJä́v��5�����������^�*�D���`^�:�\��:��唤v�8w֝����d�;����z=��I�ګI�~=�V���rK�2u�R�x���r��A��.�3��*-W��MO���ۗQ��gd�'��5$��W��/ϵp�1/*�������E�	Am�vf����R�t�.����L������E����]V���5����n�.���6=8Tc�S�/����ۡ��9���R�m��!�S�Cb�0��
?Z�g|w�*vw%�0ɨ�k��gLlbc|����3�]�o��^�#%�w������(�i�Y�K��o�!WzסQ�8�4qi�$��;�v\�wǩ15���ǟ�0�t\ݫAu��T�J�]����2p��Т#
@PNO���o�8�����L�|v��31�t�h���;�N4E�G�gգ�%&2u6�Ψ^̿d���ߑЛ�fѹ!�^�fJA������c�H/u�}�N�>=��2@���a�񮾜�ҩ�.+P���Y���V�P�E`Y/T�۫�wb�kC�b:�:���ڜ��̵��<�6�w~鿄pJT�`����ׂP����!g��맲u�;7v���`T��ݱ�z�����Z���*A�Ƴ��}"I8't]b�*�Z�fb���� �llwR�+q ���Q(o[��S��P��삽����޾�wkH�Z`����,�@(kU�B�(`�Ļ��5_ڧ>o���K<2`Z���]'��%Ϳ�b��q�����t8�Zs��7�r�h4�-�
m��;����ύ�J�7L�{�[�/�n�q8�����-��O\��%m��qU�kc�⌂�-���U:��^o�7]U�q[��d��6��x�5͍��hw�{��������<O	�Kv�kba��4�b���Λu5�A��b�"�����g�o���v7�_��a����W�VA�d�ia>}���͋�k���JP4k/��3t�Ak��AA���<=��m)�X�����Ա��9#� y:z\@o�}�\��OL��O��gB���J�
7צs�A?id�i	�M�B��<�n[�O��$�bq��u���Sq`/�b��Y:S�"8O���8x4��17��}��_{Ƨ7�݀C)���`����L��]�3�Ȯo�����I�-�ӿ��J^�ku������j��6�}��LE�*�%��z�����s��IV��ݻX����*�����$X��Im$��D�*i�Rћqf�B�n�>"�xƥ�A�ppb�1�,;�5�`�/dJX����XGh9� wm,�������)�5�h��!Ā�%�62�Jsm�1�i\n�G[eu�*���i�V.c�v˘�n�γF5F����̹��T���]��\����Nx��Q�q��f�&ƹ�X3�5�vN!�_�%�;����W|\�G?�"�v�@�2�&��]�SUӞ@ 4A����LI�uy]� �f���n�墅�JO������'?��zL�_��i�4\�}���/�w}px�$i���O�y܈i�i��� ��x4x]�n��\"l�y��[�/|0�L���cQ��M�q4nvl0�kX!�lN
�a�U�d�ފ�N�d��aS��/f��{��Y�x�r�C���Ԗ�t��z�z�M�Gd�x)��#��!�`�'�f���pR���>G-{�Xނ}�s7.�l�^���Xl�J��<.���	�L�I�7���׀�'��
��J�+4;��骺,{J�h� �C�b��K���VD��L<�c>��B�]����j{�V�Oz�λ	���!�O�)������ʹ�^�`v���p�Nl7S�7���Vqn.�ט�4�)J��:.ǽ}�^����oWw���jh�Յ�mր�$0��Rg@��޹�s��\_U9x������m���x����%lzr��y�]]�ƺ��$�@	�}��G�v4>ΰ�+�K�σ�&�e��Z���A��� I9�3"��U����f\i<�Ď��j{8\��Z��cek�"늇^<x��Dڈ���g�{��_[\Ѻ���J���[�����ЂJm���\ކ�y��^E�㒱Agf����>z�{Lv, 띶ك�YS,��h�q]+���4�a$�J �W����ɥ���ۭ���缦T��w�rsuoc��Z!ł'̿7��Bd�yx���^��seQM�ԏ
�y�m��#�z���A�s�����f��@X�����Kq]�k3�Fa�Yk�r\��MrsƦ�J����j6Q`"���:�d�$v�g�H��ݤ�p�=2:$>y���X��7���S"����i�>ɩ$�.;���G���wc�Ax���r���\B� ����k�ʲ)��o�d\0}{���l9�O�y��oM0�߉4tj5���b`͙s̈;��J��M���3��9�S��#�@�A� qԡ�����<�c��놣�n	�^�������՗�Q��iqG����k�Q�C���:�臗1\�d����={�3��t{1t�qs7�yr-�����H�ڻ���ʚz�/C�8���>'�i��.M�Rd�����J�v"�`\�6*[6�-
�	BY)� N�Ӟ�*�=�Q�=o�tk�%0��o�_��g�=�n0�Ǥo�{-%>{x�\/e%9o��v�r�t��Zvf�G��7k�e�S�

���9r���sT��n�t��.�u�2D&Y���KV�d����{q;�\�d8�P4�ds:����O��2�}~>^�(�:;%`݃��.%���}o�pA|�<���ظ�a�l�'�K*U���d��m%	�i���|�<��fT��IG���Sƥ_\����l����7�d�X��p��|y�RV�}\W��=I��������L�J0�� �Iޟ���Y>�S���_��z^�O�}R�{E�����L�.�P*x�Vk֥%���k?��E�ݪjO{{w�.d�,��Y��}J��wi9Ֆ{d&=����=ư�I�;3�kCm����s��>����9}����ڏ#��U�q����e�yُn�^�Qc<40bEF"-���̝�*��LI���'sJǮF��8-�Y��~]�d��T;SV�ƶ�땹�n�R�A��m�[ ���+ٙOwuOO��9F<�C�2{�1a������uWm��\��=y�>���uQ������C��yb��de��{��V��Y�1���ϗs�:/N��꾁�m��<���Um��g��eg�8���#�����ݳ�]憼�P`f	o��/���` ~�T�SA�c��ފb�'*g8�Ԏne'R�9z*΃�r����ۅ���yx�X�V�vօP?��;��F��+z��zfi��u���ƍ�.sT��ٺݣr9��Kv�ձ�ϲ���u�rj
6Toz�>�۸%B��.��޲/ΰ�%L�'Q��-�����2�0+z�TTh�k��ŝxw3`�ɗ�2H��Qy�Q�?)�SvA{�b�p�ƛ����%����;�*�
��P��=�u�Ⴕ� �R����4������G3��
���߹���Y�z�e�i�e�|@fL�窢�h5F��Ԛ�n=F��bMӓ�;DUN��)K��b�\�S3���-~�{u���e��:���[F)7M�d�/u^�@�d�^��͔d	�x�eX�c����u���zRZ��(>�R;N�%�_y+V�or_-/���4A-�	K�XC:�7�$��g)`�G9��X��[�;���霳���b`��5/�������0�ރ�]x(��`ď:��F�eu;��'=Z�������e�N�uۮzr���M�}%6`a�E,�-��nZ*ț?T֖�	�ٶwd��Q��.(��P��S3T|k�LZ������������x��@�����9�:8��η���<�����^�y.x	� ����(�S-R\��0J��1��.�h���fmqvr��^܈�ue���_U׌�9ҹ�@���M����ccvoe�̩?eh< ��j��î��ح��W��z��_�z��⪪�������m��r�̶ۄ'�L�s�;>��o���=�3������ F,U�u�v��SGZZ�zף�p��jD���M��q"��s5�ֲ���q��t��t�:�zo�X����ix4z���yD���]�rs��2F�<Q����O�&����Æ��]qOI����ҕ�t��Y/]�˦D8Ԯ��gyF�.��Aomߦ]���Tv���7W�ʛ;9���h�(f]ˮ��]�$-�Bp��/O���w��T���n�ޭ*4�1ڋ��j�7�!��q,j��3[v����Z�j�4�.�l���քm�Pzz�wo>��3��i~����ܸ"l��p��NU{�>�f8_uƗ�^���Ol����cW8E�PI�\���
ŨԞ{֪��&�\)�����f*].�bjk�~��u�	(���w�:�w.��Ү�N�\X�}��(�{ػY=�Zp�p\U�|T���=W��	v}š1���%c7�DY�������3S1�0=��f�̷�=,��z~��������vu|m���<�s����<K�B�ra�@�7usR�*\���g�Wu��֬�#-������Ak�3A���C����<=�d� �	�;A�hX2��\����g�������'7��Si���Y8��e�b�R1,6Kv���ִ筺����#N%ڮLi�-m��3��`ĥcA����u"`5��l��#li*��ѬPt��&�[��̑���+j[v�)p��"�٬a4rK3s����f#�2�66-6˥�W[��U�bGF݇J;���R�����*����Tl��iVhjk7�q0%�&�^�D3�Q)s����X�S]熏��?@��[T���6�LJ�sg��ӝPĭF��G'z���:��8K䛋C�.������3^��#ؠgx뛳��y����tdࠇDگ����n��������{��O� ovUՖo�U�I����H��*
��@�j|(HQ�k̬�.I����N�3�9"T/��"��$pI�PeF��	3�u�T2���V�M2���] p8u��~���<޸�b�-Rz�e`���Ԁ��d�=O�N�~���7z0FWlf=�٧�ˡAM�����\Zw(k�k=��ɕ|mE��T!�C��O�Att���1T��ţ���`����4�w���>��ݟq}s�a�meA��;���D6AA��Oz^[{Mm�v�&^�-���~�|���	���ՙY�{�"�SFne��$"��_�;f��q���6�2<�Tl��˳�$�Uls=���D"�g���d��Y�Ơ�g zG����wc�8���_�}�s�~��Q�A�5'��ƪ�[:�#��`2��7���3��\D �P��p������ۚ���[?&N�^��Z�e����n7
�d����MZ	(g���o<B=~�������k�ib�m�������vp�۷���R
��^g`{�h�uG�/.�7mvb���y��Ȑ�p������F��DV��dق9b��վ�*�twцӀl\�PT�r��t�{��70S:�ɟ y榊��{���m-�ff)b�"Ѱ�E��:��#�˳�,��Xe�A�L�~ݭ�xy:���Yn$�7�뇦�O��>^��J�����5aP�7�p��{���x����
��Zג��8a��s�ߋ�~�ʱ.�Û�iP�賁	�e�N6P3[�tn��'�]b�u�雱�~[���:9B%� -������@ '��Z�����hH\�(
�t�bA^��t���j��H�,���1dC۞ڪ9��Qf��A��ާ�w�e���]
����a�S�Q�i� �}w�,�&(b�q� ��������T��, )�p�[^��Y0����VI�Iqu�2_�R�dk��dƴ�����+�M�C iA�DO%��rI����O��AvːE���7�W|�"C���8�k�<�D��vr07��y��7�2Dr>�+�b���"|Po4�B���P)5��aK^��L:8B�@�1�Y+�O�P�z��/ �F�\=�$n�NGSRZb����R�j��$�H�s~���C������Gd�F�T1 yb�A#�xf��5�֍�� iv�M�lٵ�4R2��+��$�כݶ���I�g�B=��$D�Y$z��H 0GI�(IÃ��WT.��f�x4�����ێ���(V��pS�n�9�]�d�7�]u�:�R=����A��k&�py �����]�c��9�n*c�z���ZuS�:4=��f!q��z��A�BEfO�Q����Ӣ���5����^�D��6g@���o::���qr6��Tf�Tk=u'�G�J��?V(Q=�/۽�qFP�h'��bP�-����4�H�i��D��<������&\'B� �~��Lg��;��f������^�s�<���;�y7>߸)EP���R����i�N	��D�Us7 2{��	���u�Mu��e�L{�H#sˮk�v/��n������(?sc��EL�Nyl�&�3,ɞS!{^vUG�yCÂ�$.�y��dw�fW���*����������9�t�F�3�^�Ĺ�x��_h��	�
��2�c�c�:��c�O��~��]�O�9Y=� ���~	0U�"8�0��3�k�r�����+�k`R)H&HܖT��s]n�P���8�"�\AЕ��f*�bWh6���G��w	����/�ط(�P=r!g0 ˍ�H�y<��m��.'p�Y������\U���.��i��wa�}PP�j{�%�z'��;������p@��mg�����y1�x�M'7�?_��1��K�g��C�9�^ʙ�;���)�L����mH	��e�w�1�����ʒ�P�7���SB�������?���;��3�<�׹=C΋��s+__�$�K/z�b9X��΋ɉ��2m�f�Y���e�~����.om���9>t�:7Mj��I=�}U��F�uw��vm�y{�]�>�m-�����~�_w4�"A��)	������-=Gr�����:��޶����3^>~���&���g�DH�W����kh!��@��<{��b=���W�Tsx��pm��&��'����ɝW��;h&ھ�H�Ӓ~;VY����� ����D�&f{��I�jj������#g(-]b�0	���ŋr��阩�5���DsRmFE�i�ZlO���� S2�d\V�dy�2͇��l����\%����`ģ5l�lX��`�H�4�Q4��b����F�w�T<���~�d��鉻�Ӌ�)�탳��I�c!<��)�¸Υ��5��uw�=��� a&���N�q���_�v�q6B��n�\�y�m�q�@刢���шyz�O�����9�[D�k�y�n��=^^�f��'�;d�1VR����
7EU��E�:���j�:�c����ϕD�n�)G���w'��f_h1�,n �V��~�zU�������*�\$l�,�:�j5s]ݫ
��v�ycz�t���}��qW�փ(3�;��j����W�p3�-Q���j�C�X1�+����V<>�Ak��G]ɛ�L�1,���,~��/�U�z�Q3f=��,��;{k5��Q[�8䝰�~}���!����TSh�LR�E�ZM��	x9�����y�4��Uڅ��� v[ �4��B�5"�*)X�".�6 ��6���I4��Aap�:��:hbˉC ��A�o�Џ����+��-�KfXj�
v�m��Z�M+��f�H��0䤩���`۱�]1�嫵r6�:]�D�M�Y2���P\�3M,�E��L(���ߤ��
�u���!z���^��b}[�5�Mf���*�,��Ap
 e0�����B�Ѿ*r4瘪7×/������2tZ� 4�&=��У�-3e1j6�c��wU>�${ȹ�kr%v�\YJT_��랷ʅ\�� �H�(�G��^Q�<�H�+�d!��4՞���3�B�e�7[�Y�()��f�c؍�X�HM�Iv%
���D�>�ͬT�]��D��=q_�n���<�i���E;��o�hz4ǁ�=XU�|�DVwn�v�2AEȉ)�#6��`_i4/�G˽}���\�t@5�3{U� ��X} ���_���`[���\��vl��)��R*b��Ìԍn��ܨ�v�eUS\x�OB�˂_Ÿ&eo��p�����/�×>M2:ɕ=���^�]X�w��t�4g�fH���R�Z������}���ak	*>���;2mdL8;�3���i�Dy;~c�}���g��0H#N4ޙ��LY�C��'2��ME�����Q]�}{�
�؇-�|�E�-���������f=~x!X��؆h5.Y�חQ2.�U.9�cjk��SƳ����0�)�J=A���6hg�Py7��jyj9y�.uD����4�atPva��AvU�S���NN�@����y�e}{;w����� 9va���G+R�����^���j�T&��mC[�{9�x]���D�N]H�u�<�0��^w�r1�x�E=��L�L���Izk��0��XI �fy�o�.���~#��TM@������uv�f�Mv�v���]��SfP��1��#D�@�HI�-��jS��ݶ�\����d/a���r-a����N�M=~�sb7��̞y�L<����y��}~���7�AR�������<��u�3>��{+�ܵ9L�xZU��[k.W��oW"!������"j�|��U�Ӽ�e����GiQ?_j
����&c*� ��d0Y9��m!�\��C�[Q�{mm��mX���>�>�nL�gB
�.�`a��XH�zS �^��<GU��`�`����lX9��a���@m�L����ky�Hys+�7*q#d��&�ʬ�r�n\o���Ϧ���=��c~r-�ѵ[>_S�]�����Y�[������$$HYn:ك�vt�"zR;ϸ�4P<g�暵r���vցG�n't�n��[9Sn��A��:��.�1$���}\�}g�2f�mx�.y�L� �e*���l� �@�5C�~�W Y4��6k�q}FQx�}�ɾ��W$����-���P`��@.L�vT�ph�6�k6�̌����$)���[���C=u2����j{�Q�����ܪ�[���fØøh���#��}�P�$�9s�mp��d�Y�S�)��tÈ�y��p��!;J������� '��Y�ism`A\���ׯ&o �Wf���+���_���Y�t4a�C)���[�6L�ԉQ���*�����ڮ;Ӷ�ʬ#���#d���x��Zs����T����#:}xb�ĕY��Ί��ѽ0�m8*�a�K�%�p����6j=u�nyy�&�uk�;U���^��ﱗ)x�;�P ��jO)e��\jk��}�3q�@ߑy�����))�$m5�������k�N$pp���O�O'tﲜ
�X�m�� �o�u|�Z'6����(Iȡ��k��3�ߎ|Ϧ7�0WW�׌�Y�kYb�c�7��X�v��tnt���a����������׽��}�q�I�05�w#�y��3ܮ�b�^�U�]�t}���Y��ik���#���=���q��/c��1�M���������J_L�j�8Q�O�O>6z�I��9���st�Dڡ��ui4���e�h�A�\-&�(H%�ř���Fb�2�r�����ͱ�{�8S��W�Rq]8��r/���k��ыʞ�\���9��	�����ө�:����\p��Mz-}����vz�>a���Lb0;R�~��K��|�߾P+�8�j��즨��4lv�.��*��t��xwANXr�v�#�[η���������}�E�u�#'��<�s�`�;^A�৏[�G��3�����b�N�<%���L��n���9��}��2���$W�>u�m���D(��njŝrc�q*�� �8�;�7�i�VDf���c7��� �SzOٓ#�U�9wFD�8�w�sL;�p\`?�E�	��%�[�qj^���0v� t�7���'�w�y�a�y�s鸔MX�9S�J���S�\ͱ"���<�l��X
y�b�1}�-�Ϩ�7�t�;� �!�;�Q�Ֆ2����e��n��]���a�%\y�wKȏ���n|��r��T[�m�xgt�9{K9��_�y��{�|�o/�G���rq�^*��1�t34�hA�9kjb�fs�k��L�˓C���wާ`۠L�ӂ5�`�67)i����fm�ٝ(U�F6�B���8-���0��~�~�߿ZĎ��O&1n��������%�нS��`���rr�h4W��;:����7���ܩW���@`�D;�j��La]7S�ճMK~҆��Ui�m,����2�D��-I����{V&t��	��پ�c;v+&�ܟLl����tt8��(�P"�T*܊����bwd�싑��hw��̘Iw�<���Z�����3��f�O�h7�{�V�߮u�xx+w9a�C����u��;�+�׳����8��B	���E�UiZ�sl�a�-M����'kn�'�{o Y�
S�ѐ���-�ܦ� \����0w	���>��vUB�_��R�E஡!�UG.#�m^$WU��87��)�q�)�ZIZ\�;9#�
3$��(�nu��Y�%�by3�ۖ�Cb��a�̳.��́��`�dz�h��#���)j�������琗��5�L��k3��0"ke��-eݕ����3ے���	)]\�, Vf���0-�z�b-.��%��b&�\K�F�q k� �.��]z���y��ʄ	A������sJ��%��w�sσ����~�?]��A�J��� �u�[v�0�p4j��麻��:�M�&�&���jDg�h�홻�z�cqO]��w�/y�����c�_Tۜ~�S�̋+&G��y�"����s�uļV����h���(���@��8C��e�n��:l2�)�EP�#qAU��	�z%�Dџ*Vu�KΜ壱�� ��L���8��RXU(5���#�����lJ6t����Z	���"�}�T��4�c���f�@������.�wR�(|ϽԨ�Q�{=is���/̠�Ѿ��UC��w�A�a6�wr���q��t��(߬��q1��*�{]������~��w�l{d�T�L���ǅ���J�9�@��Nh�x;=���/=�]U؍%��̖eBN㰈�)����g���m�q�/�iB����mGV�ٞܺ)/�VnU�>g�!⭨�C�dԃ�.���{�oZuL�
f$=�����v��q��=�����DfD�P ��3�*S�d�Og��>���hm�dYK���݌��}F{�l?;�� w��`f�;D�?	!�#����&�Td Q[)>�������}4o��r	;��i+���.3TZ�����uU��U�<�A��	i�\kۛ�x�VW�@�%\�w�{ ��sjw�����5�p�u?Qb��S��:�i]tî���\�S[V�jr���ԉL��9�U�j��lfGYg�A�e�4���2G^<��+�f]��]��͠��Y��(v2�Z���'���w��]�ݙ�k.*=8�'��y'.V�w�;6b�'p˘Y��k��"n�on� j��#7���؆�L��j��!+˔��`�d��߱k���t�y�:��x�Fq�}-ݥ�z��S�u��,�M>++]^^��\��׋�_��y���O5��h�q�q�),ڍ�o�p�)�%w_��8�E��ޱ�&��:CS9�N8������Ś]f��S�Z�S���fZZ�=�F�k�{����aǭ;������HLe�ڱ^d��̽��z�������
�D6��m#�av�oC���xݶ]���:����v�s�j����m�5Nmּ-9+�Zn������u5&��s��TN���s9��`�x`3%��_,}$��������%u6��$k�a��j,|�PV�E�==s^nX�����T��<L�9�mKY]f;��^�@���q���s�g&`�ì����t-Z��V]f�LYM���z_>�
�����7�Ur�գd@��fb������̰����R��K�[��#|&�[w;+��̳?.oq,���bZ~9Oe47^;� ���Ӯ%X�M�y�����=8f�f:Ե���n�e�q�sA�Λ=]���;j�}G"o;��f��y{�8�o��_T�]�5Ԃ������j�P���*���W*�ɁWU�v֊� �� �dl���,�L+aly,�`Ͱ��,S�6�o4Wb�]![.�p����] �˕Vʒ�fg=L�.�ڢ0ґnՉ�;��a��bۋ�h=�$+XY����.(�@�4��		m�=���:�ZMX�������1���`�7c\�1�GjK��6(%�t��j�	fٴ2�h%n��[��)0��]&���m�T�J�"XWG3Kf�䡭ΓH5��Q�l�XW6[GQ�uƅ����38l������5��,Gf�,Қ9�f��a�%Y�����Һk�L�kJY�"�3�@��S7m�E�hi� ˭��$K�Ŏ�(��H^�\�Ґ�m�L6��Z�f��ZY�j���h�t2��y���[43'6�vH	]��GZѣrƷ��1E�Uf�Q6:��T��s��v���-�h�#�4��T�:e�D-n����%[��b�s.�F�lg��){C0!ͬ�&c� d��j�8���1�jT,+6^f�*Mv����8"�S)��qcm�E
j,R�zR������T�ŘI���if��%�������W�Fi�g��I\@�]�$t�8���J�	�ѵ��m��&��0F���a�J��6Zb�5L�M����fܐ��٤��`M�@�n�yûj܋(`l��У�&�Լ���K�CD�[D��5�e5��f��Mb��.�
�Xj�R�#�VgL�x�H$[�M6����9���2My�:��XW����"��m�݇�0�T�b���
]L���-�1���6hͨ�D%v�*�Pu��#p�%�j���Zh�k1�l����*�ɥMv� ����p�n�Rk�WM�f�`���-�h�N�JX页-��]j�K�!sz�� ��k�Z#���A�).h�kj�%��Z�b�cJhn8Ku�[�!�	������{z� ~������9w���0D��r(t _���&V��^��@�ţ�}�]�M/T�Q꯷z�S�S���=)-�`$��\R](���4�:�`������\�H�l�RL�ߵ{3T�����Fo���7k�l���*,�|;:���HV�ۓ;�W�0�ܾv���fy��䊤�F�a�@"_O�c�������a�;��Tw�os��"?�v�ʌ�n��w2�8Gc���'�v�ʷ�P�K��-]�W�B<ل�0����(��>f)އ�չ������1�|#ݝr����)�?h��E��]z3����@ڝ��y7�q�ȭ����棩����'�8n
�P�1G�[⢻h�*�6a��]��ǌ���>����tV�X�[GGy~��a� ��v������ ���ջ]��i(�z�n���E6�4Je��}'�{ {�߄"��a(�˭�^�����!�,�4&>OO����g�� AT:{e��²=*;6�ة���l^�t�I4���uzhb�c���M��]�^�F��Own$B�a"کO����Vz���_�J�]�݂PM,�Z@���ty�-��!�8M�CP�&%������˨m���,5f����P�w��}�,J���=���,ǁ�Y�{�[�^v���_�0z+���M��%����>)V�ۭ砘��#�&s��������:��`�v8�Yɺ���ݓeg����6,��iN�	ݖ�HK՞�[ˬۍ�y��U���6��;�Uu}��l�Z1��vg�3�c>�c^��_��e񭾼
bRb��H)��/G}�y�ޛ��zνN'$F`�ݤ�}7�`���T�m�|�gh^k�����M*z�Q$��x%�p:���J����9׵�G`��������cb�{3MA��{ˎ�2����]���i��j
)��U�|D���d�2�s�I��Dt��n��ڢ"zI�*-Gq�x	��N�g�3��<��()�ݱ����z�Ҽ����3�8�'a\�H�PR�v.̳e��m���Ot�����BCzty���9u�QC8�W�� ��(����[�=���
�}�phݿa�򪏹n��
�/ӓ>���
C EH�n�|u)�4%d�ˬ��{�>�c��v��~�}\��m6iω��lE��a��#��Zd���2�\B4�����6�����xc��vUx��]�W��d���J�U��"��	.��+J�c{��j�^�fv���uz�/�P$���0��\d�~�]����GoE��>��]|��S3×<��,2V5��E��ez���5�yʰ�N��0Gsn����ʷ1�V�Be�����SPWAD�0fE�,%�B�w@'��N���ao9�r���oWDJ�W���.xD�m&KڰH�@� �Nν�����5�Uj���:���,���cJ�m���	�@���u��<Y��I��w��-��L���=[wF�}�8+8>��K�.}�֮���a�m�-�ТGE��sh�d�*]���w�<^w���ӠO��t �;�H��F�s�M�)�������~�J\$s��=��ɥ2IM�f3V�x%�{f�Z��{��eE<ʂ������]Ԉ��{�U1���<W˞b�Yǣ�D�\��������3;.4[�u��͗=�T���c�����,1�>���a�>ٹ�߲�OmV�u�p�c9�w�k�d6�P ��0Ԍ�-�vb˥
�lWU��S�>0Q��$D��ke��~���Iӳ(py�G�LK�
�Ƙ��G|��^�7�Ŵ(���ӾunE�d�v��7���N�~���� E|$�G=�	�(�/}�J���.Og*�J�v��@[\.ˉ�'���HFJSO�j�x3�:b�W��d�K��	��%y_mv
��'Lt/�BC!\^��m+��G=���OSn؅�"�>�k�D�;W[���Yx#6\x��[N������,E�L_u꾼����ލ��!i^�ie��PO ��	8b���͕����X�\b�E���L�8��=��k�#;.n_O��b#��f^����fGv�`u!jLr�ʵ��坂�S�Q�s���k�h1p�[���H@�v��R+.���g���#�R��AP�b�P�������5m.&rfu�Z@kt�hU������:�4j h����Q!]�&j�8��Z��:&��&%���y9�)5Lg�,v���Rj�+M�6�[�f/W�[�ؖ���FSZq[(j����5�7]\6���7|��^3�-|�^�{T�4�&6�aY��̗@��m.e��������s�k�_�;vy|G��WNt�s�@��6R�5�����{��(r��	�L�z"[��(�"*� '�� �nu��j�)eȐkF��T�w��s�$ĜQ˭'���{{��N���ke��c��Y�xgs5To&l����t�����Ǻm\o�y(�|�0�u�8Y����*VVd�}����w)H,����[	���a�6�"jC6kG�]�W�`���7�+��j�+P���v�y����T����h�P�j��U�5�"6�\4�W����r ��`��mU��2{Z�n����z),�v������Y�O��
���!�"kˎ��+��ם�h�#ø�z�]w�k{��H�C��)�F�}�btIiX�foJ�=�{¸X�����4���6�uh{g�L��8�S�.&Ҏ�u��;/w�lo�=zk�.��ͽ�q��aI ����c}�'w�ɫkӪ��%��z�{v����}�*�3)^Ù�%�|v���diCƽ]잸��	�5���ɯ��ݎ*�o�6I(WTnt��j Wgހ0J��R�7�%��,)1i��&&� hh�����M���#��>�o}�cr��<!T�дb��uGZ�̴?[S�LX�o{� dr�����Z���ZY� nJV<m(����_ڪH����=&N�J~7�;P��g��F����2ږ&��x�<�Xbv���(<�y\b[�<�}n�<�u���>���p�B�V����P��a��ЏX����sђa���f=�px�|�>��Q�s4�P�ſV5'N�U9�e���}0W�\ �=��ns�s�ɭ�{Q��@��I1�/�Ӟ�{�YR`�dSo��	r�S�Ӷat��w(�/C��r���R9D�*x�2|�zEj�L60-# 3�+%@s���m�Z�S�I�
a���3١���y�=���K����B(���)��;��2g�1%g�j�W�1�P��Y��';;�'m<v��n�	�H��*�����0YP_���Z��|=U�/�W<N����ꋖ�׻�X�ׂ�`L:=	f�
G	���y�}�9S�WJ��\���_��\*�vM�"�ݻ�n���(hHZ�+����_�u��[�=s)�����V&�k����c�.F�yzL9Yr��Gz���nP��>����f��}�b����;��YԖ���E�	�u=����&�-��=��G�������a9�#�+�DX% �N"A��0�d�vfKi0�\m�]Lgs����Dt�������|��w�2���(Ȁ�Zޢ_�� ���9DQ睢k8 Pr�9�21Z���K��J�t^@����e��U�+!C�U\HO�>�}ҷ1�s;�#mFn���@�;��x��dP
�����p��T����Z�W>��"҄�^e]��AK��3u���l�O�P�_���k^��؜�\��A!�Q�0��wr��E�~��]�r�*���#g��F���
d�r���V>0�'
#�K�j���M��d{�N���9�}�i�]pQ�1�4tۻ���+O�a�S sp.!^^�߽���=Sy��VK�z���	�,V�:��U��������?}˷ֹ�ݯ���jN[I�Wz�%�J풹�uS<#F�2�Zs'0�ģ�y���wA��&KIM���A�؄u�Hϸh>Ϋz�1�o�WF��p��Q��I�6�d�
���[��w�ey��uq�w'/�ȓ��P;r z�Л���KbhAa���G�]�e��6a�|�~��mt��$g�7H�4͌
�4�%ibs�J���M���k�	�����M#��+��l�K�z���$}Z��9²�������
��׋��w��W�����a�97:����pHH��5��#�:��ufe�E�u��"h�I���*�ժ/�܉Y�����l�7����T?G���w����4}� ��؎V�Α�`�8�p0���y�ƃ&���z*矻�Ey�{i���'��3#���->�rD�'y��C:�4=fP		�$�71:R���	D�3�7;��h���(��U����6ۃѧ��-� ���u��Hr�M�Ԙ1���3b<,��.RfF����xx��\��M7Ͷ�L��{�.S"P�MD_�L
7;F��z�t�2#8��^��J7��I�:<v:$xϞ/=�F=�7[n��b�����\�
wr����Tק����a���*#>�)�I��>�������J�UuݛN���g&Mu
!tez+=�
�ƟN���J>��UQH��gS���4�.(��6����c�1�Vi9���*���1�v�Je�kV�mJe(7\ۢ]���BYc5���4~Ln����CǏ�~ƪц)�t�J�\o_��ܙ=�\��}�^y���f.�GNo�z��]�N����:���,�eѐb��7�	��a��iL�ڽ�v,�w���p���:�L��p�׹�#�Op(��qB���,�cθ�a�aG�-�W�����WC%B$&�bc8��?#2j����xM�ߏ}� &��$�q��/ǟ�����'h����ݭ�5x򺡀����jҤ�e����v(q����t���/�33��a���MÞfN�܆?Vz�MMo���h0�2ʓ���W.������;]�o���T��T�{��gջĦn�ٶ����I[WY���wC���{m\���k�\���w�������˩}��u��J��RH%�2�)���c�=1X��6)u��ؙ�m&�#*���+�.f��.��PM�(J6��@a�]����,]fjR5mIqe�Ѽm��;E+&�Y�Yf�H$�� 䮌�Z�Y� �:W%1���]]�r�v���U8����\˵Q��M#{U�y��tm�
Ӗ�6�	s1!+42]�5�5�L���БXmA<�w0�r�Ί�.&�|����y���<.i(!�}rsu�MB<4Yn�Gi���)�sc��{��*T5}XUQ���b{�!��E����ڈ�nWw&U�7<�o�eg�����+��B���'��oO��fP��0o*�XY�.�' Ua�7���5k��g]�B��i�z�e@#�]*�K6�ڊ<�WX�Θ��m������v����I����&��m��(�:3��z���c��N_���l�z��"M�{�e��	���姂ٴ뗻o���cی�ۅ�b����ZN�ݓg���v����ϣ2���GG���v٦� 9���e�uřO��<��C(�P�p�#�n��]�|�j{D�`L{������dFM��bm'��3q�0�V�~IϾU�c��nW��Cs0׮Ɍ�#È�� LtNi� z	���9����]��;�y�mI�]J�cWǴ˻����t\i��2�3�g˅I���ޱ�{yv��b��{�Ǭ���������xug�9|���ND���E��0K��髃���F�����\CKiZ�{�ף9���k����v^7.۝z�pu�x�'j^9\ooq�U z�l��6�8�]���R�\)���4�.���*`�;�wZ���.�c�jz*��vé��5~�:;� �p�9�������Ꞿ�(v�����w�����^�i����@gj���DQv4�����4��n��^¤3�	' ���힥�1�6����m���ʸ�.�h��Oy��)i>&�H��7N��j�M��1&�N�zf�;o�k�D��P��;�Zp	�ښ
m�*f1}�Y����q0��plI������G���N��KT9�)=qG�f_��*�g.�Hz}�Ԯ=��&l��(�@Z��`�B��e��^�4������`�E�ˡ�W�^d�;	��(�]پ��5�eZ�#��^�yT��̏{�w�1�D��b8D�٧����9 �I�m�Z�x;�a�Z���w�OyF���8�ngc6�O�d{���_�!:�#_eM"m^�1n�o���uSٮ�'��AA!W���U���[A�d�*h��Mhk�65�3��g��d�֗]H"z��p��$�~Ҁ�T�p���{o����\q�hg�=�95��5��t��9�꼛���PQE�	�r2ɿ���}�13|%BǞ����o$u����b�(in���.�`R��%�Va��G!c5�RV�a�q��{��%�8� x���</ދ�f�n�����e}�3KY�ĝ]��d5J������"�=g��3��i����I�ʲ��;s��9W"������:�ګ�VA+w�������p}v�\��(i�
����:b=�%/���	���FO�u����<���<3ٶ�j;�e�3��*�$ǾF~S:���zh|��C�g��.���`(M��Y����N�)M>��wؕI�v�	0��23�w����%�Qx�e1��v'�V% I��{o�U�~Ӟ�'����,]��6��Ӝ��<�d6$Y��j�7�=u&i�l-���|d�[9E�_�GOۇ.|��/y~H�|��23_Ӧ���ʗX�&���#�Kuu}qۼ"Zl��ED�0^��H{ݔ�.L	И�K��x84�|gbg�_*H�]��2}�d��]q|z��������m┺y=�Z�+�"8�L�؏�d��d6)���^�q=�X�{��z/��s	k��p�5f�$�q�$�2SL��2V$v���]e:Č^Ժ� B<fox��fF�x]Mw��ǟB����o�<7�n�Y{ѳ�Q�w��PwGrʻ��G��� �a�bU9�f:C6���p�����L�K�-��ϻ/�ˡ�8_�����=�2M����b6du��!g��U\�	�tGUWD�����!��i�������B%���m���@��ޢ3�l4�wj�$�F��+�	"ͧ����v��\�U����3oy+�v�}s�ú%�M1��`����J �`�J$Br��6]"NX��}/�t�-�`��'L�e+�'"���m�G5�s���f��p��S&�����c$�޳u&���'k;v��u5��J.��-�szK�:�wwml�W��oq��nY�����|�X�/�sչG��0V�5aGk�%���E���YG
�/�j̣s�7�Z{a�3Y�gG��*��qU�Q4���G��]^-M��F�-̘]��J�ռq�P�����G�ve�gvřj�b���|��$g*O݂_4�)m�n�8	���FmA�(h8朠�Y��L���	�i����[9�*�!?��ӕ���M l)|6���c�z�v��0�w扫G7\�p��t�aggl��㾉+��Z�5m�*��I�$��3H�}��p�:Kd�kuVhU_
Dؽ��o������������C��I4����J_K�gY���t����%!u�Q�Y�+{a������e���ւx�]pAPNS<F�j�;4�
�d1J�uݮ�
�i�Iv��V�P^���&�������357"�]y'S��&wM|G��v���wX��c�^�riο�@�ϙ�r̎��v��N�L3;\�ܦa٣�����N��2]�ڸn�~{����UUUUUUUUUUm��e�m�=�ɴ�TL[�k*���'`؄P��daw{�[��xHm����k�s�����'��mO�àr�$�@���K�U�׹ �W�T�X|:���{�9]�/1�rE��+���[��0Q�)���Q�J�qK.��'�e�8�cS�>����o2�?���1Q4��+�Y�'�;�ܧHy/vG#Ƴ���g�v��Љ��*p�V�e�J�
�i�w�K�s�S1�,�tzWW\	��-":��e,7OL�g���<�F�򨻸�qQ3hv~��*�XR�3&ٰ��ʍ���&���t���I���~'�{����Y;J3�sՆ��J�G�d������8�t^ǕӂI�5�x�7�#���Y��l�p�M�~>��I�<������vKn�����ܣ �Nq��,���蛑]�~~����e��s����ثٸ��VC���0N_rЉN.-��(b�;s����j�ϵ��^��̜�g2����5Ƈ�S�f�+ӗ��q������"���q���e�r;�=	��E9�ý�N��YlVӅ8}r�]�oM�	��!z��^>�S��I����S��{�ن;^�о�FWM�tݣ�3�B;�оЅq�h^��qn�L�鏚X��r��:�"�3��Eܼ@�eu]�U���h6�D�b-�b;U Y���ln$Ά�m%P��@��dדucNԼJ5��f��,c*Ym��FZ��޲�%�TQsW]l&��^3V)F�l���Rm"u�Y�0붚��ii ��tq���è;#�]˙�\�,f��8.f�av�h�K+\P�F�-,.�i��ݖܬU�6���f��.������4�$��aq��	G�>��Ϭ�g|]�3�}l۝W���N5����jw��&�$�j���h�5��b������n-�#������ڣ��n����N��"� ���:G��r}[gXKѯ+���9��h�Mf�7��^{�"�D)8!o�il��ճ/n��g�Jm�uGdx/5���C�p
��t�[�m�����R�]�Z�v��0M2�f�1q����{�h�L�a74c�����n��,{���ՂcNd����v_���PV�z�e紑�jM�p���)���͙{������]�]�cR|Nµ�@��Fܛ�ޮ��lc�>�]�SᙫD��z�E�x�l�d����B^Nd�s�d���P�|~̼a��U����n�.��M,�nצLģ��¯��Y�@�a�G�}�S=@�Ӟ�z�/�n��^eUZA7%�x�}�cN�i(p�E4]D��%����C{ަjX9�̧�:�)z����vڳ wuf��CHy�/h������QA]�ڣŊ�E)�{}\��{GBp�p����4���2r9��wAG�z�*L��(w�<2i�RS�I������[f�V�r�:���5N�dM�)�^\��`�ל]�Y�f;�|Uދ���Y�?^��f�����w�;�I+뼽�\�t�%��U�b4"�	���CP�΁!��t|%b��"ڃ{���K��p'��/M����yUs��v������k�h��A.�Q|�A.���M-F�V�jj�(:�։�h�#\��g��O~ϙp��<]����x5��Þ�����]U������>1�e r�s��/�O��r@����|$�ن��Y�Q�/l�����w����(�pU������s���`���*�c6�~�Ǥѳ�q�ޕ=;Fz��i(4&[u��O�_�}�&~����y���A"e���[]w�D0z�0Ȅ��g��,��Al{�U�f����	�l�a�\��q��$]{ˏA��E6 ���k��<ON��~�#�lI1o���l�3��j��w�xp0,F\�)���P%���ת�I"f�^W��j|�Թ(�r2��5�t>��ott���d�2T��vQ^F9+9W_�Uƒ>�Ԃ�g��箪�<��gw�W����ΨA˳��ų}<��C>̓�#	l��ꥃJ�^=���ש5��_S��?���~�K=umN����v{"`�`�K�mG%D���"��eĴn.m��F(*�ύ(�޺��
,��΀
ӝ�b�u��-���S��w�A����U��Mu�����V����z�VU�X*Z��jt�x��+ky�m�K�2��
� �r�/7��γ�e\#�$�� [5���V�T��b��siH�S���j�'��x��ۼ�=�RO��okb�݄�s�l�3�㳙fM��7�鮻�d��܌(P�l��j���r%��zw}�LV{}%{�#`{�Ctvq����nJ��3BO^����9��dH��.'�G��Ñ��[S��9.���˙ͩ��٨]zwI�p�,� YLǥ\��b4<�ӽ"}�_f�t�}z�[�������:����-�3�jfOz�9��":yn��-}ˌ5���m����*�a�/2&GK�3�oT^%@�'{�k�{��w�O���GM���Θk�fy��nY���c�C�z���~	��u��7	Փ����h�wyHN�ʥVj�~�-�-h.9�P����H&
p[q]Wk�2��݉Fj��+w<�Kx��F`����&�[;���s�����-'AVj�*7�REF�Xn�3�57�+���&�N�T�q���Kk\�Fn�u�P[d��uՖce�w�f�W��$O,ڨtyn8^Z+w�u��`N�G��yj�����]i�*�'��9��ʙ"ϣzz�Udg��7e!t��
GE	��!�D�l��~�W�� �oK��F�ʥ��ϥ{��f(�Fp��@]��]G��P6U�1%�t윘BoF��))ձ�j�G������cT��giA�/����Ւ`@���5�S��cdkXG׹�_yW��eȬV.�}��s����4�-��G{9���1���s���g����0�zl�[qϳ�9S��Q��g{jӔ�jB�L��v[GU����<��{�p�/pC+��6���S��/��]��-�T��u���'��;3��*{���fA|����R��8�}
+�ѹ	��lx����u\tw�{����9�7�`�ПQ٭�Z^������{ɷ^�p���@j*T~��[���YMv&����j6���Q1����r 	���{]rz���0=KS��tٕ}Dr5׷����#ڒ=����,-w�=�1�᧋)�lCH	�
6���ﯢح_i��8TF���Mx]�Đ;�����*�rԌw�*��-�A���zL��;�ڜ�v�!T�}��&���AF�u��٭yD#�H���+� P�}��c]�:�xk���Pqi���n^gX׾��.y���~�w>Ͻ\P�s�lh\�{�U��}l���-�Q�z��n�Un{��!4�p���ѰFv�k����ja�����QO�/3���Oz�}�nV��m+�h�l8756���}æ�}�[�&4ɗ���M��p��$.���A}�rU��r�m%�+����Z�8dZ�L@6s�ګ�)R..����K�p�`��؍��R��f؍`H��tNl3\V'j�����k�\ҭ���h·G�P��T��B��[3*5�ݛ�7Si3F)��],��mkR c	��-C����4�n�'U���h��0����pv�%�ec-4k���=�R1l�b��AH���!a�l{_��O����J%h�*ydک�Xae-��US�[�9s!8d8)�L���`��y҄Ǻ��c~����[�O�|�yV�_��R��{)�]>��fw�_vxm��.���T�:$���1p}��WW��x���4�`�ݾ#Ӟ�*k���������|�7A��z��!p#$��gj���:R�A���-�FJgV��3h�e�>{���� >����9���V	���������.���\<�>7�"z^U]�}��>m�@P�E���{��ٽ�-{�G����~��Aath�{Xd5�=���Z����g�2p;'M_	4c�+��'4裉t����r��@��P^5`����$X���r��m:z���w}̄M�av|���gzD-m�~��{��������Y�˪�`�vm1���o�k�����"�x!�:Vfd��Ӽjj_F�*��@J�7���h����j��Ȑ�
0+��^��xj+�O�oN���4����x �h [����`�Ǘ�*��{=�kB^$5O���\��u�M����ĭT�=���T^e����-�$�rU~�����U�����M���imHx�ⅲ�΍��Q�¸���Vs1$�7:i�<��vl��S1��}�Th_T�z$%����A��̥a���?R�҅O(��R�h�`��H�˶&�	
O2:�e�PT-޺^t�㊅@BE�`��D�U�B�Bk�&���5e]��M�4���!.�%o7wܻ�*BufI�.�{6k���4�ۃ��ݶv�M�l���<c�uR�E\�v}��sL��l4.G����1ਬ&�[�{ ['��}^\���j���r�Ә���%��jǇ��}�+5�2�;0�iL���r)�J%�	l.�
�v���ى�F��!~���И�c�s{��K/:FόDR}�"��Qq~�;˙��^:���^�F��燾��a�8���9+=�5�A4���$�[���r�T>\*�4.H����J�-�B�c�f�����u��BN�c+�1���ۯ����B}E�ɺ{z Z�%�aBI��k4s���5�~F;�	��nyp��z�e	���5��#�Ճw;k�2���9����m��U�Gv%nJW/�}������$�-BLt�F7;�����d֠�p���{o��(�a��(�9�a� �ٴ��[*�4lu*k3��̕�Mo�,�Y�U���,���\Û��;��)��%|������S�;�^B���4/�5yV�2�A
������5u���n�L���rWq4�Y��%��X������w�%���s�f��	�`6	����3�����7�y'�W��~�oL��`|�ұ1�;c��w�o�ެ.}~+���gI�^yU��Yӽ�6���ޭ�m���-4T�S%�
_�ll�y9���/E0��.���p�|���\��[�(��­�_j��BږB���}34jS���p����~)�ʝ���ݬ�核*6��:/��rbr��[A�Z3`����s�'R��m�&gӳQy뚕���:��^��_ΰ�*�<�g��#�ue��f�ק{���j�N
-�VB��9۪�����\�U?�/9�Z�u�ί
�'8�\�Ww�	�kq����7<&|���L!̈�q$�m����$Nw��栆����������]�3�m�{(6[�a3,��>�~�|x���(	�hkp��h��5m�V[��bD�mHۊ}R�g3�^�wk����k�G���S��Zo��%j�]�����=g�*��]l�F�-�#Ó�e�����%fZV&�f��!�W��B��| _-[^�Z������r�q�d��>�ɏ/g#t��rtf���E���,��l���
(�6Hx\�ϥ�h���{�n�p3����m�?D�_UӐ��y#1�����̽Z��������N�wEE��B8��A^�m����<kO�ff�6J�ܷ�iX���=��|�}C½fRٹ��V3�!�W2��O��D��%�R
p8�w�;#��<��MA��"����mG���`�7aߥ����ks$�Ʒ"�����l�-����.J��N��e^g��hE!AyN2l��I2nrQ⽷��+Y���f�=utX>CI����bh|/�,�s�F$✲��ϫ3��*{2���;�i&INvG:���a,ݪݮ���u^����<m��$(�laA�D44�[tcY{��[�'mq�*�8��%��m8$��ݐ��|��&�����6�EP���V)ل�l�}/��gd�A��M�tN7���ǇX%�E�-�dO�O�԰f�����'u	CN��A�!�Wit�svEV͹��؝=f�3�=@'W�jm�UŢD-;�
�/0O�l��N2���r4H��n���}���:6�t�����E;��/z��R3���_D���=���hwMt��(��k��vq��dq�⳶қ��A��HZ���zQ~Q.�q�mp�����^!��]��u�atL�	���{v� ���{��X6��Y��e��{}�⺕��,n��5��4�L��������u���X��WiדJxuZJ�Ur�.c]]+E!.���P�4+C������۲C9LY��ۂ]q��
	Xf�:\���Rb�6H*U�m�D�6����B�`<�q�����s͚�`�qs�l\Yp�m.� �U�`:3K]F0��cH��B��+LP���D�U�6:��
��`굨R�Ip�b䙗�,ԥ%�]Zh̻\Biq���32b��~��Cp�O����]�5w]�#�J��0�=^�t�lXp4wj9�R�_v�Y��Iڳ˰���q��}�W���JWY�S�T|����#Z �{�x���şƬ�U�t/|Y���ř�����4�j���׻noq�M$��������DA�O̓oΔu��m'�L�k��a�vٸ9�B..�qf�u�P����Ģ�#)D�l(��#l�7y��GO��c'ٞ�3l����)-w�	ˎ	YW����C�`�����O���>t�출$Yntv��KԦ�.�ۮ�q��UR4���wf�`=��"��׽Tǉ-߀���?����:���F�Y�n���px��ڹ@�[$���/#2	�G�<۷���&�?vh=�k�|Zj$��T�+;��&�˵�����l�T�;�oL�G}�����Ù����A�]��8���2</u�k��
�J1"�nmJW�o�柾�GkS��=�\���z�'�Y�a�^�o;�3�#~�nQ+��U]Rw��EƤ����{�����S�ŋ���Ɣ���Gl��"(_����}~0=7�½�J[7bh�����
c�z�����Ϩ�جbȎ���f;��0�J���a�0K%f$E��-�?���P���U�5:�u��7M�MvV�vݞ|�w	{}gX���?��k�ڟ�z�69�TxJ�����;����S6Tܣ%�Vηz���v�ɰL$�h9,D�9��9�}}=�`6w-�kJ�6��=����^s�Q5��u7iVՄ���՝���	��3�WZ��ї��y�Q�P���� ��Q�DWd�IcW`=P�q�U��k^S�k��@�]�t�]|�BF�q�%�vq �M6T�e-�f�s��w�1{ /_�,-]�;�݉�!���xJh��W:�,l�0���+��.�\���o�'V=�0��a��ٸ�hz/q5G�WnTB��x�]`F<��1칼{@�ʕ���>F�l�񺈣�7e��݆���Y{5�:=:�u�M�D���;���n�%��y�?,�VŃ�\쮢(v9)��]",57�t�z[�Á��?e�C��Pj�q72��@W'���s���Cl��U�JP`�q�7��iK�%. �$W`w���j����T�u5?+�P&]�b:&K���xP��{��2�c�z�?��������u�_�f6��,�kv���o�F��s�v��%7�<��D����whƏJ�았2�7ء]PN_mb�R�EnT�����ze�yN��u���po;��<�AP'��\��,��X� ��H5 �s�
��IY%J�I +�� ��*��l��ET2l �᪁�Ub�����5��U�7k#]��8!�e�6t�%B��,ف�ƚ�m/	�ٗ��&3YJ��GZY3\C�FbiZ�܍�2��q�e�R�փI�e����f�L�gF4Ѐ��̻D�;U���v�1Lي$�s!�En��U�uc����#l�`�5�XA����5��̭�AtFSU7Z��f[���fE�jY�"�����1�̣�гd(DÍvl�����w#K��G��&D�$����uŕ4uͭ&J�k;I�[�jY��-�v�"��,4IQl�ijSW1���cMGP�u(��t��9v�����&uջ\ܠYK��1����̰T��2ڹ!k,z����ToS��\�һ3G�YQ-t�i�F��@Lk�#���g�l�e���A�YQ����"�[��b�k-�<�,qy����Y),jR��Տ��M*f5�ƅnH;d�ZC&ܖ�c7\&Hf<I�Q�����2ْ-X\�K+n����;�Q�g4�	#
���s2K3`33F�i(+Q��"ªƎ�5I�V��Z�BX�GA�Kn�L�-��5��bb��VXB�Wi��4�%�@206�z��V�uA���YUхծ���RiQ�b!�Gk��j��y�Psa��Mb=DRb˹iq,!�!�ڑ/Z8*q�iP0�"L�(M��5+��� k ��7S\��b�,��f�bݵ�R��<xCM�s,�eB8�c���
��,5vHk��,
�ٸv(�f���+�������!��.\����&��x���Z�X��;Sgh�Z�
v���$h�[HF6�Gf�놩a�$�f[*�Yb�ά%a!�����z�L�j�S2�����ph���c"��Ѵ��ɫ1F38ln�s�2��.�G2��`�V�=��R9t��ɥ������fЃk)e�.�2���l.[j����O6�M���
�p�G��217��O�������D\�0�Ey��Xv��BG��m��с˕ͯ>S痮��8̴)�����P:�*���8e&V�`���v���uݰ��M`��3��� ��*n�I�ު�CL�.4���s�;��Px��n��mc-#�|������&	�����5���k�Dcb&���=Q,+��V�.~+��y=7&�n�֪%Jܙ�X���'�(�{c=�Pk܂�{Z�K��x��92(8��>��Z�oG�	�ˆ�6͑������"�2}�##w�_:y��7m2�	f5R�=3����կ�S���}s\�V��S;ާ�z�=���6=�uL�>�[P�!M����z�!Al2N�:P�F.�z�]�H�����l�
�����ۙ�c�Ʌu�G��H��k�\ʍ���e�	�:RI�
7�]���v�İ��h�x��z'x�u����ȃ���3�ؘ/3�4mj�4��r`��GT89�^w���Rʰ��<%dwy(:a�'�ڻ��l���+�M8i�iU�zZ1���ʅ��L'�L����0����)��
�KHl��&!QF�o�nmnG��1H��7��]=(B��БQK�,������ȱ,����<=Aֈ��cV��X"7��M5YJ���s2�X�.=R�_�z���}�n��;xҝ3.���D��8�vf>W�U���U�y\�i3�o��/8��E"Ym̑(Z�z}��z���D���ݾ��Wd�.o��O*�ty8}����+>���^?��^�[��qUTW�[�@��׽ä�[M�M���s(q˪��ɝ'*DL߉��*>�g�3Օ�0�,d�~��?���L{�E��).u�'e��ꎁ�kӪΏ���x����.O�h [��^m���s���yұ��{�7덟g��-c�zW��%�b��D<��vG���_-y��gD?b��o�5�����pA qH��693(s`�B/ïO�MWu}��<j�M"����0���C�c���ia���/`�,�r�wy�ɍ�D:�>3*��ew=
"PV� O�r,Y�X��/��
���ˣkZ�|eG��V�V��(Y��t`ir��f�*l�j�i�en�-���á~o��Ͻ��N���W��=�m�oZg�|kl���݀.��?�����V5���Ս��dm��6A�w�%�g?���^�/:�2Γ㈿��	�̊��������j2�soFJ#�)��L�F�GzUv�c�>�멚�e�PZf��W�?A�+��w�6/LYCD�
��ֈ���&�ٝ�;d�]t �4j,BGc��hd�BD��[[�����N�w��~�e���鼗
cgzr5>m���4Y�8(t�mW�=��9D��ɗ���+��������+��ޑ����^r����9�}���К-��}���]�m�mԭ;��	�(��TӃ~�w.3���P�ħ�gc�A��94("��=���v�3�U�U�~��>G�@Zp�PNCUj���MMN�q�x{��J�7�|m��0��ګ�ٱ����|�z��^SWs��X���m�����z��B��b��>�����a.0i�)B]N��c�;no����c�I�� x��E�	��֫�W7	f��\��,u��Ў��ld�=�X�n���Í�}�Wcl��q�}Bz�]�[��=Zr��졕t����:�U����g;1�{ݩ9�Y��i1!d�M��3Fa��\�Sz�,��!�Ea�ɺjz
7��tN��]�����w������;�U�ٰ>������~{O+7�K�ɍ��Y���]p+o�9�y&�v�%8N�Q*ov��RO����|�^yDޚ����ڦ������'3n���<s������Gʀ&�T�BXt�'�M�x/�uC� ��3�H��t��<�فpJ�c�6�u���'K���j�v<�Sq�j�[FI�LsE���&f��!�ȹ��r�@T��k�I	U�*�˨Ic!��E�v��#/]�.�4�4��9��2K�ڰ$^V�ɛbےR1 �1�l�V�ƌ���0�]�{pYXR��e�C���53�	Q��Ƅ�(@����۸��z�æ��[������K,Ҁ�Z�WSi�YT�1���Sb��)q�cv�)Q��5���޼��b�
0�45����f�H������i��(��f�D.�[�ٯ�����n�<,�t;�>����8��I^VjEnv���l�	����5��+8S<�tF+=�n��P�����%c���g��_fa�6�Z��j	>5���v 7E7�r������� �	@mҩ g9c��'ӱ>;�<|��!��0����f��5��c�A�V5��5�vvM�V�����4X���Bi��J�=뎈��������O.{׼j�?*&L&o�3;��K8�4�{�Q�]�� �`A	2ҊB8Ʃ^\���-��ҝ�v����陡w�쬼���)�C��[����O"!�s\���K��ϛ�lnC�뾢��n���!�Z�S�f\�z6�=]ˢ�+�b���@�Ț���/g���;���pKU�Z����Te �%��gM̞�Yi�.QC�^uyЄ�TH �_J�n�,\&\�Q����w�퓼�5c�{N�1����-d�W�L�͛�޳�O�(�_T��ȶ�����(�x�����E�e�Z�bt�`zg��R{�%\���M��Ϻ���V*�ݛ����;w#t���J�ܑb�ہ[Y&�Jj�ڠа��mc�
�TV7�%X��YS_l�x�Df���0G�jO�2nm��<֊<�*�2"F��<��;�cK,d2ώn*���ת6�^��U��<�HI�[ք^ύ�׀�L�І2�^��BfW;n���2�\=�0��+�{z����8��4�h�n����"3��5�Ig�u����?�!��IW$〟�����G�$����j�A1/��j��w���o90�����:�{�����j,V�	�t���R�����ݕcޣ�Q��ٳq�G��rG�Q��o6�}�x�y��*p��{u��!�h�-�W
3�Ù[�L�Ww��_Xxs9yOo�E������2G��"�+�0tݰ/�^���6;a��ZpYE��!��mL�r�<��crZ�گ���#��'R���R�à��P=�z�P��_ĳez����B�Xx]��^��g���(r8d��&�RtW��R���VT�Eer��\N�Q��ۯ2p8R�;�B�%�S8dq��[�.F�H�W��a���-�Wp�2����J:�ܞ	�#b8
���/qk�Vﯶ�qԈ��A��u|�>�O��Z�}y�u��HR7HǴe"�`�!	Zf���ڗT`b�B�D4�{xUsڻ/�H��92w�7p�-w<^���yɞ�S�������m:'G7�%+a��V�Ą	 ���0�q�p�*2�^��v;� TB|)�o��ҭ�u��
��+[U�L!,��u��؝�n)ޯ<�$���G�c�,�p��o���T��"5�{5艞Y��Sw�~��
�¬��j���oA�{~�нDf��q���mo��ܔ!W����P��: �%�
���0����5���O�$[���꣝�"��R#�������,;���}�La��Ǧ}9=y&����K�>��'��ҧ���]1��N�d��=�&[&m���&�ږߵo���3�#ݕ[�S��jP~�]y�7*��,x{mGOa-Oy�7K�P�a��	`�2�<������m��J
3�yG۳�G��e_o���tB�\OC�Χ[���^�5'��rU�y�v����K;}�9i>�>�jn궽ݥ=�	n�c����s�8J�N\λ���#����!&���|PcF�s��~��������t���>�w�{&��$���])5����a4
J�FV�i�m
E�u�V�B��M�~�}�>����O�c��hݺ���n�����M����]O?fܥ�R�U�&<W��*NT�V귑�\[i� � ���Qa���M��d��Z&x�4�<=��`�'�v�P��ǟ1�-X�W��&�uv��"x������TVj�P�[I���� Ѱ��G+��d2�f�u�
�<˼���0�ӶG ��S�V�
庰h�e�ܛ�;+��	��B¤d-��N��H%�s�z����]i}sm��[�T�b��L�:%ݸ��¨V�5�D3�0v�z���ˇٹ6��]_�2����/Ok����i�6�)C��]�w�5�°��N	/��b*�ٌ��]Uu�n:�����=�#~�c3��#��y1�pt�2��8ލZ�6Y) �7}4���+Au��[3��~��8f{�8�ܯ�R,�߰�������Yy���y�o2OcX\C7C�������)�'�x�3D�Zk���r}�\�0PSh����q�^ �2��8!��ezvKڼ��h�#��w��f�͡�6!��̻���I�^�6fZ�5�5��JR�2{%�N��]X�ẞ�����T5^Ԟ4+�Q;��e�u˗��v5`'C����A�Qj�p��~���Q���ΫUgK*}���M�#j�:1�>ت�H��m�p������z��M\� ���y�s�2�}����A2a��X�|+3'���z@��Qk`���c�c�ƪC\��1$���)cki_Ed>WKcN�w�&�'�<4��鲄�E�>��nd���|�5��X&o<���؅/nu�n
]�^�*�������U�;��U>����w��+�	~�ג�iT���k8�*�n���+:S��7B�dz�Ě�dL����p�I[��&V�y���q�ê`�L��b��Xi����])�v��LX���mW���t*f`�fW	�$��`ճ�Z�V��f�43*,��в�zm
p��kl������\��4V*D��-�a��1Z��(�$��u.�KP�k�,��0����59u�h�Y \�)�SKĩ�E���1
�	"�b�	zV�/�wxM�ݴ*��BV)���Ώí|�3�u�t����d6�n��`'2,��~� ��qa��ݥB�3��\�p�)����ë^nu5*k-�l����>R��i� ���<()��.����:�y�bQ�^�����(��j��nd!��*J����*�a��}��Oq����i��:���B��.͏a����X���!R�,X���*��9�OpޚL�>˪�i�e��]�-�������皙���<��C[�2LvإU�����I�$A�P�ϔ�9(⼺i/q�A<��4�F�2��Ǐ��6�T׹q�� ��,9����f�ۻ��å��I�g;�u�!�~�|�?�P�h%;Q�|eFl��=[�r����a�
�P}f�7�;���O�+�t��Mxn=�B�=�.��P��ӝ�#�ֵw�������{<k�_��-'�L2�Z�,��O�=}^᳙9p�4}w-N*�ŽR�yw^���ˋƴ�W�m�6�R����Z��o�=���ǆ:�H��*w��:�{Q���B���:��s�g*f7�v��QC�Ǚ�� K��W�3�����yD�=
.}f��I#7�l�[�\Ĕ �I]f�e�gy9iuKyӱ�+n�{�����:���*Q�-4�ӥ�D_q��ʊĘ�'3�e%;h��|�|j�q�԰����I�!�8�9�NfD���� ۹bɛ��BA��%���Я�*�Q �p�? `�LV���*3h풗6�M1�G�s��2���__B9��uh�;��"�U��'����.>�s�S��nR��J{إ;��|���(Y�Y�#"3'LU��ғ+/0����K�)`<�^�O�xaVB\tf�Ⱦ��aW��9��>���/�#1�9��Q�:,�a���8��D�J�Q,�!Gg;�7�p����ܥ��ʿq�.f���W����.����X��Yb�f��<_4�� qچS�<|��˪�]�S`��
HP�ي��u�䗁[Y�O@<:�sꛍ��e�w:5�n�`��w"ҕ׆�R|'<�Uc��̹�U��;�	$������jn[׹]�eCw�h�h��$?mtj��l���᯷1l���(E��n��:)wC���{wՒ�)f�S�1��c��K�=���I�`$�_Z���\Mz�hp��Iz ���z��H=�H����RX�������t�M�vh��l�]�[�uh����A	�0�(f�,��*���5�X|uP��u:�sܥA�VWW%i�}3&0��0I���>Bһ��6C�R$��W9�A9�RV6C՛2)9Ș���Oބ��3��V�����/���q����42䄉!�������*B�Kf�Ɔ��<dW=��L��j	�.3T���z�a���⺑�;�q��k�O�(���y�v�y�:���,�Ӱ*��,͂i�{ƣf\��Ra��7>"�;�0�}S�~�v�]����a��=��T��qH���׏:k=1���g>�\���'w�׷U$�{�ԏ�+��N�;e�i�I�>����k|��5�}��������� ���r�z�lT_�a����K�#��u�٫<�{�__{*Gw�0S���&�����X�3%)��#hFY"_���q��Bz57�xg��0!�$_A`�wJgs�(�܏t�� ��/�߬qիwQ��D���W�j�3����H���Qo�0p��o�S��Z��[��_[ǿ<�������\`Z,���݉v �W���J`�Cb,+����a`�I��ș��\ō�P�%�Ċ+�x��;F2���um*�1���F�D�+y_n,�r�'7'5��R"�F��|���̾~�M���񗘳�T��列q���dāGO���������wъ"���|b���xB���;���o�Q+�4�p[%��2���|���]����ᤨ-S�;>r�Q�g�~������k:���:n�b��m`���]� ��f������A
�k����kv�G{���&Nt�����z�:�V��S�8��+K3�����;Oj��̺��̣y�������P5����ٌQ(utws#�m����r�������*��wO󵨙��7`ѧOxv���mgq2����Af����$5�m��Ԥl�8ȵh�zQ�˫�z���Wˮyפ��nK��!JS˷[��5����^`ε���нjN�9S8�̴�;x�.��K�[���fp�d��6��Y5�*�`���ni��YT��Y\�ˆ��N��0��锩�葇/�Y@S���m
L Yq�]�H�0g,�[LB�It�;[i���o���k����F��JU�$ZAR�{�i*�4(��Bjƍ���QG	"�5v��z��T_l\��Ş���dO?-�܅7�CS��
�3uZ��'��]����mk�B��{(X�"����R��V����̗(Rޜ=y�C�K����p�/�/��Q����Y�:��.�h�̻�%�n���ՙW�:W�+&�ɕ�e ��ȠR]Hɥ�ôd�$AY�Ӊ�����YEGMq�X�$��3�p��<��gwsU�[�]��Eo��%�/+(���*�%_q�9�2]�OcyWLf����p*9��>��t�e���u �w���u;B��ߎ?!�/��r�&u�5a�J�{��ё~x|'矊�������������sT�n	���L�M�}ؕH��cl�5ʧ����Q4FW�k��'�~�9���g�we�lP��<�m�U��kGp�i�K!�h,a��.�zH39��Äou�5�]]���P\��j�E�������>/�v�E��V�9ɮ�Y<3i�d�ZW �T�K���a�]}�t�㈄�<�����8�𶶫KZ��>�W�Љ���<R>=y�&_.���X����3�>魊�����N����=�v$ �{�{T��w��&�,��W����+y��:H鎄��^&�7�8(�jA>�cH��#e��)m-�1�LZ����3@�Q�aa��#9��k�����[�/S/Py�S��ٮ?b��3e�>����qiz[����g���e�ۚ����T�G9
͈�z$��÷̪嘗��n��$+{oǢrpyS������7���ʂH.��Uyv�3Cd���4fT!^^�\�.v{�#;ݩ�"�pM�B6u{��P�U�cq<<��~��ŏ�Pڟx9�J6G"�s�7��zz����ڤ�����t����d��:0�O�z��_A�ַ�v"U�w��A(I ��q�;9���{�Օ���?Vx����a?znh]�z����������m;I�٘��º\��I6����p[<$�n�I��Z!�c{*���│�}M��Ё}�N���%UEWU�kV�-o.��\ۦ\��b�S�MJ�&ȷVƣ��͑W8̢�W[R��[,:�:�@�Q��P�vI���YO�����08�D����$ٴ��(�GP��\���aE�Ѳ��.@��e�k���n�-�L�M5P����(@J��HX&��%��\]�duҶ���8��M`��#�pkB�$]j[�Sp����ã9�~�nm��Z.�^�=�&�nuN5�����Fe�{q7���BKHD5��싁8�V��3��y����9{F]��<hD�d�n�==���C�/���3E���6����79�XW9>~�I�aJ�&=��и ��_�R���g�6�l?<�����r���k�7VL�h>bH��5�R��˅J�&�e�)�i���i���ۂnǧ��}��8u��!iB̭��wB A��&̯{71X=�&כJu��;�#۽��ŭ&D�q�U�*���5���;6*+��Z��/o�T��꥾*n2�:t�i�q�YK7�f����W?gdKƎ��|��<�G9KV�2�,�C%U�O�,'���nL���ށ9 tf
$���~y�O��B��#)��+���=�ֳ_q���<J޳9�q����w)M�R���<�L2�"�eQ�Wa�OҫϞy��}�m5��宛�'�w�\�$����|f��v������������:-].��K���y�����Y��R	!8.��^gN�6��E�;}�g�?.��>�����ٳ��[�/��+|x�n�Edj��q9�Bݝƻ�=��n��-mY��̖:�q�л��)��}�"���i0�O����nķU*��)[��1�2*�W$�A��O]��t"Q�!�EA	'�Lo/��M(0���MW��+q[D|��0�<y<��F#ջ����)+��`�Q#��U��)v�0�E3M"�����R����mCv#ө�tm4���,��zr���+�W\Փ���g������x�춟�x��VIV&�]�uVIOU�!o�>�X�녢�u�P�h,bʤ���Z�T��=�H�Eٿ{w��;�2+6rp]ձ��κǼ�j��6�,'�_x�F������k^P�E=�w"X���DO;p�}���oAv�/f-��j�`O��������X��ʍ�q̿L��c^�=c8.o��i�W6�����������u��c�B�nr��]��q��=��G> �}k���G��L<�ƞ^dRx�*T�o+	\�����
 I��x�]1�m&��GlQ�C�f�y:X~�/�n�W=��x�a����g~R���]�C������J��X���'��=W{�̾�p<|Jͽ�xj��-�Al��9<��dˎ��k���(��V�m�OcX���4������T��eC]�<�J�9pg:m3�2��(\!.�q�#FE+xNn-�ʪV-1�6�l9���X�6Sz�w��'l����[�>�s'n�&A�P�1�#�q�-~9�?E����H�Lv�^�f?���M}��8��b�uи�a�.vx�V`���(�bD#-�J�b�a_�����z+��x�ݎ�칚\%اsJ{WCӷV�G�u�f�i?YB��<,'�S�v�͕*��͞i���0]f��C`CE��pc>��̶��)nmh��->S�9�vU�C}�]v��:����o[u\�.累b�8�nϱ
���\Z��W%U��*/���6 �Aa�1Cx�&}�=g���XOd�:�B�ޭ��/����ni��=��bf���0���q���l�N�L�J�B���C2xN�=D��a4Qu�+sY�&P�}B\�{E����kǳї�v�q2J-�i��9���ª��8��^D�Wѡ�ǎ���K�#tt S��!&i��,���$�s�)�}��X�[�O|}~�~�ǫ\�h�la��t��]��JԄ�F �;R��qF�$�I ��f�Xsìd!f��a�ܾ�ܕ�So��M������X7�'X�.�w��xc�i��L4�e�11(���s�?o��Y�� ���k�]K���*�95����xz����%�'=s`B�u2}�|4t x��*��Є���H�2տ�TԖ
����%��'��s��M *��gi�j�,Ծn��ݦC��^ ���_sB���2�r�bm�ty�N�����cԒV=�݊�w����¯����*ww|q����%�/�d������T#7��ևؒt�3��	�a1 6�*L[�ӏ'����7"z��$A3���|n�w�ɨ�V���4_�C�ylj�-��EZ�oYBv�>⑊��n<]��w	숵�79�^^��u�R�#Uz��QT}�+N�+V�ι&���|"��R����P�|7�V�X��Ml���v4ៈ�2ib��u*b�|�4SpS!?�̓�½ⶹ��mmR�t�yY�S.���`IYWn��DP%*EQ+�v14бX&nZ�`�s�,�En�����̲����[��ȓv�N3�ɸ�����[����K�0/���N�"qS�QΌ=���<�g��}�ڽ�GF�6�l8-��VszhgHV�	��K��a��:'hO��S=�g�ֺV�-��u^��BVUx߼_'�̙�<V窎\*<�xv��k&�;|��\��A�y��!4B�`�;J�{|eg2��{7��uKܛ�5�q.;g��Y1�J,���|6v6w���w5�V�-��G����S�c%Y���sy{r�j+4�Is��1Ϸ���7�-��a
a��~zL��Y�t���M��>�S�����͑u�:�H���drRX����b�Q�ɕ|3j��LSH�
�:��I�9�M�_����� [�^S6�Ԇ��3�K+��LD��Fݫe<H�
P`D�e��u,CB�9���1�H�a������h�.��v��Lv^]]f#j	a-5t�eL�;BT�2��h�\�	ki.f�e�45��	P���͒�M��glm�@a3,��q�6�[��]5�jmUW+!�����Ѭõm�����5����1����a4�d
�"�~^F�_��+�[�'��1�yub٥ٛ:���M�<��]wnz�=�;�E���\K��&b7�μd��Ю���~a��5^K vT�Y�ŵ���Ρ1�W��){C�_G��$��˵���!�.�f��{]SJyh;��������R���ʺ��3��\�֒�F��!�/mo��%	�a�a�����*S�=s��lm0�Ya&�cj�f2K5ni3�W	���/�v��������X��T�x�:jY�s,�! %��c�Ͻ�y�ބ���w�2$���R7�٤n�^�%U컱 G���wU2�I�*ӯ&�)n����h�U�z�$=ސ@k����zǯ�J<]�E_�}rN���ʭ ����5�	���fN�&ؿ �0Z=<r����zwi1n�|�s>Z	�����w5Lъ���!L.�3���L���S^\1��W'�{�$�E4�F9��-^`v�S;Q�.I��X�M[�Tk�9]"}���&p�ź4�˶p�����X����-��X"x��!_i9��ٔ{;���t�^W�m�޿g�e��v[����ǚ}EԮ��ЌPL�ჷ)T���ʫr~�*�%���x�M�pu�k�ҥ���tt�@Km�Z�p���Un���;k���B\�L�9t!۳y{1Q�#޼��#�cͫX)��z�����ވ.D��=�޴M/:Vs.�ʪ��x~'�7x���M1�B$�@�M؀�"�f
n��V�V��"V��7j#]�o��{���|o5:��@��������Gu�ܸ ��?w���D��,���]R�;�U���ѫ�M�`��!G��u�ٶ��`��}�E���\=cI�T�
��(�j��zw�XoT�W5���>�Y��ykv+Z^^]>��Y�B)��ġ*3:yy<��m�����ٻ��)||1ϧ���_]��n��|i�Ԣ1ϖ�ݮ�S>SN�r��=g�^��W:��UO�����2B�iI1��Uʨ{�����Ȝ	J��A��r&lv}���>�o4�9�=vu�B���ok+�\�°�oӺ�-+�.?>5��oAp�V��Ҳn�2�åL�>�|�=Z1E]�C�9�x��&����Tq}f�;��;���wn�ѽ %ɏz�u�M�˥]�pD��Xc�ƫ�A�	A��1^6���	<���w"�\8I��P�q1����3��f����qk˄�,h�-6��.��f��$�}��#x�&s=�(���t���<�9ϸ��P/)��Y9����V���n�A�v�:$ 1͍�rLcG��2
�:�T�z�W^���r"���<��Ł�݄��u�;��!/�?9Y�'�.ޙ}^��"9��M؂_�p��AmmC��s]9Cl�[���VP�k�'���7eV⎷��Z	"r��]�v���Қ�K��S4J��f�O����$�TBl�*
cI�< q���\= �=
A�����V<b^�`��?�W�x��e�eC�	8�a���Q�%����;��r��*��!��Í�s���"����62!���\�k�T��*uSy��ן�'ޥ��f�N��ػ� E��dq�F��nS�/㊇({Quy�"��Ƕ^�ep�;�8��8��4n�Y���^`H�׮6\U������B��9!g�����՞�Zyr�{������i<WU~�p���J��{����E��iL���	�BP�J��=�Ӟ�t�ҫ��@��e��ò�aDxA�q�[��j�4��`s,հln]-nZ�8�~����v�:H訳���R�N>��$���
�����vy3F�B�9��ٔ�c�їu
8ǠU��[½̖�0Xm�-���^:�	�5�EL��w}ׄL�Fx:vO���f��j��;�$��OI��쫻E�H�0"�����ڪ�r��$i@b��7��¶w���wX�����A{1���$����A]"Y��W�K㘹.]	 �w������lg`5;s�vpz �7\��u�F����^R20R���i;��ܘ�,pG�ʐ��6Dֽ��}G��`��������w���W��ݛ�f�7s\�����ﳳi���Y��L�\p��">+Y����Z���@�����u��V(��.�ɼ�!��OI ��[��}~��ǲ�mʻ�Q!vS)f�&g�\�+�� �����dug�N��z>!چ}�B��Mډ���UWn��ČC�ܧ��Sw�nd�f���|�D�!=<��Ǯj���	S�7HN]7[���w�g��n2)�wqa�'���O�����>�2�eη��*[�[�'TlD�ZTʀD��]����MT�f%In�ّ[X�K]XX	A��-@��n��#����'���EZ�5j�zBT�s��O1p�GI�8�������Q<3�mZ�m�!m��Sx"@�r�9^�5��=��͹k|�ǰ�ۚ�˦��7(z��>���v����d�I�0�Y~
k��6-8n��g3<"�N!I�$t9�'��u�G,C�Y��ppr���v��J�J���uLAW���=�	��UJ7�-�Vm�wxߣ���&lv�N��XP�k���y�-�Ќ8�I�����dF����O��8<7-xB�~H1��:��
b�u��!�]�vi��2�7�w:u�H7�]f��ҝ��5�[�+Uog^��,�w�"�3_Nx$p���x���Ymb���\cU�2�P��:�u���փL!h1�EXe�g��ъ�,,���>x�x��Z4�T�S^�-!	THٶ%��t!����e�LT[k.,�ˎ&���ʫ*cZ/:�[^C�G��2͉�k�ۅi%�1ՙ5��U�	�%Ѫ�0�[u��$��Rc�c�9S	�gd��`���jl9H�����X��/V��v�
�_�>���E5��=?��o7���5OƝ��UC\Ĺ�O��]^��ҷ���	8P�p�؇���s�6�z�^����M.�n?^Y�(x�a��&�j�>
�
�0�&��ߵ,�Z>��}��b�P�ׯɋӉ��P:�rCŹc��BBdȕf���l����f|{}R�t/�>��~�|�����j7\d���4*Ǯtܕ�eb�F�P.�m���Aa�wI��ޒ�T������;=3Y~�{|����}�T����b,{�W��>����{�@��K�BWtmŷ�k3]x}�#y��zz�Ϥ�ϤACHPٸ=�p�[=��O�(���V)w�|�v���>^]�˫v�&{ލ�JL�-���'',7����}�O�'�*Ǵc�a�x���׸��1^��X~[��<�(��{&���?xT��Ӟ\��=V���ve{���З�a8A���q�Q�)]�s����p�������:��Egq��.Sa���)K�u0�r)�=q�wHt	赣�6e�795���`T"�0J,�|:���g�v�,���[��\c�����M��	㨇H��΀^''�p��o)K v���䫩�C���|�ΰF,��YCf�ƅc�g��'`�Y$L���j��S��Ss)��+-Jmt-O�$��K��u:��[��t��a��R���	|pN��#�H\Z�_]2`��ڲuΘ����ckW*��5FӗwP��EԶ��w�`���`Rx�/2��}{/-�T�\7Hi����4H��|A�:V��Ң���۶�u���/�;Ts�7�uս"��A�	RPԲ��� ���d$��$�� G|7{WY} í��Z�Hޫ�G�3���8JR9F��}P�v,���{J�Q�tX1�l�Q6H#� �f��g�S��]O(1e���+눥ԝ�7J�ٲT*�N�i��sl�jt��3v��7��c� @�ys6WKF��z�Բ��[MMV�j��9���2��1�ыg\&,��S�}�qC�T���`�����m�z����Og]�n��n
��u��_Z��d�p�*�e�&�� �{F700M�m�=��ś9D���ֳ�M�a{ίjq��/P�z]����s���c�4�\�EN�*z������
uE����9�,��܎�Zd��睐�x��t=�Vdu{ռv��m�o,��y�T��hv�w�S����åiL�UY�Z��������/1(�f�G�Y-�M��)��*�q �c�N ��g��L��M�rҶ�9%���W%z�����C�W�Y|v^3�!�n����@5rji5wI��[�M&�M�Qb�]�6��Se�UT�Rl�h	��t� eʪ�����@ڶ��T�UA�d9��&����뮭p���.�]+t��"Y���Kw��g���ib1)5V4vn�u����*JA�t�
��![X�`���܄�uY��<8����,L�1� ���7�ح�6uʒQ�u��e�A�v.�qX�K�T�f��^:�,��I�+�����t1U�R�&��(̮.��+�f�,[����ݓV]+l.�;@�����e�Kn�a���к	t&��M�2�-.i�,/#���9�m�+\��lƔYeՕb�P�B���Dչ�*SW��եɠ��˂V�$+�%,�?��^���V`DE&���Zay���F��<Yu�i���.U�a�-�բ!C 6��,4M���h#U
�Lj0K�c�m�uYaAm3l9:Ķe�k�Z;�+�3�2�vm�5m�Φ%�h��H۳�d�V[�������&�I6�\	��4)�������*LX�R���[s&�������hSWf�������j�Pe0�lz�e��4�j�9S=��T��[]a�Ж�32b%խ�٭Å���b��N@ڍp���u���T���ukK
�[3v%�B�^l�u�m3CG�`&�u�f3���T�;3U�flM�g
E�Ձ6�®yX�Ԏ�2:�ls�F9�#��P���K�굷a[��.k�� ��]�|�o�:��Yb�e�V�-��1��)��I��%������L[�F��n� �6�PX�5ATMr�`f���%��V�	K,�H-%��͕�f�g�R(M��Ypeέm�$�5���&#hb1u���jv�����R�*e�{�mT)���j[s�Q��CrƖ�j��Bh��ܒ�XÜZ���EծmLG�����:�dX�]f�M��nΫ�Mĉh�ڲ�A`��*�k6��X���
V,	4������ �.��	p��_�pJ�4�e:��r�����`]�}Wfs׳;G2f5Hh3��Rך0\	�Z��!���X���ɵY��6ٰe��m�h��CD���
)��s6�iJgS�1{5F��q<��RU���$��k*�w���W�}�V+�:D���H�Wn���}�� R��V�{u䯞�����髢�<�u|a��^���B%;
�LX��`�ūkl������>�Tb��8i�{��<n�W�g����F�%���*�D�w�a�0���{>Gps��~�>�;�����I�d�c׬�����rql�s�Q�[tyy������WMW6K|�m{�ISSש?�]C�����A��޷��r����vY�齖��Fr�+n�Ӭ��(�/m������5�����X	��H_W�����,I���ϯ4W+#~�-���sjt%Q�~=J��<1�J�ͫ�s�W�\<�fe%��'z��>�΃��+���S1ܢ�z�1w�L�S��v�?,{�fTw7Tb	��R���4��z���wv�q��#ఏ�4Vhe�i�ϟ��	���e�t-�f�Pق4��l`G��Z�(�N�4$j���3~�)Ν�y�D���{�^T}�do�a+�9�Y/�}r#�jw��j�qs�ё�c�9����A� ��~����e�i���fu�5�^X�7mA�ΩW���Ri�iJݩF�Z�;k�7r=�J_�xk����n&_4��&c�&Q^~ݣ�mx� 0�{ڝ}0+���^��:�;�f��;b�%a����@4���M7r����J�.�>�4��*M�D����\t�l{[������:��p�2<��2{<�srn�UY�_J�Fv5.1�����dc�?<�ʸ���G��X�g:�t,m����6��h�� �[d��j�xT��.��m(Y뼫�*UY~��&������=��>��;��W91��~�\0R��\��=%֔F�}�燺9���%�d���+3K�+B^2�������P݊~�4��ʰB�)xk���6vC��+�x��!z8EU��	�w1y��m妹��Q��y7������h@1|�ً�	񚬬<�x���a7�t�O?u��g�kᘺ�T5�CR���v���7.��b5!7"� CD$��>��ن�|�27?y*X���+��o$�KZ�{d��!ź�/���~N�I�
rpˢR �0�u��*ܯ�y�mԸ�%��"�޹��^|�\�}� }3���bk�-Vx�9ϻ��	�1��S>��3`��E<��Ða&!��:&�g��,�ggn�8/.��s'�N�d���]s`P2�t�N�V	i������7�5j���f]�vi
sp���/^��qw3fZ��p^�%A=�Q���U��m�5�,&�zL�R��I�C@���s����]�A2�i\CB�<�t7�7T#���r`�A2�F/(txFl�2�dx�o�nB�=�}�E��j*r״-J�j���Q�v{�.'� q����S&}��y���J/'n�s@�1��&&1nK/�׵��&���Q��.�;Q6"��O�,ڐ0��"�MjX��ޖ�s;]*����q ��14���};���y����8��1��˞ګ姺ۇ�\�(���j�' �^�'Y�avh���.ǎ�Ad�}�z0]F:1��P� J�M
t�cWf�Wul�A@���~��wF5A�i�B����]9n�)�n��j�z:^[�JN��Q���F9��]�$z�w~��:���$�	�����@�6�N�{/%��}>��'ӕa�d�v!^2��Ƈ���cD��y�QP~�ڣ5���8�\�]��vd�/3Ϥ׫ojo}�~ԗ8�-��L��q+nŁε��me�rxY��<�7�n��,��|�6r��I {��S>熈Ǫ
�^<"�,C\��v��*PI�ł��;��~pe�o��ne�^�1r��d(n}v��Q ���!S{��S��!��ka=�Lͬ�����>�ֻ�/:Z��]v oxq��"�Y
���&��6�P��^���KH��D�M�2���)�s��G>+�ChL�Z��j+hf6m�!Kf���`���g2����2�u[�Y��V�����^����v+��\�i�U%lu�;x�| ��3b�F�XbW\L�r��դP%,҉aIK�e�[�aq��
h::�t�c��!n�%�� Ͷ�����JƤ[�%�c�GUb`Xb�飝��n����6J�D��ԁ0K3+S=�n�6)�I`HK2�+u�X($^ֱ��|>>��پ���hW��4:o/`U��ծM��e��b��n�kǏ2�'��4�6׻�ozJ�^��N��*/���F,�V��^�\��Y�({+����m��Ң��Mѱ����]�;"�Y�� �������j]�Ϸ;C�i�����n�"�u�V��K���rG����&�it��>[e��jC��`�@��$�u��eԈ	8IA��-0Or���[S*<�s����n�O�XM�C�ʵ0w�J~@@�2����{ށډ��vo[���1����(l0XE�*��ss%����[x�qQ���x�ψB�8c9�vr:k���Xll������ ���2�N��z�-�u���H=�b�}�&!�M���2�<*�����nb�|{+'������\Nӝ@��ԭ�S�盽3myY@���U�#��S����8�z=Y��n�Hw7��Ȓڂa�����r�Rʼ�3�P��'霳_S��L��5��j|�{&�I�f���d��>I������*�wt��2R�Hמ��Ț�7x&�I$�4�dD�ؚw
Y�����|��Q�G{.{~y��}������`=(0	]�|��P�t�~��O.�/p�b�S�V��\
�n݊o{��ز�9����^�z�[F��V3?&�6b]��{���*���7��R��>�7s~�U ��������wj
F�-H�z�2.Tz��-�#΢�ϵe��o��O����'��d�D�Qԛ7.R�����ٛ	sBi7��7��?yO��m#]�\f�X�L�7���ܡ��5U�����%�*��ӣ��w�mvV]V��5P��m��f�~\[p�Ҽ�\Q�o�9F غ�犻���x��/C�+߳iv�V�n�e߶;>�eKW��gu\�n�ԛ�S��Y��d�3��1����Av�F�ާ����'�*��zc�y)��,Ҩzf�D�<�3+�R#���jf)tI��;�3=�飙[�w��0��oQ�WϮNe�u]v�@��@���3`�P�{�mu���Tu�����L޴=��B<����1��:ç/�<�ΛY�����r���x.U�5�+�c�߯i��[�^�^׹���x8$�n|449bf\��=Y�}5�.aU�Qx���WKK�zߟ톌f�Q�Ӝk�0T\'zs�r=x�Q��~����2s�����*N��N��xl,F�p�U��w` �����`��<�=<�-����D]�-BQW-�L�\b[[��1]b�uD���Y�Z�矡̍n�c袏9���d䭺|a�\����R�;��&��4E��\u�;��Bl�����N��C��:����e]sU���@UЇ	T�6��ă�mɝ׽�t���o6�T7J\����/O��p��L�)H!��]W��gsv�u���j�Aa���5}�ލ�*O'eق��9Dg���9t��F���َسy蜿!^f��,};�6�g�9G6�p�%�284=\�g��Ԟ��h2��vN�6^��T.��T�7�����g�o=�w��t+���K�1�Ih�,��?+>�ϥ�Hg)B{�';�L$���q����.}iXY�Ly���i��} �2����R��M��s�>��382"ho<Ax=��Z=�$v�_]�6��E�'"n�����^J������Ih�D��tJQ���jy�p�6��)+�ѕ��榇x"yF@2hd�s�0(���߽�#O��\�
`�)�[����S;�;J�Q��H�`��b����P��n�k,�y�0k��թ��
[������_�_R�z�s�[k`:1,�Sk�	T�;c�� ��(l��a0���6Fg�ua)�˿y��{��fb��sR]�.f�g;�%����x��cuO��g���FS+;���D���֙I8-��i���\u�DFks�����r��;�:ws*�)�1�d���;A��1� .�R,C1Nz�'}�s �͜>o��U��=��6�`�	m���6�����\#�V����q2�{��OJ�	P�ǂ�Ӯ����̺ʅ�;���f��e�[���dE����qg����m���2j`��~:�/;9I!�=
U�7\����{#�H=J�,>��	w������#�+�]^��3466<}�ю�Q~�C�1�����٫�D@�V!���_w������2�A��*���VfL!���{��bf��ݣs���\�Pn���1��?q�ACYM�%4�o��Qϭ�Ț2;���O���[����as�7���ozbx_���9fV��U�������93����	���������cQ>
S��[�C����!�o^^���ɠ�jF��b	�B︻��<�'�l�.2��y��R�{$ݥ�7CA3\]��ι�ZV:�S1�C8%n��N��{X?=q��j��q�I ����y�ͮ��k��=-�o;���ק�F�J@���]u�D_�����G�ܛ=�Xҙ�`	��/��*�;�yx�*ѵO�t��U#�W��b}��S[����`����z�֖GA�O��WDN�7�<+�ANб�L����͐����L1�9m�%g./{ޛb�8�?s�H'�<���e{۩��n5!�A����KJ�{�4�	6_��.5�� Z�R��V��]��(�T��k�/��n򙇂m�^�����ھM�+�Up}���V���][��� ̎�6N�߭����َ�D�n��β�`ݱYF:2�8Օ�Gh�ˆ2�`�L�7�$�̀Ռx�[�q5�ʎ�Ѯa����f��Z��D��a@�C�bf�u�G�KeS���b�)��p�)p�;mf��0	�6�FT"�d�Z!�M�ƪ!^]�Xh���ib�,c5�F��A�F)V7b��3d�v@�X[W �V�[�ZIF�Z�Av����p��Lg䲹�@��pn^�3���B�,�k��h>�u^��Sdj^T����ٳ�mR����A`�q�8�:����O��޶����}\���b勒�5rrd����vB��ܜd��B�MA-�b���V{�+�"[�8c����%/�g/+��1���>k�5��"�B�2�@AR�7;Dv&�^b6�ju�ct��-`�9��N΃H�m2�����G�=�$�y��q~]��z�*(z����F�#�c�j��2�q����0L"ݶsN={1P;��W��V��v����5x���+օ�(i;4z[M;��[ۧ=󔟐*����ۖ��n�Ľ���̗������d�6Ue���5�L�1���^Ϗ�� 0��UɃ&��s�S+1\�ꆧ���L���lQ��6O�z]>�9��8�[�I�M�1=��=+�H�t�~��|jՠn�'LА���T�h�n��F˭��%;~�봕JՇ���ǣ���R�>G�'���Q^:����[���ټ��zo������&�Jm2E��3���JC=��w���r��/N����AkY��F��e,T�>ּfs}H��a��]��o��;�G��E0N5��kYpsf����n�7rR��=�"��m�����l�G���ǉ��lF��0��[��_��}k��QC�
ӂDk�3T�g��>!�
̨־0x�e��7~L����+Mm�U�G�i#���0�#n�-(6�.��v���Y��؎����5ݲ�;"�⽛�sv=�g,'<g��o�Gq��:�^ڮ���q�d���j`��y�����W`?�Cu��HީΥrӇ��uS�@>K��>�ِ&d���I^�hkq���V���s���p�b��5��U��	~ŔcF��%�q�{��A*AiX@��YG(�,5ҥ��I��Uȋ�(KHg�ܟz��b��1�u<@�4mޕ2�TJ:b�T9�k�"��<�1Z�dH��Ì�ܺY�Fw����BnL�uhq�J�O�K�U�;Ƽ�B���J�W�rߟsr����|�l#{��;�ݮ��s\<$C5�Z}|2� T���J���3��Q.�dyjD�H2�AgH%]S'c�v��Y��߆����φ|;X�/�F�|W_%�W1�j'R\���u�K9�Mͩ��^8|䔼��t������*�bΑ����vn�Q�v�AXA!�7#FĖ����Z���ʯ���x�s�ם�9�H!�6��pu�56 jR�m�k �����d��%�;�����C\�y��Z
<+=I�FW_��ܳ[�!b<�B�ѓ�(�x^`zF�Wn�!Oe]��؈��;�+}�B	����O66�'��f#(��y���6�w��6��i�WN�D��yuｘ(_`���d2���$TgL�gwN��d��J���PB��y����3��!�D�[�x�_�WnO�v�V4$e�%:�S��mr�9�^S���M2�$�,s���g]����E9�:�O}6�ώ�r��]���!�sx���b�= xz�۞���Ϗ[����QW�u2���E��Ӟ�^�+C�&�>�=�Y?�o��>'`C��74&=u�+�a�oƞi�:�o�ض���zUכfvv���J`\��F��:�c���˯��4��׃��gt!&�������Vi;�5"�_-ݫ��/�+e���'�o�l�י�h"���Vnt|�Mw9^_�I�h~� ����3�.�e�V�a=�>�]���c�x�T"!�ĝ��B�>ə���$^����:ݱR�G<21�7��\�.K��M���)w_%��l��(u��HUm�&."Qj��qwoM���U�jJ)	�}��|���"c�5$�V�M��Qc��R��}t~�*>x�?'�M��$�D�2�E�Iw z�h���S��h�F��2{��M��
K .a?K�/�Ș2�MO�z��X~x��n���xw����SyL�x�����	J��V�����x���%�)GGg�V|��ɐ�b�l}�(٣[.�׊�=��!um��;��9:'��Ʌu�gq��z�]W`CO����}Wn��Gz�j�[t݉j3|��ӽO��:��W�6ky�3]���8������mɏ�Ηs�к�����Wu� 
wҞ,��J��Gm^�������������Yx�[|ӝ����j�V��V�F�)\�Dn�Fb}v�#��ڷz�N��{�rux�ǖ��\�Y'�u&�fdh��Vu譕��2�.�w����X?bGm7%�H�>��CZ2u�����+x<V��{;�Mfs32��/���ݲ�
'na�Y�u��fcr��/��t��ӯ��t�쾩�:��:�`��賂ď兙x�2I�v�bμW�:�
���[.���#�Ju�ǈ]�c�W3���zR2�ͼ��A��g��St���=2܋����M����V2k��7�v��ռ���N�B����ݨ?'OCAȥ4)�&��s�rTL��yCN6���r�;�[���*tI}�=���JwRZ�-�й���57W���r���]����1ÒY@�ɘ�	��sh�|��Z<���wfr��N��gWu��W"��S�Ӈ�fh���lt���i_M�aM�����Y{g�n�}sodo��xC�������X�.���g<�ȗd#9x��,��s9�˳�Ğ��poNdV�gc���	�ڎ>�+��빃��Gu��	�DؒJ�������������.���\�����q��S�.Ͼ�y�ٱ��D�a�я�X�����&�������|���8� A��b�BK�W��7��u!z�k+�t3"��o;I�!���0mz�Zٌ���N�\&�����p�rw�n���4��d��y��;Z��y�����d�2.��v}�w��@���������&�.}2:f��N;��oi�{zlnz�<<6�~�;���꘸���2�E������Î�7��؛�E�}������n�IF�C�bHI!���kM�fL��2`�[�����" �$�ȓ�~���z�0#;W�N{�,Qj�:�{��%��Lw�J�W	
a����F��[U��{�ZAH3	(,�ip�h�۪˳�W�wE?cW����[$t��x��H����4��uF�-
/�>��>⽍�LsG��;9��v|���~���DD�����U!Me��hd�
�_{\�{�D�]�f�����L��[]���3�l^4�u�Jy�X��Vl3c��d��;9~��f�� ��Ca�Fڙ��y��~��"�m_n�<^U���IA��z��'����i��e,�)��y��F�1�V�|��d��K����5&���e�U}8�<�ߞ�O�=��Gޞw�l*�� ��"�X�I��J�W]4MWFծ!B5�6����j8�@���\�5�fm(3����.8T M��ݫ*\Yi�pv��ka���4��&B��))�Z�f���ù�p�a�6�0ץ�;���X�Ge�R���b$�@�ˈ�֡4ID.�u��lF��R�20nqKM�#��#Y��V��Vյt�&B�8P� ۾��"��"�`�I��m�o�������΃������0S���a�Uu�d��,��V�}t�S�����zoDÐ��|�3�Ur�,�P��S/���Q��I{׸#!����R�����pg�1�LL��4�m�;�͕���cq�aV}�>��}�����Ľue�@�2�Hb��:0�j�-0�	4�(3��3ZW�ܜ�8���<y�7���,�D����޷C�c���f�|�czr�[v--gbL9#")8$_˔Nw�_���t^�o�r�(V������PԲCE]<(�
ߟ�o!u�e�l�绛�Uc9D���p�ϖ�kskf��(eS�'3��[�_f!���U�c߹�����1���lw���Q�#�s�/[���n}ơ�������t��Si�x}F�T��Jʰ1�7ɇ�8��j}P'#����v��w�||��G��1��oޕ���|m��]Ll�dʘ���g&�vg�~�'���j	��?	g{�:]j��g�T�g���O�N��;ug������NoL���>}�=��pb�����繆����/%��v���>��]-t�/5��pqŷ��Β�����2˻m��}P#�Wc����]䕎�p����*��9+��n���w6�'
':9�S�:f��_�\�����w&oд̞�0���p��P��Il��f殽�Qk�J�3sq5#]k/\��������r��gB�� Ƌ���K��S�jtv��O�@�KM��Ζ�u��d�XN K�r$$&vG=�_�n2�W�����3۴�gIpK5��H��-�T�,�+(}�j�����>k���f��%�z��^��K���H�ỵ�q��{[�����6�c���E	�\1~���ѓ�+oK��r�lq��_W�%�F}�"my�eu� \�q��~�����%�p���Q�����B�T,:������C����af���5����1�k,Ь2��+�q8�v�<c��iw�ﯾ���7 �VwKǐ����V��)=����d'���o|�R�]c��~���#��ɣ��ٵ�[�Yh׽U��(	���)������B{�5�\��H#\2D�[���ߢ��p"��~�m�&��/ď[�#N\��1+�ō�*v���9a4n�[]-V7��3��!�[�@�����}�Nq�{�s6�喸��<j=��;�=@�q����y�m�X)�0_��H�mI���k�T�
��ao/-=�`u]�&=�bN�Je�g5e���h����K=]/�*4.��ۧa.*b�{�X�����O�>�8�m��������P�J*l��qį��=���s\����G83U�r ������i�����Vd���� .^�S�*���~E>��=���"i���ʹg��1ӑx�W����&𨪸��
S=�F�q��G��>�;�g���f5S&�z��Uo����w��/��_���QBs[9�VV5(q��{�9�����Gך���_�����=�h����LBh��i�*�l6��nt�;/�����#��v�0�Ǆ���75���F�f*���pm��ہH��z�슣�1�ힺ,�{�6�+�H�I�R��ù>�?.�<��U��<-�澃��m$ !�!�[���Q)4���� �]��5&4�m�Z�?����7�~��M���Md��1�Qy*)���OE%�ym/�=U|I	}��g����T�J���-�����K��C�O؅e/vnM���>"�V��L��>}��C֯LHs���:�q��*#�X����`;��N��`Q��an+�.k+����>�B�R��?��`��G���f�4ԡCdC��MӇ�t�����z�~���ٌ�D�L�J߭�V~9��Rek��ڱ;7r���J�؄��#x=k������i^��=�sm9O���fg�ِ���f2���ݠ�:����)�n���R�{ƃ�f�+K���B&{3�Ю[|_�#��l�����%�����Shժ��R�=~.n}	w�éݱ��N�k��ep�|�=�y@L�I��u᾿�G�ޑG���"�9}v���NQ�N�2+:B�.�9>˫Wz��u�Y��^�O���]�Y���+����8(n)&A�7�NVVX�v_l�^<�����Wu�YLq�R� �-�c��%��m�6I����p�D���(�!J0�vug�z�՜yQZg3�g�.;�p�U�5kB�q=ޘ���J�����&����ACA�Ubw3�p�^������z����f.��������ht �MEzT�w)�@l���p�9�V2m`������_;�ނ���(�IT�<�$y��]+��ky���U�#��8`oZ���U�Ѵ���}~�yR`�+��Ń�f�	=R���:�E�̊�1�#0�יXV�w.ij�W|�2�����}���n&�NR�T�	1Rue(->V�l�,a�qu�rs^"��p��t��uq�x�d�Ӛ��s���x͓�>ArT������)l�i�R�e�`���e��X3X�L(�-��Թ�X@���x�Ǌ�����֠�,ة���5��4d#v��6�𭺪��u쁪C	.�	���\V��P&�S�@] qԱ��ɷ@`� .�B��5��v��0���[P���b\1أ�J��H��Ɔ �Zokq.F�ؙ-ؙ��J]��H��l�!�C�#�Q}]����x�`�Fd��o{v���r���;���LĖ҂��T���U�9�m�߫�h1�4�"u�,���V}}}YPO��94���Dw�nE{����[�%�S=�?^d늗�ㅚ��]/:%-��>?#�;̙J�!�ɗ��ެ����޾���ءKIj"��j�Aa5��4���ա��:�ܒ�k}���_�>���=Fɮ���L\�>�c��~Y�'Ҿ�kEpb�ݜ��??f.O|ǶzU�9��B�/{�9�d樼;���nC�?`�Y4Ѝ�}�c�;M z��	�/Jl��n-��Z��g5ۤQ���?�Z����_���f�� ���*n�����Ē�d�L�z���e�c�f��W�U�vX��Ѹw�����XM37����������O����^s�B��R
C�7ӎAŕ�����v|��"PY�@7��⿯��
b,(�B��v���veg>��@��^�$8��e_��_H��I���S���iN�}S�d}�0���W��a��~�1��QȾ� "F�	p��DG�~;�U�/��R���-� ~��>����2���D G����f<w{k�+%��?_�<5ϯ7�l�.�n�-�WSh���4��e��m��c9������Y�/n�ܤ�l�}OCn�5Q:��}�Ǹ�/:`�p�y�b��Z �~���>�=��p#���xv���ҌE߾$m�Dt�� M�J��Q��#Oc�=^;�x2E��ؙ���)V匭4t�����ڇ�Ѓ����Cp�`�!�e�mW�`�'�x~\͜>�c	���Ᏺڏj��1#叧�xZ�"���5߂Qj��~��}����/�x|Fl���R0c�>�8lс���<~�����ǁ
X����>C�b뻻�h�Y���<#Q�;��O�ˬ��+�\̜?a�ç�s�}^����!�����}x�oz~z�z|v~Jd�� �Q��u`�������[��j�ڭ�\@+�=#���'W�� v���L��`��Y�"DE���>9��>�?>U՞wH�՛�9���}�Sy>~DV!^���E�ì�m0K���#���C��>�7���F�f�?X��!��,}��g�x}"=QZ3a�^Ё�?B:~�廡�,��|=�z2 i��E���2=a���8h����V���p+�%��Q����M>+��/�7<�؊C���}��s
L}�<2>��oOт�;�w�F��_�`����(��� ��y	 a z��������]uU1_�gߦ[�X2(�߼�@x������c�g>�0�#g=�ĂF���݃��(��4Gj����	�?�6@�!�����- �+˞2��C"�@�-�����`ķe��,b��k\�΂�j�Ke�+��_�����O�@���mD�@�c�G�mKp�+�Z�E����GEVԑ�(_������ҡ��GE^�6�eh��m�_�|��CJ�V9�t�F�P�)v���8����;��ܵQ���n�M3�������K��FQa�J	�_p������8Q��?WyU$���xF��L�>�?Ftל�$�0�O�~�H��Dq H��y��
�W���gf�B���7����-��q�1�n�o8@��#�g��G�u��	�>���-6�d?f@��>�� B����뭌�ĵB`����8�E�4�پ��\}�CC���x���$�3���Z���r�#�#�!�<EE��|��>[\J���o
?�����_x�uݮ"�#�歉	#I����w_��d��c�g>�<�R+�D(�,�-��A����H���Y�:���G��u}Ix�95F�^��G�W鏰|�G��(V���l�G�"#��gQ�� G�1�>雩��;{�i�`F�(.D 9�𑼛��#Oç�Dfz}��/��8���V���vЅ+�{�{̮�?a��GH��?���o;y�����a��Kw_�1���g�O{�����#����@9��u]�Ç�7�g���FX3�N N$<P?�~"�9��������BDu�=w�^�ϲ7Q
 0n�JBl��Qj:�X�m����Jaq
VV�F��"�/��׾���}�?>���`ik�X���������6>��;?}ؾG�g���7����Y
:�h��/�P��u��n����H�����K~0�e$�jX��־ҍ��@�^m}˻hDB�~�� }�H�S̟�O���|<a�2(��涆+�K�|U�� ��:���u
#O�!��'6{�r!�_{W׶��6>dD��r��HY��s����0@��������M�?���,~c���g��~��m�Q��kۥ�IN���v��ˬ}:B�w;���)��(O��c詒��w�μ��-[�;���I�xXI��u�0�ȷ^nc�q�	��Io�;��? � ������6�~�>�(�1L!y|4�8I�;�|꽅DGI������i���������g��s,t��(���B�;VG<~���>JC�@ٯ�@���G�?QGܮ�dU��@g���݌f�(�oHq|u=��>���\���$t���s�3����#����`�mlO���0�}���9i<x~Ҹ�?|̺���xE�I,H#l�E��/;���A���ݽ��1���ާ�c�:X|D���F��g�&�]�z(�,��dYO���O�r�Ae?Y��@�ݯq��_���~�|˯�"�� <Qg�|	�|���p���c|�0��"2����t������Ѽ��B<��$�P��"��Y�32 [��0P�?��!eWFK�jಹ�a�n$��8�qDr3���~9��Ϫ�H�G�Φ&"�XC�1���#�M�X�c�,��Gó��ʗ��_ v�?�?���a z�*i}B�U{Ղ=���#4j����"䐮|H&��\�"O�"4}�3g����>��t��>��+����P���t5_
�����xx�=�����>y�pp�m!� ��ؾ�󁟺G��#�����X�/���������l(!i@�>��kWĉI��}�0���⿾����e������3�O_]�鼝=I�%%;��$�đ 1:y��B �,�A?}�9W�>}�{>��ͫ� z���?z�w�
6@w��UYwβ9�z;�(��M�Ą@D}����G���x�=W��O��4~�8~�Q��׵��-}�^v�ToO��-0�w`T�R��n����<�S2��]	�{��7n�+��&�+�كj�ME3t��!�B��uG'�t���Ϟ��}��T�:Ԕ2Q[�z��׆�@�3B"Rk��ue�/b]xI�H��jmt
�dJ�L�5E��c)���-�أ�ɺy<��Y�%�q����Ɖ+�q)Hm3�kZ�V����T+�و&I\���M�J����ŭB6Pn�`Q4̤��e,�atd^��j�=lfv�� k�$���ۣ@k^Ɗl����(��D P�u��}�Tp��d��s��!���>?H��?`����?GmN��}���c�QR�|"C�~�r�πD!����4�dl�1�H�.lߕ9٭z}���}0vb`s��gw�7� �}d|ϛ��}��>����>��� d3� G�F�������#�ھ��$�~�9���S׼�2��t�����!=�ɡ�G� ����?p����H��jş��{��R�[��<#�+��+\9Q�(2H�!N3�D�\V�DF�1�Ɇ�i��jvΪ�)q��ga�'��Ϗ��}���!~���� 2<~D JKn��@��f|�����l ;�_�W>���H'I .;�>F���k�N����p9��4k��8.�i��(�A?Y҈�p��J7*�أ��"�d+�g���;�e'T@�G�ud{|��朲�}W���d�� gW�d�p�}����#����~��Q>�f$E���{�X�nx{S��74 a�(�0��;�|�ն��y��3'�>#gW���M@B>����}R��� `��>�f�o���}0"���$���̟�G�܊���S�>�͹#�B=�ϙ���D̂H`q*�	))��̎��D�wϊ�A����T^!�zQ+�b�ʏ�>�!ި��!n�0H#���ŷV~��6���h�������S�r�8tGՍ���jb�|�ar~_X��]�w�����*6��*�r4]U��*����o��	c�u|�Y4����Ç;��1�Hyt�y�}�}̾p��(���ᝢ�a�������9|�R��{l�P�9{J	Y|9����+�j�'od���ִ<4�͸����I��z�c��aW���X��r�cV\�m=cDX��P��[S��i��:����u�C�zev>������U�u�W8i˱%���WN�<��|����3�z�R!\�4�����"�
\��()���چ��.����l3-B�,Ȕ�����/K��عW�
�НF��Y2��Q�����1�����)]Aܙ6Z;/9;��ɜ#���E��Ya�a8J�}}����q[*�j���(���������-lk����HM��8^�gB�a����U&H0��Q����5 ��G+*6o+���QK��_��m�����]�e�/�|88q5������7m���)*��ܓ�L&�-f˸����U�_�9���jb*
,�H^�o�8Ib��Y�}��=%�e4�b��]G/Q�є�Jc���NV�ۻF��Xֿ!\������s6��
�f˼D>]dY����Q��u��B���n�gLe�F��n�P��찄�o�껜�]jr���F޷\[Dӎ.\�f�=�(�0�W�xR���nWwr�-�h��d���E�+��Lޫ��hU�*DK�b���X�dl�q�m���J�*���*\�Js�\f7n�
��j��Ԁۘ��uc�-���:����O�p|/V��"�iet�o���� I�2���Z�*�*��UUP�+��
�uʨgl��mc���j��۲d2cSQa��A�l�[#����i��ZV���shRҹ	��5��s�AIuHRmlf1q�oZ$a�X�i��){cbd��I��E�2�r��.c���o7`���y�,3�2n��D�Ҕ�k��\�Y��v�[fA�K(VE�e�cY�9�1B���є���	��H�6����s���yo4m]4kf"�8��м�����Ki��)��n��@����� $u��Ύ�m+GX�z�Q��"��q7!�Y6�m�Mpmk֑����b�B�8@�]��jR�K@R�	��5ΐ��CRH�v�#��!.���[J��6:$��
�#f��fւ0�Ke\�Cfh���.:��Y�R��em5�5�����F���f�r"�cE�X�ԩ��+J��%���h���e������0ѹ��0��v��֥�4�GeȫCce@����n�(��Wa[dc����M����8�6n����лM����`ȕ��њ7eJݒ�ER0�ƂSf�k�L�p�,�F9F%�])��mĚˉki
e�
P�YS�;X�k�rB�et��v�D�d�m�Bj���edHZB���I��Q���$^�qqebL\1�Tк maSa�hi� �Z��u����T�P]���,i5��-Ф�lI�,�[wT�A&��*ʹ�ҩ��p�*Rk�cfm0�ڢ˒����s�r�i�j%�6�4j��4��%��fʌiai��QhXݰ�챖��V�]���c+�ˮȗ��m��K�PK�;D�:'[��fR��p��jC,m��8���dv�.��`�)rb^]6����E�ka�6F�C@ 2QZ��hB[xګ����SP�e7i�Į���Zd��]�Y�t���T���
/R�n	����F��ٜ�[����7qR-��6��� a�Jmd�31�Pq�s��"�����=Y>����S���8���#F���=��|���O8��썇�A��>��Q)�q���ݜ�Q�����d�����-�=�v��
-��l���%��%ֻ�Wm&�,ke#Q��,��Q��+��i
ye��>�������!Z�O;a�	 ��(q��}F�~�o���P��Vop���n���_��2c�F+}�P��$Q�p> �v�Y��)�ܧ�KY`�8`��HP�?1&f�&�1�鴈���d�7�o��7�6U�N�������[P|<z@~�祖���e�>�����<>R5��AS[t>�����=[~����f�_����[�}�������ÁV`�����S��#�#��hy%&"�O�|	�ďrQ�ŀ>��t��unY�h��5G�«���^�i������ܙà���0T�$��G��$
$Ϗϋ���P�l(~@�{5�U�;�� "76A>Y�u����$Q�3��=��fu}�'���q]G�#G�8P�Z����2�������C%@�Q������_�R����!�~�f|!� ����#�؀�nO\��!�E�_D�]}���3G��Wz>Csn�ꪨ"���X"A&�hY<��d���~��	"�ԓ�e�k��G6+2��}@���Lcg����F��&ڜ�!1s��nX6����&�����Qs����a��p؄B;w�u��}��N^��!��*wf8S������=n��o �L*Ao�l@W�$��g�[Tgav���Z������7����(�|�>-��X��v3N�l۬�`ܕ���=�2# ���3�S�;�ys$���Rd��j
ȐDSZ�b(pG�Y�.g'�#���!�����FU3���"\��9�g؏���Ueg��Q;�#�����4*�;�������>H�D�}���d�>�DH8K$��� [։��띿d�UՌy���H��s0~����@�'ӛc�{���؎G�
WaHLp�@�b>\�ؕv�b��D��g����?�躟q�Wv��?�ڣ���n�&�$E���ۿ�?B|�ɝ�8�������U�PFcu�pZ�4ۼ�8D=$/��N���þ���$�l���z�s���6�w:���p�I���H}�fdU�����y	�.���{�n�:߯��z_ك�|�管��8D�ܜHbDL�o���%9�L��<��������R�J�eEb�\�8}b<-:������Q2"$��M������>~�z�&����!_�30k�i�1)[[�+]���\�ڭv��?�|D�"30Rj��TT\����'������cÑ�0H�$$�v�r��@DSYzD�Iͧ�k�AX�CR�a1�U5��y%K�^���s�Q#6T(DYf6�<EX_AІ�i�/�BY�Gs�n��w=�ji����V�]=g����7�ށ�O!Yƈ>�@}>{u���omP@Q�<p(��;���z[��Q�' �B�i�wu����,}�=	˻ֳ�ﵾWQ��=lKP'����)�NtӃ&��Ƴ�]o,�r���?nSwf��{�g=�K��$������|�w��+��ج����t��Ϥ�ud��x��Ϩ��0!�_yM��[ٜ�.�P�"z'�?0�nnj	�)�t���/�v���mz���\Q�;{߱�2�b��U�]`!I���oϹ��	�����Ǵ-w^ҳ,�.h�e��$@�r�G�Ʌ���_�b=���S����f��&]*<n��m݄�X�""��kذ�|Le��ȩ�UD�8J]��_N>��Ctfr�6!��L�	���S�EAU�<k��)��5k��}-��F�+53jj�Q� �e�`ۥ"	�wm�V��&)b��5�"̌�Ii���ވQ��^?\��[��E�6Wң�hn��Xtp�	#)U5Χ�V߽\yv�b7�8�B	���$I'D>>�͛��aI��K[�z�S�(/���:��3=����m���Uo{Ie���dø�I����%�`pz1d{��g_��:�Q�#(��/;�'LvZT��G�[ڈ��D�/���������=�C�}�
d��!$a�δ���}��9��k�5���~�z*̋1��dKsi���0
"�n�$O*��n���1&�8�c�=T��]F-�A7�b�\W=��}Վ�e]C����b�R��:S����Ә��b����e��Y�=!��Ŕ�'�38;�%d�I$�����2�vك��5�bX�Z�)V��u(QX�ۚ]w8i�gd�G8tҢ[�(�-����)���m"a�Yu,�]��C�D#[��4,vš�XM��I�n#`��՚Kc&�t5����fc6��L��lWq�+�v��86���n�j�q��&� L�q�f�X��DJ�:� ˙�&� �#� ���6�� F��LmT����Q�?
���p�Bp�jq���|M�d4pkI$��9(x�r����׶��UA<A���O�V9i�2G}lj_?��m8��z��p���[��a���j��_x
��$B���껞{s�yP�i��4<Bh�(<���nD�/�c��u𮕽Y�X�C�U�ءi��N�e�"4M���2���i���u�	5�Ä�9�$�!�Y������!c�TB���{��Thv>������\9QJ���ʳ���o�mLy�~��PDSk�bg��K&�ɖ$tmO=�'�C��T�E�V�82���f�4����8�I�%�]�����s��߽[�lB�x{4��(g�J��.�����.]Ѧ<e�1v�z����f"pî�fa\���Ds����9��LWҁ4����-?�S���W�Uw�!���q��PrU^S��|�"�(�NRg7Z�I�����?��]�J�#�q�k\�^{권q�F�?�k���~"*��)�{��kLC������Xy����MQ�"-v�}�.��*�>�{���
���\���<1N{�B�pε#�y�
{nH�Y���zΦ�E̻��;s?	���:>�$e��2�:j��v�nj��,��W�-�6VX}�Ve*vZ���i���N}���o�I��E>�>�'�g�<"{ܧ�L�S�2v�l���!�Q��^�T�z['K��/R2s����B�A�:�.6�9�6��c0�Y�M�Bf:]
^�čҥH@(.#9��x�Q�����l��<��f���s���k$>ݥ�s���`�;���uA��G�o�!��%(��e_8�A�ft,�_�7'�9h���u�cp��+|{�X�׀�+�8@��Җ���9�.C|��K7�h����w�ǟAA��P�q^�t	6O���xB�u�]�5#@F�$ֈ��3��;9�� X�H�����w�g6K�g���>JhM�k#;W�Po��G���3t{�ůD%�H�m�!42���T�ϙa�|v�w�0>�����u\��Mw����4�����s/j��KQVa]OW;�T��{���Ya8e���Y����ח�Em{f	�s�H�b7�~�V�m@i4|e ��j��>1��"/UE���4�rSB����Wؚ�o��]�#f
D6�A���ˉ'�Y,P�,���ږ�ug:9'$*�n�bY�W��#b`�]CF�
�n�&��u�wo>� o;��*�>~�ю#�M9��%D\�;�6���p�	�>6��׽�cKC����.��x�~�x:�7��w�f���YϺ�du0�r���H�z�Z�-�2�1�}�F�D����C���[$re��s{�a�l^�$�6R�Fј)x��we)���>�D}կ_�Lb$0�X\~�5#yA�<x$�^E_d�"G��NeÀ(�,r<����Q{���|�&1��٠�	"wA�[��Q���ߺ�v��"G�L� re�g�ھ�~"���츖=3�հ,��;������Ɉ�i{E�[?
���v��ť�،��<�}���;;�RfJ�*��r�ƚ�o�|����>��� ���~#=x��)�\sIg<�Lw.�W0����Z1Xaoe�����-�`�P�hm��wc�>ٶ���_�?6��s�>\����M��F�i}G�f�$�*a*K
r����٬A�8��ʖP�TyJ�)��9�n��Dϊ��U�.���������u��6 z���lR7F�8���4�1�]�2űZ9�(e��M6�l�6���u�5�G��"�|vL]1y{]�q�La�#�EI��ɸR[��g�3>G�y2[۬�g��h�C���w��������sf%�݃�Y��x람w1�i�b1��O��ӛ�K���}�������ͮM�8�L��j���Y��aBH�Z�(6��	���Q3w�`ʢ�צ��������0��o�gR|��h�z��"���Aݔp�«[{�m���m��zR����NCtp��[N�ğd���,�q�5cn�@dw�R�$�:C��ސP��ix��}�`@;7���ͼj����I�|8� -��(o�x�
/��5o#��V��t�"��p����Uϝ�9���[�:�Ϯ}���Q���O�X�}�k3r�o������nq���J�a�w^�� �@[�Vr�mg+cb�uRuM�����dVJ������h|�ó����ˉL;Z�Ջ=q~�TH4P��ߜ����Qzc�5\�Y���Nz�q�Lq$�?VG�CJ���j�X7�c砺X�y%*�Q�<⣄�"٩4�˞i0�9`;[M�ijS���i,kF>�3��Hnf���,��ޜc��|̶����1��bnWQ#r/�*�^U�5���w��2d�j�L(�8a$�A?X�z|+Ӟ~�_0E�����w�	���@t�`��`Cئ��W�zpu��ȕ��o[����_K�9 ��"���9������Cʂ�)Z%Q�lcހ��/�|Vq��TY���o6q���'R�1�׏�@���no�j�X7#!l�?�n����93�T� � _�;�Nv�T-��mA@���.H$��'�iD��5E-QԮ�7\<<V�e���ӦA��:?��nv�`��w.���9��B�����������y1��6�w$۲�Q�
י��>��ڱX������f@��䨪]�©qfSQ�,��Z#K�hGT�P�\Tq2KZ6��z�l�˝��M�����p9"[f!��bB7���R��5��Wh�p6���-�s-��0ԶB3#3b��ZY&F�`����bV[l�MIX��8�WP`R����K��%�76�c�Y[fˎfeC�.sX�,Қ�XP�ȑ�ߋ	V���d�v9�"=�� �j^5=LG_dP�?Mâ����Gt�`������b�f��c��~Έ�o��u�T^�͊��'���>���Y-e���K>[����%� X`��b��y'�p�`�
��X2�)�e��G�^�:��ug�]�������noY��VT+v%)�ڭaB��1a�01���(!E�w���F� ��c\��^F�4�g����k})h��#�eQ�u�שW��F�	��ӆ��g�|rn�E����CZ�,mOT �*��������JԹ�gĊ�������5E��S����q���j����H��'FP�_Q�lQ��~{�
�ﵓ��f2�VUw����
��pkV��W.,Dr0(��.^k�T��;z��D��n��+�jB`"�)��C�/��9߂Q�{ػ�U�~�D��黯Rq;%�'�ǭ�ӿv�����F�1��uD�bLv��Y���Wy��iϢ��tf������i���A�rP;�scW�dv]����n��zV�F�T�����Ig*�ŔM����v�
�3�i�W4
�b䏨�M:7��*:d�r�os�Y}��ZF]e������TE����tna\�#�G�{�Q��ׄm�{�P����Ĵ�
�F|����_'{1��W�!�bG=�j�T�'�B]r���0Hl�X�n�gq-�!H�M����WR��\ɯ�x���O,����.%�Kg{��7u�/��u��-������j�r��ɣm���&��	$�A�&Y������_d��vE ='��U��}<,��n�����Y��CJ�:�|M�½��3ܾ����8��Z8^�d��ބM$a�!Ի7_�fI���7ۥ5����x`]� ��o��+�+����%:�{k�Kʽ}R�x��&<k�5v��r��gLe淋�מ�'�$A'���y���n��]�َ�;��?7��[�����QaϷ�ǳ0��.���<�峾�^�]��c4tL0����m�Ay�g8$KU���s/�ط܍� ��c
ޚ�u�p��úo�v@��dß yǥZ���M���wJ������8d��JBd�3��~G�
���c����>�F� �H?��6�4�	sL�6�l,���ZVm��eiwP�f0�HB��9���]����u+T�e�O{�^5x�o��U��+i�R������"�՞�Y�u.��+7�>���՝�PU0��3��V�nN���=DًK{v�Y�Ol]��(ں��c`�Y��)h��y���wNR��y�U���]u�����xni�U��`�6�E��cy<��G�о��;�l���.��I�G À�71���1������8�Ϯ���΀�֡Y�u[�.V��k�6�%�Gn����������2�b���������%��3r�����}�U��~�]Z��|2�
�+�OK�݂���-ޖr��qGkH�}Q��E5S�&kk\ě���0�-��,7�2�gq�#�V!Y�0�����=*c��=y��$��[�b�p��+��ή�����x}��ze�ʗ;�ގ�+�,�e�	W�~�jj�Λ[���3�M,���
�	?���-Ձ�i2���3l.�b�Z�-5]ΪA}�����4�A
;c��w:tY�7����>;�$�
ɋ��G�;����ʍ�)/�:����
�� 8O{���ޙ�����1o�%;#x��)�{=z]�s��2�Gz�h�N�	7v]аY����zy�����_�I�wwwt��ߗ�t��ӻ�?����I��?��|��wwN�����xzO$�N��	;��;��,gwwt�=�!����H�N�޻�Y��9���;W����I�?�N�:N��ӧww�_���ߟ���N���;��N��_�������������/o�����3�~����?�>;��Y�����;����~���|:wN����g�C�wwI���)ޟ��쐞�������?����ޝ��'ww�~���ϯ�4���?�zO��^��?�>�����㻧t��ӺN�N�N���:t�I?Lw�>Ϯ�wwI��|g�G�w������|}\�w���������wwt������?���?��ۧ���S����������K�N���;����I��>���>�ߌ�I:ww}�;��N����M>�t���Ϝz}!��I:wwy!���O"D����|g���3�e�2y%����wwo~���>s���N��z�����i5�?�O�|!?|��������N����������gwwt�����w�|���}��?h��C?(G����������ߢx������ã�������Ct�����?K�8+�#��=���wt����z�����N��ӻ����O�?'���
�2���o��������9 ��>�v���h.��::b����Sۥw���l���شwpWj;��uw��[ޞ�R��������݇���s`�ݴ�;�r�̱E^�{���]�s7a-��v;4��o< �)�^n������ӭ����mv�[�{o{�ֹD��!͗�����u��޻vm.��t������m�=�j��ٳmţ��ەv���J��%h��ڢ�v�U���)K6��t���q��[[�h'���)�{y�j��=�u��u�m�3c���e�7w�=yW��{ 
to��M���{�Of�U�^��ٷ������r������O��cc�{{�>�j���mm�o   � �{�   � {�x�\���H���M╣)��jB@�X�mE�/=���4�Y��n>��U��B��6�dﬤ*���}�J�i^ؕ.U
I=�ﶹH��K�IU7��%�1�>%�>��l��ޛMR�]���M���%/F+Ƕ�E��R�|�^� $��m��Uty�d
���g�x=[=C*z<>�^Pz>�z�hʫ-l=���{�u���kl�9�v�K���N�k�L���
��pU�t��}������tzr3W�iT�΍��
w�^ر����J��oz���Yրٶ�g�m���V�hh���ݺ�^���3Z���7�po�4��.�8���P��<��2��^�^U(�ttv���h�Z������:��_Fz��[��� ���+�����>��}'m(_c��֭��}�s��k2�Mm�f�^�;eH:�ۥ�����U��h���F���t継�޵يݏ�<h�6���
�hu݊��ﯬ�5ʤ�w���<�m4:4���}&��uli��_,�����<�nm�7�s��t�j�nFQ��}:�t6�=F���a�����A˺�������ܪ�Ӟީ�:	��*����۾�Z�u���i��u,y|�`]�ӻ�x����m-[e_f*��||W����Ԍk;��B����ɳ-�sk�FM��2)}{���{7��'�l�o�}�:�,ι��sv��>�B��k��}�b�����Jz��g�zׅ7`�A�e��M��i��m�cE�X
u�	�}S^=]��׶����\c[aӏ����`��;�kU�ݚ�c�/�7� �fSK/�����Lg�z�L,ȌB���wڕ:�ض�t�Tkl�v��a�S7��M[��s��@ͨP�_`�֩����}sml6�ԭ�Qm�J֞����c�V��G�f��vr�Vǧ^��}�]��c�eN� E?LT�@   S��$��� 4 �i4USSD�##��T�R� F F 5O�"5R��0L0�II	2���2x��_�����_��?mׯ(��ڒ�[?l�ys2+���,�1�`9���kR���Y���`P*���]��P��UU�(
��UC��
�(UU��
UJ�� UB����@UB������UW��*��UU�P���������?������Di�{X!=���x��Q3&��Vͼy�6�=O������P86�X��p@4ʼ���nۋ�JE6I[�iF�̽�1���B���Ё2��}��=`�H����;����h��؆�WsݖT���A���LXj�_^�N���\�b6�
���B�7Ͷ���mi�ŀպۛz�[� eK�M]�C��c�޵����Ț�#�;K����Xأ��G�p�(	�J�.=��]}
�q���r[���н���V]�\3���S�^_=���緕gb�p���:������W}�x35O��a2�b��qPjgjӼ�%�fܓF�&`�+x��H�1�Os��^���KȪ��
��
f�ksvA�[�S�(��2-#�3Kq_vk��Gu�C�ͨ$��zewY��j��:�z!��N�e��bU�s�[��k�m��<���n<;?t9M�ڹ�{+��M:S��kq���.�VMEy;G*^�!�sq��b.�`�r�f���y�����8)��֬��P�uuo�ѓӬ�k,<�Ԯ���o���Ʒ�2V���[�*�%֜�d�� ���4�f�N���n�j�G�j	F�ގ��	6���%�W�)P�s���u�8"z�gYV�T�5����]fmK�4��jN��k��ͺC��]M�g�}�aSI��y�Ƃ�Qo���p�la�PX�/��T���x�s��*[�E�V������OڻuZK=��A�0�{Qݢ��kF4{s�:��Z��m´���g.�r��6�"�sl�/V��lQ-�D	��av �d[ׁL�њm;�Ed6���I�,{F���a���az�]�ç��.���/��Ga����0�;y�n\�w
�Aۦk��r������@��^}w#���?'fN������Pn�i���p<����n+o?'�c:�Y�i��89!��]2>6K��kǲk�����HWj	3N���-a��	�A-~�x�l�T�)M��$aK�T���������<��[�s����ћŌFliC�
�6C5�⣿D���м�XE@EE���Y��'z��X�fs�n��Kfc +����窿h��j���<@�gkoU���	�C�4�F�CMi6�,�F�g'��]W�]n�+7�L�3*{��/�%OU�x�!��˻GvSpf�d���sd|��C�sE��6�ݖ�E�� �qbX�٤�E��P��a����E&�&އ���]���@�����V�$b��BՂ��+^�D���ZD�įo9�o.,��N*�ld<��jɞq�]oe��s���pۻ�ʧk���0V!e-Q9ي^�7*+�;n��<�a9ZŮ)�7���ֈKvfl����B���nd�vm+C�R�H�a�β<��F�?-�]&���~p�L�T�M�F�\�w1����۽�W ̉A��i�v������2~�j�IM�F=^c�m7f�����{��Է�S�r��(@x��3͞�gz�dM/v4r��a>6�q� ���947�ʽ���U�QV٘63&GoF�ֹcB�w�-H�dH�Z�c���9��8.6���F8^QWf�b7��4�UĀXY���<���ݎ@�WaT�Y�گdX��!Z^yJ�]j`-�lJ�n@�C���ֺF����BR��ήZ�ދ��Z-��T�����3� �W���l����U�s^���uH��u�ߚb�:��LJ��4��j��d��w�Z��,����+�LWv�
 ���Ҧ�X���md(mӏe�P�*�P��%�	�V.V�Y[�7O����˕+O�z�U2J:{��PU�%-��z!��\'/����a��;%��Ɲ_Bfmݪ�
�eT5CK�r���X��ҁG�
�-^���$�k��B�����vv\�G@m�-ЂN�z�,݉r=K��D`��!]u�4�L�{���R�p.����pxa���E"�"�5CH��ƨ@Y���j�5C�P�P�@x�"�"��Cƀ���l6���}jtE-�R��x��e�nw,��t��]Q�����6��i9]�� ΅�vt��fs�ߘ�X�`�މ�˴�=j�wJ���_<j�5\�.���at�fK�K�%�bԒؑ��]X� W�����	�[EpMSS�g���&Hs��P0{j$2+�B�Kmu��=t�ܾ�>��-)ZB����ju�7]%�M�������ANo;{Z�c1K�-t�m��r�ossh����`P����9��2vX��^�òU�6fNU���iu��4�9vv��p���Q�qm$�0� X�r���h��&�VVfS
�d'�C�֌����kq:���k<G�Տ_�M͂�a��w�;r��r9�a�,�z1�&�w�x��.�Nƪ$�R�⹧'-Ь�	v����λ*��A��eh.�܌ S��T;P��yjP�����U��%�E��Km�İ���ౚ��}��VD�(���Y)xDc�̉ץMN)G����n�'����{�������u�7���B�ȯ�����Il�ej�1�`�3�f�v�^�'6��[\:f�
�v(�ܡn�����m ��nZu.�,v���m��zW�C�@" ���<��5�c�$�l��nr~AyV]7�33/��Y�mлX�DI3�ض1�ĶÈ,_����N�뽼ݓT��s!%��{��9��
X�F1^�we�4�s����E�[6���G���,�lf<���M嗇vƛ��ɭc�]$�Wuw�St�c�?X��������Jud͒����J�y�P1r]H��u.`���2S���R4h�-�Z�h����5�M{�QF�76�3QC�R#3.��6^)�s� �ڛoUeL,�(����V�:F�]=FV8Uɥ���$��7wLf�K�G@u��l'V˲U"s {�4����n��Ib���E^V�wk�L�w�s�����f���kj�ǪP�nA���
�R�*���T�&V�n*Z4�؛Z%�bF�����ld�'P�@��OYSZ�T-��-"��6�N�$bgN�E�R�{�%�����x+ ���\׷'�q{b�ˬ�O�֋-�d�&��߽(��<��|�zn8����֏���	�^'�f�$�=S�W��i�����hY�RHj��]�B��m��;�@��I+��leM"Օ,��&<�Q	ܬB�^@���b���l�G�ja�kw�[S`�%�2�ъ#v�B��73t�[��J�ý�o�X���a��{L �)�"oF�n�
�6)�������T�OY�!���)���E���7d-�'�۩3�Yӹ6��O%�jñ��y�vL�[M�o--A�A",�WH�p"�s"zVjy��34�����i]�l0���ҵL�bB��í�����_8k��P����Uq0�E#��f���d����]WBWI��L��ԣ�!R_��]8L �=iۓ��ɗ��������7�;i��3^Zj� QB�>��u��:}RLܴf$&]���\@�Qb�.�C��f&˘�,�5�m1�c��ɖ�ofv�E֮��Ԁ$NZ�pFlSy59VwTaj�W��{V����6Q̔�C���NI܉B�S�9��hlu�5|i�~�J��]�%��SY�kf��M�o2�H.�i�]JFP���"jұ �b�m�����r�iIt��(T���Gf�cr�m�W*eƌƥ��^IxU� Ml���!��1���Ԉ�	��k�����P���F�M��`����*k8�5wK q'r������%��v3�����ƫ0P���wgEڴS#����9y M�̲��nb����1y�M5b{$�s���u�KF�}�*+�ٷ2d�~g�hD���4c���Լ����n�SF�ՉS&GF�oDHcg��$3��b�,��lN0d���4E@�Z��+HCV�k��/:�;.�͖�rh5�j��t�ڏF;�)ڻ2��]���n�e��%�.	��o5��t)��b�N)�0�Ee�#$9wom�*3f����<wW�[h���B$~�2�	MV�̀]lw)k�j��I:1@j�p�)b�������(2 G)PU{�Z5{(dE��K�a�ݒ�۵��(ջ4mj��"����b{�*
�;y��xB*����ؖ�ۙ��	75�O�����$���\�&=36R�iP�z;�N��*c� �W��dP��##�BQ�[��2 �L��Wx� @"ۼ㏸R5��U�� �}�����fu�=�mjx�#J�M:�}騶���LZ�劎�1��n�(�b����ׅ:���\^j�tp���t�������Y`����:���Li,0���S�'X��3KJ�:U~���(����t��\M!�C7B�Mw]]�՗�Z.8��{qvA�����I����+x(��+vj�[8� KK7iK<��'�KŻ�Jj�7�wm���rT76��-����n� j��J���6��x�����=��1��u��/����Q�Ҝ�L}ʀ�Gc���«����ZjҸ��r�=����)l�E�4�>�Pur�e�㐰7��}<-�+�a��/i"� �-a�#�Vʫb�P�Y���k/w�Mo�K[��f۽[+9�j����;�N�e�'����(Z���R��`��ؗ�=�0���s�<շ;I*�?��������e���VʸJ,�4.M�T���%�vU	s7�ȊE���5{x+e�jZ�g�G�8��XN��=;׆>c#�D;@~ �GS,m8�R��Q�m�p	��z���B3&�O��/�X=73r"��4K�{���o%�f�?��hU�CN9x�cZ���b�婝���MV%���3\��Й�D��I�B�J4�1C��Y��K�ձ��ӭN���a:���*Lw�/�ï���{t�6 ��y֢
rh:�d(���?�D���W0�F����m:�<�G�g��D5�\��N��e�3�z�	�s%�f�:������-b�*%.������ڙ�i(py�T� O\��ؠ3زJ'��]1�ɹ"�s�,7J�ntY =Ǖ+ZFխ�T�蚙�'�ii]@�Q�ek8��F���\����,���:�w1^њ����{xrlФ����N��\�
z/��ouiĻ��JLH捣{�S/Nэn@A~F4�g,Ѥ#�(
;���!�4!��)2�m��R#n�Q�v�\E�c�4AN���+���h��<�l2J�3n�T�bY-`��:��je�	Wb�Y.УG���,��f[
��iLȅV�@J5j��xV�Ƒ����sz]�e�K��H�s�:���,�3<Q�m޿D�q}�O�:�4x�-��������M]�KZ��h`��0��po����}c�.� ۷�T�<�7فQ.�C`��l^X����P�%�qwI��HF�rkl�������ID3%͵�s:P����<da������9��ݩ���p#6,�wj�;��uk*��A��L�I�D��
�������T;*	m�X)[z]�8�(�qe�/Gv��;R�/18ɕ5�E�[�7S�	�J�=q�S���l��#G�fAL���5��[[��4�ͳ�DyD��JW��Wu �1�+�!a��d��Ź����0 Z����� �Y��UmA�H:Ķ�԰�6
ģTm�l#y�A�Hr:,ʦL,'�KK?
x[�����Z��x�M�l�:ĳ���5���Xە�9��鑥z�i� ��ȝ���{,��)˥��.DZ����G�Pd�����i��uA���gF"T5�jⱓ8эw
AI1k��
�9���t����(w����Y�{�fI�]Y^��wo5��t�f�f�j4��4�*\��{ו�u^�v�6���f�I��l7F�cv���5�㇭��5��״��`�>@Qٵ�V�%	�����X��Xf�k"kO:�Q�F[�K��A�gfp��K�8��S4\�����-Y�	��VU=r�N^Vi1U�&�b�h7$
�1��(�R8��G`X&@y@H1�m�n\/�S]�-h⤝��8TN�q-D�X�m9]�s"�ڦ�ڼ<�:,��
��~Y��$����[����(�6n=�on	+1^�=�Y���O)V"Q�m-��Ʊ'�
`)P�n�+Vݽ�nk�����}�a�v;tnT�y͏�h�������H�<&z�Z�&���kI��۷4���Y�q��E��x��)�"R��.�?��S��RזS�� �yfEd��Qh�sF2%e@�L6֊�����k�H��6�"�\�0F��1���EӑY�i(�sQ�y�9zі�x�x�ި0a�SB���GcA<]*�pU�FQ�n�P�;���ҿ�;w�����N�ʻC8�ܦR0cK]Y�k]�i���`�3*�o��땱e�$#d�~R㣄�`ÖFB{1G��1��xȼ+��V��[�g��w�X7�sBe8�(�-�d��B�������7��Tm�/n�%S�]��W{7����sV������S\B7	}�^��1e�N<-8C2��Y� �-����^VR;:�B\/m�����h�ɻ��J�f��8��e8��RKT�ι꠻�H��1f�繐Z#�r����S��uj���o�   �@   �ʼ_�� I   ��{� $��G��$U�t�<��*?{       �2��/�0           �                        
                        C���f[��sf,�$Ӭ���w>v`i���j�\��sN�7*-��U��&�Y�����hI���͡�'R7�"i�G+���2gL�WJ���]�[���#���8����N�:�>���r�X�>�⤯w�*Y�vTo���Iu��(L��ӝ�4�>��WN][Ir�m:1�_r֜��$�{�ހ��RXXM�%�#����΍��ډ.kR�q4�GS�ee�g���-�ff,�+�F�mԒ9��2$�*�5k7LhcS�Bu"^�[)�Ќ*e����Ƙ�*vwb��+md��o[�.@ʌz��8¬����f'jI�£��������ǥ�n�J�̴t"zc)��T���ǖ�Q����dis�sp��T��1�P�D.�0\���-�X�چ̶��j}k!������ߦ�+@+�%r��vx)� l0��G4e�M"��o�l�Mzl�gm�I]��&ww�Ӝ��G���{b#�聧f�,'JT2�^�Ev�]��xOr�U��8�kr��h��Dk9_x��mTy+��������6�;�������QSs�}��5x[0Ǣ!ˊ]���	��Q4i*(�ޔ�[0����tN�z�"�MQ�E�I18�8f��%QH�徹�_p�E3Ș�fm�#E�>;b���Rz���i�7#��(Eb	��{l��{���!'�ex/n�p1�1�,����=~�	Q\�Q,��q�M��:����3��P`L]q���뒶�<��%ɬj4C vb޻�I�޻�-�E��Zm�]P=�X6��m�ˌ�C�庱
ʺ�^��[.����aP��3�`�g�ڰ�����X͠�x��k�E~��idJBZ������	*��&������{����g�׌�G�Z�v���M�[��Y���W�"e z:ɓ�.;�v�2km����fQݬ�]�m�]�TzgH���Mi��dZ"2��#LKZ�Ԕ�~��Z�X[źa �U �����f�S�q0�]�7��n�c쀛6mI�Kݫ;7C>�d�8F�	��{�Ų>�Q��ga�����$�����i��d�6;fexγ��\m�D9�L�5.��.ACv�?ǂ�"�d<ӳ�H�HG���A��gC����΁j:@�=ן�dPE!_�
ČDW�V@
)]֩�d�M=
�ab��t��nP!�.�
�ǄR�cK����#oɛ�&�:��JcI�����.��h� �%�l�F�BD�L׮k�ϓ����Y�	��2�,~=k�Ln���m6��� \M��-#djQ�_�;(�X�Xx���lf����a�c��4ˢ:��4�
HR�A%��r�;l��o�q�yl�Y����tgj6�M{
�«�CU�і֤�0br�J��#J Ll���=���.<*ҽ̦�b��S͈XP�z��㍠SG2�]o���Ol�r���%��?m�v��\�!)���N�ݞ�8���e\��r���ؤJ����k��;�w��ޫW��Qݹ�yM*��aMY����[d�L�:k	梕�l9�P�(��g�f��ʁ�By�U>�W=�s9��fI�;6���$�-ز��9��Ⱥ�rn΂�0)s=%�h�l� �PD�wui��W�GAi��*n�8�q��7[V>U2�_X��6!�cŎ������_�>(�$��n-$���:���S$�AI5�k0lX!Sx��lX0��N]�=��_�%��5J�;>�٭��ֵ��1���yO��/���w6RV6��%?v��7��.ڱOO�[�ܬӈ����, ʃH�R�r:�'Y �m�%�.!8��o��X-�]���o�`���3kF�H�}�Wn	#�l�� R�#F�ю��s(t5��O௱�ͭ���Y�8���L��U�n��Ĉ�|lC�şYnL�ǌ��86O�>a�+.�@��Rgj�۞�,�E`��9�uѐCkw-���<&0��p�D<A�vQ�z������{�R��v�Ԇ�H�J�mc�r���.����^�]�`��<���qP� 楴�f�@����������U@e��l���
�6螎B`��'LX�ˣU�垇 ;6SbN����a�l3a"�Pwg��#?\��ڻ��o�$z��%1�Tw�A�d]���ǳ�֢ʰ�K#��YZ� �qj��eq�Nݭ�����#z���X���Kˇ)o�J%"�1)��7֓YZ���JEb�C��@Y�U�2s�U�Y�#  )�'�����#]!{���z%�~eK^��\0���"os���7��1jە��)-�<��i�]*I��9�J�C7{&�Vw:����Áb�kM�j��Q��|��[��̌ݐ����i[��3.���B'��9rE�0z�$x�1G����)��Y"��6��}م���<i���I� �^�;��;�[V�rF��Ѫ�n�v!T���F�/�?$�d���~P����-Z��䈆�R��p-�.�YѴ���0���aY�k
�9�Ag�\����qg�A�FXR�Y���Q�SM3�������G#��W�xE+7��'y�:j�r�gE[��J��m�dp�B$���� ��;z�b;2`���OG�cJ�&z3��9�0CZ���*e+��9P��B���=�aY�����Gr�~���y-T:�B��<��R@4B��^ZE�;"�=0�51�?����*̼;&"�[w�i�cQ���;�W=b��v8�=��$#��x=J�ukUg�p�!P����֘�VŁm,�낥+#6%��Rם^�A�SӉU�z?v�4SZ���x8����E�ݗ|l;�M=B:rdf`���4C��aS�l/E��/:�����d���Nb��>
l�V]�h��v/�{�0bqOL��YQ�rV+(�F���;�ȳh�����(+��0�ؠ�c�** ����X=�o+_s�~iW@zTF=wNv7g��@�����w��b�4����_h:4A4�E��.�ܚ��ât�LU��:>���Mn/�r���&ო �⋕Uv!�т��Y�k��Ѽ�DC�c��^��[�j/�qU���H3|���lF]m�dP�v[HR3�,����́žf���c�!Õ�ȧ���mK+����3�*	J"�v�p�#h 8Er\���U���q�4F��q�%�K���k�⚞\��z��B݅G�[��6�i���j=�j5�w�Q�=�}�]��E0\%�]tV�=������MZ8�}���+��8�RX2P�:JU2�YB�u�e��7��-�Z�,��f���8B�sX?�����c�qA5�3�1�7j���+�:�U�yI+"o��6̓Bq� �v�eՋ
ھ�w��)yT�Ih5�Rm�f�^�P�7^�[�(i��N���^r{Z!��}�T�Xa#T*�b�[�֫lN��tF�z�&�~���6�X�K���
�΢�2u3�iQ��ggLkt���7�sB����1����F�eI{����B�F��qXANMmɶ�1�����`�Ur��^���E�����e�fd%Z�*�L��w�������a�m֤J��.
��߲č�03غ-M�JÃ-U碒�fhV\��!U٫&�aA���K�B�0�[�&U�(��f�#Dj����!��Q�s{W����F��[���-�I�pXGI��-l�g3V��7�EF��P�bb	J�!�v���f���v���!�-Wف��S�H���PiJ���(ee�[uj䉀96��A][�ܫ�t��^s�ӷ�h��|�����l���V/&�+��P+NLv"��6��F���/vﱙ͉�z�Н�2�0D�����f����p�vs^��/K��B�h,�!���@������R2�v�h,黦d�o6� %A֖T�6u��sF�)�t�Ҧ����מ�_]fT�*<:9��,�^`N;�0EO1iu�5j�^�í`�C�ᬶ F�:4�Xr<�A�d#aF�1.Jw�\d�5d����J�k2,��d���.^�]l\�ɧ�A2n��y�;WD5_['�H �S�jq�&ҍXC�52�$�8�j��Ef�!�Ra���W��Q&rHX1Xܫ˱�Փ���l�4֞��7xD�`$�w��t���wB-�r���5�K�j[���p7�e������f��y� `��9��Z;s����Z';])Ӓ�(>��_�^�?�^���b0�om��yU�Շ�k �R���yD%ˆ������{)\;+Y����טF�̊0'�Tqe��W.P�Ŝ�Q���3�pq�4�1��*m��^�f�qd9 h���)N�]�%١��ݓ�gv)c����ʛ�,EB�mh��CQ��F����œ�!�*�S�a-j��U���v�]�`*�Z� /���¨5��.�ȸh�z̭W��;�a���C�j��Z�sn�"�^��Ľ�I٦D_u�v煵I!���9{��Lxg �3$��{c!Ypai�F�����\N�p�Q�f��,fD�I�c"��� �B
�9�~:�m�hDEa�&�ij��j��B9Q#�K�:��6����o��O�#8΋]}����h�5E�!����B�٠��jц�(e�7��e4�P�.ug��C_=��*��&"���ody�� I��ԏG	O��ٮ9ah��+1��b=��\��ǹ���c9d�w-2��k�8g�&Khv��}� ���R9�Fa�J���	׃���r=+3P������q Y찪Û*�\�EjU����ݎjٰJ6$k�\�[X�qcO�ξA?5���=7�s��Kh;8Z�!bv��ӛ����ڸ��c4ll{k=�:f#��r+����V���Txa��qmfH�+vrүQ���a3M��-�b�"�pEsX�w�K63L�u�,������+�F0T��WO��v�u�P�i�pY86��ټ�'v^�'�bۼ�:�<:b��K�L"�4��vV봺�.�������7�*����	V��� ƻ�b^C 9��{V@�SV�b��v1v�j��
�x�]�w�T��5�̥j�q����Pjña[}���6��)5GL��Q�1�d`Df�1}|��s�!�Ȕ��ʹd#�TE5� ������(�je�En�Ҏ��j�O��/]�ym��M$��t
��؀1�ѥM�u�� ���V,9�测qಶu�VsX��t�dK2/�B��<�(d��V�@�F7rm���o��b�(ZDՆ}3�=��$�p�	�d�5\�i㐪̵P���������<]ɫev�%�OO��	8є�[��5:��9-�"|l��:b�?��DG�l�����ZFZ�U�,3��[=	�PY�!͛��2�"ީ���n�E^7�Y7VN;��N�2���f����;"ֲP�0�yBB}+�X]�G����rIJ��%��*F�v]H����#���V]1�9�[wu{f��e}aٻ���m����
ۥ=��٭	�p�e��s#s#�1��eM���T�Z"Y��+��/*Ӿoz9[ٻz߶�ݏ!�� !)E���51D�D6O��*at�%��������*�LBf�^9��=�o�[v���ogU�)��T������Id��h�`(���X�2R@�䟄�v�Ы�Q�\2����9?lݸ6�T�"�G��m�&;�h�m��n����O�׹E7U�����@�(X��`v��p"<�g��^|(� M.0�F�ی�#�t���h�,�����)DU�r���u�Qgs�r21�R�z�ӘH(�כ�
Џ�s)��@�2�v���ܺ*���X�ʰ7�"��i���_��9���v�`�a�r��[�Lu�p�*��qe�]�p(��T��Z��ˑ�i��hn-��	G�EW@�%4L�����u�̠5�á��K�3EE){i�F��q#L�@�#��=�oV�����$�ykZ	^�Y<Z3B6_)tY�-R��(V�vئDqL`�I�r.�O��5ffB��8q�[躧�z�G`��lJ_*�{R�/w�7�(z����梪K����hzn`S4e`p�g��Ҿ��V?w$*�(rj)���MNPMtn� b��%�3"dy0��y`l4�팗%��c���W��쩷/�	T������H��Ii�8~a�5:8��%�"jiܱ	�E/�K/�Q綵h�Ҕ;�a����Wʻ(+�#�gN�W�-�O:#��E���O^Ǹ�6FQZ4Z���څU��tn����V��!����@��Л��R��|�;��]<��]�C�U���S7��m��toţ�r*�H�-X&�re�a�
Kݚ�rTF��O�Ż��J��N��{p��/��U�7��VmB��r�c�n��:7���Z���V����k(�8�0�W�-���{���R�3"dg�_�u�(�V��laI�	9�;zU�����ȯ�=�>:���}|�� 
U_��P*���+� (B�� *��UT�ـ�
���_��D��ɿ֍����w�0]�̬���ך(�fR�{�[+�P3M�G��k܉ĈN��[���{
���rZ�NV+� �Z��	l�U�ɓ��#��yuw��T�+�.f����/��$��7�v�b�#{�;��Z������Y�t�&S)��1rV�2ԑސul�oll�N��>��,B��޺�NR�Y]�����C���-I��uJ�S��6!��3�]ٗz�v^�
Q�,B'��H$&���Kq��bȃ�ɥ��"Í*4/��Ը������#L�xݩ1F��R�q����R�k�p�W�T��T*���UD� P&�Q"� EP��~w�r�/�;��.8XV3˫(����U��n��n�s��Ov�a�IZ��F�f����G�L�Qa�J/ZF��й�i�a�/�����6��oН��K��r]$<�� ����e�$)
��Dg����y����XMAe-�.�Z
rc+Q�>p	"��B=@���A<��0��<� ��� �R����r��p�/�,ձ<���c�EJ4t'K[8B:�����8k:ty�+R>�}��"�=cʳަ�4�/tCl��o=���9D�/I7�6ɱV���M�][dU����V�hT�1���f9B���Uz5�&7�R��OPb���l�G,m��^���X�U�x1pc${շϚr�ut��
�rb�=;M�ܴP��Y��x'�T'G
��N�^'�V:BH���J�[P⬮�53�R�ũ_Fua1tϾ�x;��0cuq��X'{�����,�:���K%��Lӳ9����!t�`fD�U=�нFyW����+�h\)�R�D��#�����h�y��h�xr��%�c&GG�-Jn������Ҽ�FJ�s4���2��9'?w.�M��39˽F�h�b�Έc�m�$Xk,',���S<�pط,[��Dǜ�
�����={˾SVڠ@�T� *ˬ��dʀrW�q=�2�� �4�dir`�օ���XJ&�+%Y���K �vh�dQ6���˦��G�7�DE�n�Fj��T�C���1>�*�Û��f�=�I��ۡc���J�����b��2�Td���ol������g�����1~h;����3��@:�⭊:�K��e�T0D9(�b'~�肋0 0 ܰù�u�`���P=h���@�^��N���K�$�s}t���wZ�]����]{B���7�Юҭ��v������@������j�~�,7�̅��?���bk轼����`߇X؈`��m�!WvA�S�Đ��4�&���o�Tm/
�һVt�Jj�d�R��s�K�օ6OWz��'T�&�iѾ�\4I$A�8rs�kG�$�ﲀ�	=������W/r��R��4�Xe�uǤIR�0Q����N��a�Z�1��(!n������r��4��4Τ��F!I�Q$��4O]��Px6` w�OQ��n�q�t9�=��4|�u/�̏H�r�|0�<!n��<h���"%26(�Ё�LQak�J����{x����yG�j�_��T�+W/�p��'���3Bf:�V���B��$�;�|��H�^��)��)[y�o�EC���A(a5è1�Q8X�����Ux��֚����Md�*� E�yK��
��v�:9"�w�����������\[y�-��5���2�-B/���,�����E3�v��N�ɚK�-�+���34��܌�q#�&z^w����M-�f����:�o��և�������^Y��;���,�Ŀq{������Ga"�Ր˃P��h6�p�@ �<+|��e�tpǏʴu�m����:9��D"�yR��7��]��2�B�JtϺ�p&�p��I�Sخ$|��OUN<5�"cD������7��Xz����5�����ڴĦNI'� �~���MF§���L�-pIx],LN�!���գ��{I$4�;Ss�<��qi޵%��h#��eA[�<n�ݚ�h�qi[�vV{��nQ����W��G�����J!(^��)*+��> G��^fix��%�A-�X̅�&�Z��ǆ�x��������� zthx�x!ԛ�3N������]��?:����X��	��m��+�JG.���!B�%���
�3ɭ6�.֭���E�*/K�U�����7�L�FM��칕�u�U�.�D�i�4D�c�Yr��&(��aS�qZ_��>��0Q���՗��_q��-N[0�!�k�xV�h�Qҩ�0�p��nW7�������\xmm��%���ƥ�s�YZo�9�	�����.n��MI�Gmv�s�9L�j�m$Ⱥ��:���d�3�z��g	]Fu�xa�j����mL�m&��B�h6ϵ˔z��ӧV�bs�x"�>H��V�x	I�N��������N�<��P ��G�'e��E���`,�뫊2:�,f �`���������-b�+C�p�8�'��b�F+����jtX�av�~]�'��b�jxV�ֶ�e�#��h�A��H)V$�ath�;�x�D���{^F��Εؤ��G�O��{0"���H��(
r��;dxd��$�n�f�R�0za�D� >1آ��G3��Z�OT�"��y7���ifߘ�s?�X�y���uk�:�nic���]l�'�	�8�Q»�T6mKna�^���zRv�Q�M��J�/D�~"���d�ւ&|�h뉕Z8�#?>m� ���"x����%֟IA*��爌�\�������U�tjt�q
���M�ThZ^�7t;C�;���YZ�)>����y�v�B��Л�p�-;��O����m�!#{����ϷR�P���˹T��,LV}&��%��Y=�ר��c���Z'�ھ��Tr��hxtT�޸LpJP���K�]=��):���*��;q����g�Gt�k�;�E9�����-T�F�Zx��vf��Bx+��Ȳ��ug��M��A��`XAN<r�:�j��xRg&%~PX�8a4|�t�O����ex.6.k�Ax=�9.��7F���#o��1�X�"��i�;F�QZ%gN|���f/���� �[�c<@�}�{\�xb��Jo��D2ϯU�&�sn&hi����;��Ut�8s+���`�Ǜ|�_�f[59�j�$����G��.�{���h71� �;6��Ґ<Vp��AsIx���
 S"�3($(�~�pcr��%�.��|�k�:���:vg?8%�:A�JO T�& 1�\���J�$UZ���� �Q�X�f���WOz�?���f����@�yB�~�sa�[�}����E����yd+�w���ḙ_'Ta�0��/�1�����q��C���f�٬.����]�VQi;�^����v+�^�P�YE��R��8�Uۉ���2�Ve�*\��<Yj�w[�:^BqqXX�7ܫ�(x4��i�;kZV��se�|hw+1�H��T���%��7!c}����/�Q���T)`���3+��@��z� Ve5�� ����y�N_�EWw���4X#؈�h�����vH0t&�ww%�Ds]��)w����T7�9Vw���E|x���\�u6�@�����ċ[�CF��d�N�lS/��U��!�f'�YF���H��|V6��.�b���.9��Ю :�P�c�1b���UuTF��
�{�����d=JMx����"�rj�l�S<��M�H���V*��������@֝���'�{h�ݶm���ՓT(�%��
�>TDF^��+�i�Z����_%�N�%� �R��Y6J�zxT��.��������܁�,弍��n"Q2*+�@mxh�9�7u�jE���i/w��)dCkv�TG�B����3�	/��!�n�Y�B�+�����绮�&#�[>b�7BUmQ�E	#e���
�'\�S�E��Q��>.����=0f�*�()@Tv1�h�"/��xT�O���P[{`S�/Ll?*?2����N;??�����K����lm��ͳ|��3��
b���KD�2��I>#�]'��x����	7�aS�X@�E�Ye�&[2�^:jc��5bx4=4۹앎�]�u��e���jyk��7j_�~~�&HVFi�`�܏�>I���`큘�z����;�3��{���>w���](=Ķ�=�ί3^fݵTdv"?N��,�5f�%C��3�j�"����v圧S/5`y����Gu~|���z_�G���C��X+�������B;,���v&]��u�Aj�+�H�\1�OO\/{F�+��E^kV�3ʹޝq��i�U��N�'�z�0�)]r���ui�@A9ԫ���Nڸ7o9�-wT�H�w����Z##���>K[4@';��Y��¤�i�e��Θ���`�V��2K�f�҉��[V^�4��"�^�;Mָ�C2��c��!8���9h�!!�H4lhVC���=�T;���:���%z���ף�C�޵M�v��;�g�4_(�ړ;�*n�*(S��͑�$w�״�n�ƴo:1�:�u�E���	��g��o�Ռ�����$@�r�������^���V�p�]\���Lf�A"@��,�4M���@;��E:�hj�6+UF��H� +�]�D]c~sQ�XO��\v��]�*�Y�k��'ǡx��;���~P�v�bf~\0k�mCPW`��k������q�#H����g��<��!x����k<o,&0�Z=�F�Bt:����Ec !�e�[�:�+��	�F=��bE����T {LwmV��`Q�<�\=�ٷ�ԗ���p`���+� :��6��2�u�(So�j�j��y�?bo��ƻn����zn�6Ū�T�R��%��7`�\������R��BF2;����L����K�M�!VO�����$F�1�ʉ�+B�kP�;�l�/c�`&k5l�yÜM8�����R�in>�#c8���+�j����-�-�1سz����YSs.����qs�������@o��0W�uv�R�h�b�O9��T�}uP���ӛ��'����7�{}�x~�i �ķ�t�`�[g����R�-ۢ�"�krـ��u��k��N�x�p
pnn���Y�b���
)��NnOeW�еp\�f�/���u9u�	�1X�ɒ
8礀���hڹ�6{^���f�~/�O�6�;��Rb�Z8e�\|NWP�^i�<��(��3��%yqؓG# �K���t�D�t/W��f�<�ˢ�M�skE�e�M���_��~g�e�zZ���Lr��ӅQe!Y/;���!gk���+��=�W������8���k��˵��8��I�D����굯�����؁��t���*�����<=~AõyTN@�&Y4�"������+.�!�Qԩ JF�`�{T�z�.":�#�\��P|�wF]{�рd�~�.�loE�< ��G'8$>n��-PE��N�ZȽd��$�[^���P��i���"r�5ش�6���%�nl7�B��z|�n���.��=-������L|܇��`�UƓTJ+�(/�@Qp1����,׍j{��xt� tn�+��VL۩���γ�P��[�2�َ�-{�B���p3t:��a�����wl��k���ڷ����㇦���S.,N]��*A�v�Ƙ@�9!�h�Gƌ{웕KڰdJ����qC��:Yl,�x��+��D`*/pVsn�KCk�V�S�N�I� g��Ek���ܦ1VoM�M���n棛����Kadm�}��W[8|+B�EL�	�
C+݄��1�YM�H����}��E�vU3��H,�K����8�\���ër�C��M���\ݜ�]�Q�͉C�8��I;+n��k,iB�#�`B~�$�o�P(��<1����+����GF̵2�k�ѹ��
���X��@#���Re�`�Sq���+>�r���3� ;h�>�Q��\;Mx�½����ř�����cB��)�:���W��W� \[�b3]ן��򬄜��7G	8z�"*Z��T�C��,�(�r��\B�f�!��b(�F]�X)�� f3�첝j�;�,�Ԗ��N¿\y�[�����fS12��$�忘Q�]#f�v�v�	���Su����{��zuB-aZ`����U3���s���Y�d�j�%o�^�����+p��0��f	����P!y{��r.����]Y��n�꾫��owr:s�-�n���Ē�ֹR:i�a}����aN1$�Iܻ��Ki����,�r���g
v���lJ-�>r�4�B@�tV؋ٙ�����,u��.H���K�be	R2�Wv5F
e��Ș썢���W�Th�p����E�w2�w稖!�ITeuGiE�L۰
6���\X�?��� ��_����o�#r
cNCA���'X��p�|ns>5뵕�b����Z���'���a��P�k�U��5�t����ZS�@��whTͷ=b��]��>��/�K^����{�D޴[�Jb�4a�*m�����+<~.ڝ�h��E�7>2����`F����ʙ���b�N�:Ӳ�
H���K��X�E#�=r*f�E���2iBv�iM[�(���k�6�H�I�yx���Pi_hc�4a�-r�խ���؞�N���;gЉ�^c1�>y��R%;�kt7W�^�87O�AHPKu }ej'�`g���N=�b��G����E��V�X/h3�m�N����i�$YbJ�c ��5�Kqÿ�0U�8��BEj��~��-�($�����ФG�� <s��,�s���1kcP�����VZj�m�'��RZ�r�|��W���S|n�q�´T�A��C1t�i�,f��f�ˤ��5��P�H1�Tozt��$�C�����T����Z|�$r���b��=���?J�q�Uwz�y�Ĭ��XʳZj=�}��bq�Z9�n�.����NS�'ui|:�����\V�J�?U���p�YF�um-$&�	��Qk�/��J�J�Emur��yf���n㮭y���Z���X�u��[�8�l�pB��'�VæJ���xu����U���+��*�����S���x����mг�ÕL>Gs-U0�wpZxH�fO�r��C������Y��(���S��m���%��M,G��C^S��i���p��鼯	sA�wm:�t(+.,}c�阞�[�equ�]t�Z�]&�*��|]�H�����ڒŕb���'y���]��R�4.�]
� �*�W�u��WDH�@�L�j?vGx���Y0����N�9q^����۽��R��M�jQޤ���[FX��wWywZ.�G.�'5�H��W���D�&����n2���������c��YߣL'�|�r�E{O(L�'cUrn�W��q�d� ���y��P�㖡���}7�/2q0qIn��Y0��(�k�r?��@�A���>6�8o�-9�b�Qg�nDqtk�+��.�SFbĒ��|�nyXDc���F�r�vu���<���2���Z9~�Er��rZ �CT�FY���������YOr���]F!`Lނf�B��^T���=z�SNK$�@�;��شw��y�����VP����׽A��o��N?W��9��n��:�>7��,�·3�񞿆��,]�l�L�nmAM�/�      �@   fY�=~��J��,z����I*6��8�u�A��n�Ԧ�9)�#*��{6# ����nA��6;���U�&���*������:�u�,�V4�L�E��A�j�˓1ǚX�=5ּ��ܖ�X���q_�B$�����t0-TOg�#	%�����Qv��\�LU��V,P�b*�
f�̨���W��u!�q�	�e����{��R'@�,�FF^�Α�������T,+�D�i����A���]"/���XE0rѴ*�.�V��˙�0�����ڋI����
�0�n XhIFפ%�C�Ea�w����Ŝ�⭵X.�(Ucl��<���D\'������H��w�q���vж�lq(z���[;V̮E
^J��������� �&�b������[Ss�w1tGB�!��d��Ȯf�=�Ը��M3�l[�7%<em��Z�uF̴N����u�J*��9�=��yo��i�D&���Z���.�B�1b&��iѦ�㔉��='�t�Q�<ݘC���8"ec��NNmI���Z��ekx�655��6����>B[8%�4]�+��#n�\��ҩn!fKk
g	�c����F�{�n5�G0��(9�5�ct�$�(��H�<�ߪ�&��!��Ag� 5k��Kۙu(,4��u�B
%��j�����*i6H*VJ��Y���3-2���������X��m��1R"Pp�}��t�)�ݚ�H��%"�Ud�cƛ�V�IA�1�jj�kJƶ	�ɪX�Չ��2�2�H�A��'D�uL�JA�KP�
$�q��u
EF�f<�īRRRQ�I)Z��H)��? B6-��%+�B"��!��X#�nqcv���3J��2≃SIwc��$1[�V�5+�u�z�o7+��O
j�����X˨�igK<��Yj���Я5�Qˇ��_9������Y�z�AR��b�7�zA�L,ٽ�+}��_��O��UVj�:�4�|p�Z�!�?8�i�y�p~ "4��5L�0{�&�B�3T	�5G�gCT���$~��4�f��D\�#�A����^����h"E~#ޚ����`������UvѶ�i���+N6lC	MFIa?���"������ 0��W��=�4$-�� &�P�����H��Q4#C�B�MH�hO��(y,"�� ��En ?��t� �<h",�D�}���d��ǨY�����"������� ,��ʾ5L���4 _���@W��"Nj�3m�||G�1 j� "��>�a�"��B8F|��F�$?�OF+MF���ogڿ.������g�٪�A֩��H�|�5L������@�Y�I��)�Q��ZˠMW�Y0�<io�E��ֱ�%,f���h~[޿ƅ�4O�M�@�� 7>aD)���{?}cN��#���4Oƃ i�4<E�C ?�<˩@~HP[�	 q���5H�D�Z�x��dd5�4! �^"��L|��Tm�(~Ϝ<EEI��4 /��*��� ~�,�g�n��㿼-������&�U2	�V�"�� }�%Y Y�E~#���e���F�"�|D0�"�:БPW?j�=�cuWD��n�f�_00٪��T�p���������a���|�#�Ɉ���M�2Q�r�0���_�,�>44���P� f�G�}��$a�dR"��!�gM" ,�ƪ�lS����ZT����#D�Y��P��45Ay�_.�"�����K�D	�e$���o�>��?�|yq�?E�����S4�G�3@~��/W���]i����7��U�i��CV1�@��P�*�C�C�f�ƃ"��&����F~�V@f�[��h"�y*A����#f�=BϱP��_�GC��5_5A�7�0?�(|Q�5@�����d_!M�D!|
�|��5�XD�4�"	���h(���5H�j��\�Z��AYj��zn@$��G|~�z%�?�߇$�n��{�f���T\a\e��!$GϾ� ؀X�D����D!�*~A��H� �s�*!dW����� ��_I�Y #^!�� �tH�j��`B �E3AL�őD
�~��������h1/h�O���!�h���u[Wt"��ev�S+7f��m�0���4]7ӎk���3�� �V˶�j��7$�e��Qvr��]Zn�xv���x�x�}	���A�"�Q�f�dW�B5@�j�사� qY�@e���!�U�UXG�C�T#DY1�t��A�C⍑A_~��!����]����1K\%��Z��(2*��p����4>������5��B�Eq�M#ZhY����n���r&��W<��W�@!b����|���?�^ћ�fO���qM~T!���T	%d#U�� �D�F�!�El@C�4�!�_�?�b����bC5P��<h24���Ʒ�����J��Ɲ0��v�_�}�X{3���4���~W@,BET	B"�ۆ������B�j� a�ӳ@q����V0���#"�A#�B�V<�4M~?����"�MT#ƙ�Eh|v�i"�W��~�[� �^�Y�yz����E|h���4#@#P��~T:��JȢi\E#U�G��@���B���"���d/ƙ�E4�C#|��D�DR"(�C;���B�N���PG�x�M®`C�Z�o�UC^"�@�ĕ�@��1�4����[hV��R"����ek�3�*�h#�A��E��D��?�����_���@�!�|�@h2"�\�� "+��Y�9E���[��E"+��@dNn���q�qg�DMqF�Ƃ"��^��C�sx�����b� ?C4./�� 0��Ő8֐6 �t�����4 �P$n�3�j�m�#��P�)��P2DĂ(�E�7��G�����P�F�����"�^UdVj���j>��3@�H��	�2>4���"�����^n���<CHF��4��b�P$�xt;_vO>��$��>^2AY���,��a4/��e^5�UH��:���c�Uf�5@�R�j��7�Y�dR4�p�t�Bƀ���!���!�5|�CTʳ�m��w�N�؏��_�z�4�GƯ�0�-m�0�T-/�T(���Z��G�ʡVj��|�V����ib��"�����\��� Y�L��8��g�U@��D�B��|�Y����9��;��
r���>�W�q\u`+e�kֵ�ݙٳ���T��-x���pCyuW�ӦOB���C�	�Ϋ�y�\ �K��+�J��U��j�Kb2��3���w!��6:�z�M���BH����g��C-ܫ��hg�0��гT�����`B͑L��"!����DS��Y��
,��sg�a r]�;A�*�\�P$U񡟵���{���󹾽���~��Vhih!��84b(1�	Ң8A����'),��	�f�M3���B4�"��gñ�?f��X��UL��P$W�|��B %,�9�~Cߊ��ECL�i�������ښ�}���Mi�;�f��8|��@���+@���Q�hB2�"�F�Q5_�$5Ϋ�f��e�_�G���T!���zpъ���d1���"C	3"1C��GۮP�I�����؀r�d�.A�7h����WMIV�rWҾ�3r]߫u
�#�`�a�)�u?�7�t��o9�nŻ~Ȼ\��o�䭔��S�:Y��=��h]B��{�����͓�Y���
%^�ʯ�M@�M�\_��϶x�HCj����d���B!XW'.�HɃ�3lU�g6ߒ�"Ӛ�N�-5L�7�]�󷼳{Y{�d�XAO%ױ=x�ʍ�����g�}��H�K�Vt(�R�7�F�V>�����+�X��.���v����*w1�i��ϳU�xo�EN#�؀Ԑ&�Ѷ�,F�lVQ��+p]uJ�X~��E��_�����u�f��~�P&=�vմkr���#UR��DcaԮ�|#&?IQ�x;&Y��1���.\�yu�+�[��Ro$VI^bʦ�_��0c5���3F���y���3�V�r�F�������j�!���l��������·�.���۟w9���m�C٤Vq�\�*~���(�6�]�����wR����el��+5yj<��Y��ʷe�1,����ߞ�P����U��Ci���[?��~zg�iV�l<�d�8���46��4�j���/7m���A�G�Tp�)�L�p�Z|3�n��E#�zص���^����C��"�Ab��N�L��a����A�ןd���< ������s��IX{jwq���3�j�ѵ��B�PS]��1�^���w�A<�%��_�&�5DU�F]��T^�����d	%���t, ݤ�PY���{V[��~�<�+��F���n�i&�_�D1�w(�2S~I��f���d!zf�ץ�]2�s�ۍ�������,�J�R#��5�ΒP�̹w�=� �`;�l=�o��+%�ۭT���e*�UZuIWgV����pb~pP�Tq�l�K!Z�2f*���[;FwR�UA�Ex\9�)O��:��WY
�@��l��s���tИ�jI�4	�R��¥�qy{;2�a���9"�B|���$�Ƭ�����X�NJSF�׃E����,���of�_��J�֐w�X���:�Zi^�uu�[�#���/�u�jK��vKZ�T�]��\��T�j��躭��"!#��t�O���"G�0���s��k�-���� ���p��C�d�f�-׾���ukϥ>��JǍ�T�}-*r����������*�n�8��`�\2��"�D�l���0�NΥ ��U�l��Ji�u4�΀�^�k���U-�m���9t���N=]*nM��N��oY�E��җ(�{��w�en��xe6HM�┵s�/�hzv�)⟣��y��~vb0���l"���xw�ʘR�����oF���ZqJZ���K��{��7���tf�%�si/� i~;鬺��ɾ�+�_^�p�a�}��w�#�Nyoj]q�9w�t�3G5� �f��d��gV�봊���P6B�ΐ$��U�M�T���o44;$V�uV�*8��c�b�	���q�=�S����S��#I �Ó��/Oȼ�q��D���Ȃ�,��g2D��V�����B"��Q��XW�;>�j���t� ��^S�#̱�w'ƨ�*��&�t�9�h�Y��7��zGt�蠆�;�o~��Q���L�Si�]�W�.G���KmfG��ܡ�o'�F��z}V�����	6[��~���`wP�s5^��l���`���{��["B��9���//�Y�Zq��T/C
�9=�/1����QE��+r.��xj�w�]�UoTY�!d���k�<G1c�H��_Ц�������p͵y<��2fjk���zA#>�;�b]UtT��DwAX%Om��2j�G) �N��L�^�1�Ψ�Nu�0�3"=�
�{[� � l�F��I�iߊ��S`T>��E� ��20]��9йH�����l��w����=.���_z�\$@~{+6�%�a�4obM�w����2eFێ0����0��v��\l)�I�?}�H�ɨTG�!��9<�K�A�藖�YT�5[�X[����b�YO�Ľ�HomI/�b�����T���ԍz;n����I�����mO�(�V;�#W-t��d	9��|��]�7�Q��0CC�	��F���8^b�dV4�ɷ/��=rDq_�G%.�n�~�&�Z��N�%L{
�ź\�%�Ϊ�"�����-]��o��`�_��
PեKKn�.�W}���U���_4GW@pg������F�<���̋(�]��7c�$ʷo��^#�|^V u t�w*I��º��:Sݾ;Y`�"4Zd���S��k��((jh�<�/z����]?q�/������JjJ���zR����QG�^%�K�M����A%�\Ð��id±�7X�lL|vMw{|�(F|�z/���nW$w�P�\%F�-��cE��t��p���7��PnI��~��+&Й��4��QKo��L�Q��dFh����$�Ci���q����`U�85^'}���3�/�-�uN[�P):|*(�{�0N��mܵkT��]׉Ȑ�z��y��l#��Wa=��Lt߃�ln���ˢq��K�'د�jN~&���G]I��SV�۫�~��嬟�!0ƌ�WZ�Rt�H4�?��]��9/gw��`n�%5��U��js��Z�~�*�|�K�M��@�4�,�Ὰ�'�o.`���&1h�&�qࠠ��5������i�E��,4�H ��#��nC �6�e������?�wC���b��_�ݺzl<P�j��HW�k�o�s+c�$z�+ϻG��Mfz���M,�� �`R�`�)iZ;6�ŨQ���
M�2R��ګ4%��i!J[�^.�d� �ļrT���ưZ~[ēQ��6Oؗ���gL�2Rq��6^)���Ժl=�3ѧD�u癮�I
�^ڻ�i�<����_`]
�Q}q����d�j!Q�췙�ZZIlc;��w�_YF�Iك?^*�(��Z��d�+�Q����ϪuE���aθ��]�|QKK�ͷ�o"J���N{�'�:ƪ�9(�G���F[o��A�f��ڊ���{,z�-���)EXZF�*#N��Wȼ����p�;�3Ws35�I�ߜ�b7�4&������jXZ�'bd�]��f�z�����a�ή����������Sj5MP�{��^��vK�S�) Ww��蓶c����5���=�Ա��iw�uM�/6r[^��:��*xk�gg2{�+��6Q�3�y
d �z���ެ��2}LM�^}�+�u�3�_��}�94�N��%�}˽̼]I�S{�|b[��:�ۘ�����tk����溗<G�+�f䩝��Z(O�����Ew�{t�( Q2�#jKC9+S\�<!-v��-v�v~�"�U؄v�e(�ppͧ���xA2�5��BVشQ��$TIj�QyV��/Զ�}�0#rB���\\�|�)���0๮�k�u2�Xr�v���j�Z���t�:��H��z5��P��`���!N<�|z�[�}��H�%3���-�l	��
�[�38�r��F���m4���2�3	y��2��Ŋ�y���a�O+��Z�dY���2��j�Q�͖�5��ܢ�$���7R�5)<�!�i�q4�ϓp�X�?��梬B[�6�fC�����d�u�n�{��Es��-Or�/=�=^��:�$�h�يm*K�f�tt'm�\���h�����������бV]�&k^qOP�3�ͩ3�I��i�֑�X�Oh3�[m�֮er�8�ټ+�m-�O��	�ڤ B���+�X�+�eP#j30i�x�����N��Zz�6l���K��q#`6�1�C��i�Wa�]��7G��2*IA�iej\j�'�'��OFӡ�}!���)H�թ��+Q�	e�^�\�����Y���f���Y�v����>$!�G��U~��B�<
�M/B�(����ƫ��i=�Q�-��ä���0>�2	u8c����t���W(�"A?/�MA��bA����܄]��A����l���G	������TQB��I�U��s�A�R��4[ ���[����@�p�T��� ū�,�J���7���6����_���ǈ���IUTߓr�@�͸�`��{��ws����!.`����m�8�9�T�Ķ�k�1�Hv���e%�ƣ�or��K[���a^<���d��/�+w>�`�R���b �����>��,�H;�ʉ�ʍ���e�y]��@�=�C��w�MB��C|�^P�<�L篳3�� Œ���s2�Iwx�d>�Z�Wc��Y>��
�]�ck�UlZ�D�v�7o=1pߗ�ނ�o=_GB����&����:|��╓�33ԑIa��Zu+2���;���J9?t�g���t�I�y>��p��~����PYs�6&�\�.'�%q5�#{�g䶶���C�)D̓b�
��S?س�W��r7A���R�\��Ǐ��'�(\v�&5�F0�T�D����n��U/ ���?U���=)�LJq2gJ���Ra��*r�rL�o�����^�"���`��JK����Xh)��=�ĕ;�������Ɏ�k_Tr�XRV_e{>�x6�%:�.�ln\�kzP�llTzuw)K�ͨ/Wr5esB����y��L*wy�t��^4��&3���%ή'oGiO�ͩ�z$��nu
��cΑm���;�#�W�Oڵ �|dSR͛2j�4�I,f���Y�5$����܌��̩c`�ג��U\m��*+�4*�6zb�a���3K�yS��Pd#]�b
GR��:]z��W'����0w8�$h5��.��_���j���u�YЬ�K�W�.���$��p	}����՞lC�j|�^��9�l�*{ѓFc��/J�%ңy��h�,4�3'��Ҷ�CAhk����f��_���ے�5����)��yH��F�1��x��,��E
�0EH��q�G�c$�g�:���:�B�@~��ΓW3.uA��ǟ�L-�Q�%D�������mv�2��=&j�ӗ_�׹WF�o׽�*�� <�d�ҕs��
�stJL.'�ԟ�>>{�2��V�{�rg��4�+���Fc4��H���g��N�r�
ZG��M��+7�Z.ç���MB��r.m�!v�U�.�X%y�7d�q�N��V6��)�H��+-�Ft��K�lO����u��5�}6^�|��{;8�kC�'$����p̄�J�s)bH�]��ɡ�^�w������`�r�R�*�wxy��6��)\[d���Y�Ⱦ��%>��R]uUEM$?i椗F�?�`ܖpc�o6f���@����2���\4B�Hug0!L"$�6/�%F�v��NM]Z��ܝ1W���d�ɧQKSc��L���̄a!���-�ݝY²|KF��ruPG�λ|��'f�4U.|v�^f�j`���t4w����	���*X�:t2v�'��t�en��y�P��X�{�S)�hɳ�����x�K�Lj��#��vFH�Ẓ�AOӘBa �on�V��!�X����ڍ��=T�>�W{n��K���k<�w{����j�\1����o�m����/���/nl�9I��9�ijQ��Io�"�%���Z�e^�����O©o0��Ir*�Fb۹(��`��G��;ӭ*����ηr���� /=����V�z/ۆ@�*l��R�R��GR��5=��`�,v�3[lՄvW��h���s�5���
�n�FçqA�ˎA�+�a���_�o��y}毥�V9�VDc�� '
Y�驾ㆪ(�*ʎ`Nu�����]H_#u�#����R=��z���\tO��w��9����Z��@2�jM ��Yk1���xkf��R��	�eN�d��Bz:��$+{r����
b�/M�ZMEr�y�3�cQ����}~�)�A;�XK�Ln�G��*T ��cl����g��a*��g��J�S��r3	l9(�� "F�3�u��g|���B�^o8������x�|&�T4)�X��)�S��v|.L?slE�����@��My-��9(��:GC	���5�U�����e�}�r�q
�l&Kp�♫�3VĀ��V�ĀxWݸ3��!G��d��q=�	�V��`L��� �p�����ǵ�RL7��ηFg��.�m��8"%j��H��`�$z�>���>�]���V��_��d�P�ל,��.Xd
����V�ff���Rx�f��ì��xiܩDDɛak8�ul
���K�W
�{iͿЛ.�ܙZ�ָ�skJ6$���7�Gٴk��N.68�5zGs��K6���T���x���s�~�jlɴ���']���t�[w)��Yy��oZ��T�{f�ozn�(���zJ����O���_*"͈tE�ve*{��f���lnhw�tۇ2����3���P��F��[9�_��o�\j��{`8o�j�H1���{���c�-���T릪�M�`V�J��)襵lѫ�e>ʁ�Z����q���4�o)^
���g�Cvk��5��ݨ:���
��Dg;	��\��R.p�0.���3��ל��ΉB���3[xJ�*i�8�8{@룪jY��77�N�QE�tV��L�g�oN�2�$�[��ӭV,O�W1d͔t�N�ua�pج��Q��ѝǂ����:�wPP�uE�%�Wl�H� R:(b���]8Ą0��`�J���902-��Q�����Ih�ݭ�6�x���>�ߟ����6�:V��uKT��
��⮛<�Y��p���
���m*�7����ͫ���ZSW���Ҽw�Q��Y֧Z�p�t�4oJ����h�Su�&+V9ڵ�̱g�:I�`iE�=b���@0ќ�����em�E��nG,��������Ba��a�n�C4W��<��⽻�s���ʵw.���[��@�H$we@x�\�X��ԫrNҥ�(6Vj�92f�X�V'5�TQ�R��M�adN�u�?�x
P�[Ϣ���C7R�p���`AY3
����kv�5v/�J7�Ѷ�N��G:H�N$�I�&%�΁h/W�=�i�:�ٻ���~8��M)����m7�C�	w���D��+^QxU�8�"�9q����u�|�N��{r�qq��,
h!1m�|�6򁽣�SlՂV�|>#	��Zei�Md��fB�J��fve�"�&�ƈx��6Z���4�	�u�z�,/�	�`�/������?z�j�d��>��*�t�B��R�Vt�;2,�3ؙ���v�@3/��i�����GKB�,�����Q]�n��IH)������|����M��|p��2���;�B�Ȝ�iR�Rb�N�~�{���I(��⹠;y�z۟A.�Q��5�G�k��C���t�gZ[���M���q��3�fL']h�1�b;@ǄJ�-�r�- �g�t��Cħc��k�NԂh� �No����%Vi
%�S�ٴs�Aj?��s�,�yv,�'�a"/��ܭe�wRf�$���9H���Ϸ7��<����}��Dwz��I!��R��/���>���V�;��{ѷ�3>���K��ACY3:*���cZ�������Փ?&�^!��?K&�Bj#PA}dϜ�]�����{���tfI*�)LG�/�Z�l����!/���a@����&�{�*}"��;�EC��3��j��O���`�G�h&�6����M��%�n
�=�>erK���k͵`kˑDy�Z���5J������Χ�W�e4�z�,�yc�G�cd����a��wb�#�m�Б��^zh���̥��O�ʙg��6�'͏�"
��#\��H;��g�x�~P���zP���B�R�����=eo�|e+�C�{y�f>Z7&-^�l`����-~w�Ll�"� o�LZAi.��o�x�@n�T��wjⰾ�驗���Y��E)�߽y��������o-:�$��|����9^�;r�<�]��ϱ
	2����T �G���W��Zu�քN�;��՝7}��5���w���[����kj� 
�5N��,ö���$DQ	�g+��ɭU�+��hѪx.9� s%�5B���t�Hip���ff��y�pц6����ʴ����Ĉ�_�^��)�I) ��0�o�r�^�8]r�qL�@Q&�Zv��b�)j�F:������x�\��mQbk�r^a�\�/��U�n�[��䑢wۧv��ƾշr�W��f�'��PH-������o��60���������P��y9�:�T���ٻ�cؠ}�?@E��9]�����U� TA���:��J�� *|��N�j\�d�uS��T*3�7Ԝ�
'U���n܏��.m��8}���}��g� r��A@n쭺���1N�i:���������:���:�cC�ݵ{*���
���X��u.��3PtJD�S��q�7BW��6�XAN)�+��fZ(��wT�cQSBe��R���
�1U��Q�/x��;�����[��vP�I��e�
��%��q6|����u����&������׃O���I�N)�p���1J�^�$Ψ�鮥{z;o3��4��X����9r���;=�F�؎��Ǎdv��-�Q���)��l�Sˇ~���B�ڴk�J�b8�-�*B���a,8��q���;�7�
h�X��6��XE����싒Y'�f)���qs�QF���&1�V��e9Fo`�m��O�̈́B{�}���}-�X�����]���0�x�DĔG�_\T���q��U���w�fhY����4�*
��U �r��n���X|f�o�N�e�Ŧ]K7���_�B��s�� ��6��vܳ`
ϴwP�,-�6A�tPr�wq���%��뿲��*��A(ef9��(���(a���%x%q�����v���	�n�aQ�0���e�*��d[�m���`Zq�E���f���W`ݙD��82�����W[��?�[Dv���S��9�{I:ۮ7������n���1v/Q%����J� �w��I�u��Y/�y����dά��Hc����@cw_���E�)fe�
���W-���0I�i�=٨_+5����M z�FEf�r�2ۖ�E!�m�E1�M�}&����**u8U���ː'��پ�Si$i&������*��c��ɑ<��
G!dAT��~��,� �E.�gɅ�ٜMb��dTaK�&Ĥ�mȘ�ED���P& ��=�`� h�� K-����DƧ��c#6��4��#�,��ʳF��u�MG0������,�8������Ѽ��s��t!�l	mt�-w�K�{�MwЎ�Oi�L�/3��*R5��u�^oq)m��0kny��΄������1�3f0m����7�i^<������VFa�xK�T�MI��j�=��)�K��L��q3�qڻ�̱������U]f�t���C�B}�\�	9��^&cl���t��*h���(�YS��C�o�Y�Xm褢�`ư����3��4��t��+Uw����x��nːx�h��e�ܧ����ߊ+��8.U���ĽG�6� �1��P��P��S��P�� ���յ�/y�O�X����܈���w����B{��+����(�Vu%��w�rb�������H�t�cI��<[].Ȟ��Kmº�Dղ�(�Qb��\c�� �^�o�"�f�ݓ���̈́<��	qdws��(��"JV�<���q��Q�DY0�p����<J�K�����#��me���U�� ^�Z��֠��a����n{�P	p��JS��^�lǌܽ閵l�4�gd�Έv����MH��ۆR�����U�UUV,p�u�E��q�~�y��*��6O��g37f�˚E��'���8�w1ud8����Ѯ�'�:�n��h'C纡�v:H�C#�*'ٙ"��O�(��<#����	�^p��G-"i�?wZY[�.�]^�����#��"o���n���1뭻p/v�����Y�׳	'r�9I�b[����r�;ُ]��S/ƵjsM�ۖ7���PÈԭ�������)�h�~}�n��	�6���E!U�5Xd��	#H{@�Y\�g}�\�O7�zc�|8jV�&�?
w���ۜ��sy��DT� �M�Z�� �Q4"g�Rq��H�G��fK���Owv���5}���	��C�f�7�܉t<yY���	YLA�LA'm��k��ͥ��fx�%c�˹��>�0�7�/%ey5���l��ص��	��T$5X�t�2�0(H�2r�6��s	�!>��5[�W0aZc�hC`J��?�R��A�
���ӳ<{��:� b6�-^��L��g͟]�*��A�(�o��8]�9��/�׉�L�K���{�wnA囥�-��S���$BE@o�e�Q���Ynڙ���6ES��n�}�{���������z1���7���b"2;�n�f�1-��rV��3��y��� �a�h/��[��]�ն<94Z�F��qٷ�"��:���]{<sŝ#��&o�ƕ]�$,�n�Ӷ++t;��	a��u�
���Z�v���ކ-�no\�\��yF��[��6n�H����::�Q�LO)t�˷ԫ���l�L:p���g�-9�{*`Ƙ�7�_C�҆���ڀ����R/3H��+֮"��5eFǷ8x�7���{I
�7�j��J��Օ6Tl�0L��L��9���ڥ�t�m/Vc���
������Đ�)��J����W5\��-BluEz�;56洋B�t�N#[�=Յ�;�Lx+�=�?x�oR��艓Y�j�VW�$������"��k|/a'�E2N���X���a3�7¦�(U�+����H'�л�[.:o����QN�Em��F�������3��'�+����WO�:�["i	ETdB$����K�T�j;�;�4S���z�M��y,�ҧ���U�������#+�Ǫt�QT^���L-\y��Zk�p]U���0rWԲ���3a���ON�V���>ښh��n}$��	����t��}/
�Q�`8��]\��4���j��6�rlTj_@=�Y�
�P�Iۑ���d��P���9��voc��ό�o��,��h�w.^z�}է�(5���5��#;L���=0g|G]C�*����uN�`EA�ۮ�4��"6��u���;�Ʀ�&*�,�Mশ}��j^,���x���WS§�O��F;yO�~��S^�wL�U7�'ԙ�����p��r`'Ay5Sz�	N�kQ�7As�Ȉ�ʯ#���:]娷�.��a�m�>7fw�Y76v�==��r{�,��	�m���+c��"-�^J�cl�" bqԂ!lJ�s�+[�5�!&��3�[�!L6��R�4�0�o�F+#|c6��ЃJ�*�Tڀ���R�Y	�r��R�9�R��g5<ç	�۱��Lx��v���X��\��d!��#�8ǱM�<����T�������oO=ɲ#7�1>mGEy�����P�+������R�=j��P�詃��xou�c���e���.������T@�\��)�>M4Dg^�~6�ʊ����Y�o��X�k�oZu+�/��%�4=@��ٮ(����	`i	�\iM�t\
�H����eqKe!MߝEj��٬�Og#y·��Lo����!����P����6�,��E���s���a�E{��* [T>vx�<&���W��zfR��o�D�wU
c�svj:&�f	�)du�����=�艏��	�ߤ�6�6�i�X�ʂ;X��J���jD��2��=\��Q��Si��T�*o���3��&��_-�Dz��{vF=�	� ��/�n}3�>s%	X�f�����d��%��T�^���'"��OE��#+�9q��ZT,���`��!��?
���_��B"t�*b�6��Fu���Vl��S�#�x�]��0`�+u�O�-��f.��<�W��q�?ZO�$fJ1���&?lǑ�-AS�_�{��F\꾘##� 硞�z$W_o��",�|.@��c�&����o>�v��9�N����%Y�Ǿ�c��O���tn�z ��^��waε#�g�]b�>*H��>�����<i��Ur=	��Mʈ
���&iy*�#��^c�	h��t/�x�ÿ}��x��
�YVb����(�F�Lr��,o�d����w>"�u��|��o]L����z��)-���ξV�Z���=ٝo�����g~���sāI��m�Y���H���n�8�z_L�ڹ�V�d�y�SVR#tҭ!�������s�)$I`�ƤeC0N����$M:�P�8<ա��o���\�[;����Î�B{ȷ{�뉼��\`��#��'����S�)�&�����;�0ц&1�W�fz�I�1��Њ+M�@	*[t���r<�@�*�C9z9�;�B�"z�2 ���)2=�n��>c� �/�א]�ݫ".���U���p�W&io�4*�
G�� �1�f��L�q<��(#U�֋��ݦ湆k�ܛ��e�e��	��}]{&]�;l����5��A�h"|�ݞ��^����9����-ġ���{��:9�O�"��{��
U��LD�C۩����ĚF1w�V�Ҕ]����@���
5�O��+�uI>�!���ힷ$Y��`$#�r�D�WI��u���/.PӾ��������4�ML,�ĝi�֛k��F�~�Ab�et�7�b�H��H >rw&� j2�usu���kB�\о3�G�&���C�7R���z�i�e���P����Fα4��.�@�(7�^UfR�R�h�מ�u>߷q�S�%��]G`��z�33$Na��q�VZE#m��"��?b��M�ݼ"��p���ˮ�.��)�I%}�ЙP����{�Ƚú��4����C�/�̟jF=�9U]R��»�yct����Ve����<۩�b�H-n�n��tל��k]\�f�翠�J.�p��I��S�ڠ�٧A)"�e`�y�cU6�D�&���V���M/G�����?n�.<�ۯ 젅#y��}��������j ����3=�J^ql��ӥ�'�*-|>�[�{��g�Qm(0E"K�5}䊷8��LŘ��*��r�c���.��R>�쩯7@��ԋ�����t�$�"����:~�,TS����-x���D���ӕ����oqU�:��Nvxt��2�+W�t�9��W��E.xRw��a5���ģR�0��l�I��K�[=�I�_�4Y�KsGF�t\ݝ�I����":N[@T>����Q��������-�i�zT�%�?��-E:I�W�w�^,ҕ�Sn�`L��P��ɋ�m��ԣ��'fa'o��F�\�G}�����E�^D>l}���)z.�l��'=PE߾5��ϛ�KCa�Fs��D4S¾����^��j�i�'v8��	2nl�i� t��P�[P�CH����B�Y[���-MÚ)P���E[K*��L"��
��A!(/v�[�T&8TJ����1���9ϝws'���Ex \LU������7�M�P^�ܗ{&؊��,t{`v�D��f�|S�v���Zp���t��"h�9�d��K���j`��YJ>O�b(�'�{��y��0JW���>�y��rXJ��#b7ڦ��f,i�Z��?�<��&ŴȞn� ���.n����O`	�R�t���{�oo4e��\��e�!��=3!���R�'bu��uy0�9/3Ћ�˗擋"���K}:X�����[V-kX�#��_bQ�b	O&�(�����fޙp�ތ>w�G{�e�U:�@�m`3�s�LxS�S��N��La"�=BUA��i�|��}�Veq�\&�V4���T�1O�R"=[�SD��� ��z�n-���ֹ�����5���%��Ⱦ4���.E��E���ܵ	9��FP0Sd_L�4��E�&63iO�o���4�C���.�R���s',�������Q��rY�}�����j._Eq��{���:3\,^� �r��dLT�y-��ߨo5B���BR#�<�q�.+���S��8��O:�����L1-�Oܺ0�|_���a=ٜ�~�Ψ��CCt��I�&=���~�֟���m�h8�\�Yߣ $Xd�
�ߧG�6n�h��tuF��"5��j����U���8l#ҝ+��s���[j�ᆫԯ$"tO){�dql���yyd��$Vy��k���r�;.�5�"��5�c��il�%��״��F��C���{���<n�3���u��o��f�kzɷ\-�g	e��;e�F݈���ŀ�͓�!�'�7ްcuzon��ߺtș�~E�Wg��[�q����0yo��[8Q��L�qB~��G5���zlR
�κ��2����@�����bt��ڤN��^M�F��p�Q�Z ��"�Jݰ]�M�O�4��ԭ�ۢ��4�b�G*%m��lVVrpV䩪;�,8�eA��OmgmL����[Dn~�eٚ��ԁo�+:+�MN�����{L�(+Ԁ �Y�+naV�����nݎ [B�d��g�vo��N>6�d�Ɗ����9ҍ�'d����BT�8{��f��0Y����j�|"�cu1d&5$��ۮ�Λ]Bn����E�����Y.��d2Ocac/:s��e��M3�`����ϭB��4�İRD$Q�9����_�a9Ό��N%[)�,�6�{<�,Dq&�?^ڴ@.C�)�/p�����&��pnD!���5��t����y����3�A�'n��˩��ƹ ���$}�)�`�s�'�Ĉ��o8±K��9�^i7|��f�T��?H��-O:����c�y��j��QZ\&�^ }^ts ��{�a	�x?g�f���>�]����˫�g���J ��J��I:���L��o��,{�xP�(���P>���^�{��ҫQ�l�[����m�j=Uį����?]곺�\��q4�$nq��dE����&�zj�V��=]�qEz �]�tu��eN�]*;���g��\1�} Օ�6b��{4���-(Fn����Y��ά�24(�\���A7?�q�q`ȑ��!����yͩ����ǀ��J��F�llI����ۙ����|�Mz�wջ��J kQw�Y{2���!{��\��Ԉ/Ǘs�<��x}���g{fA�(���pr�Y]���ݵ��Y/v�����Ą�5���ρ��^��F�2�ȓG#�y�xZ�	�p�O�����M|��5��dfYz ���hBM�L���g��ՐB{��;U��~8]��/Z̫���ȑ�啠��q��1��q���P��<=T>�����h|8ݖ>u�z������U-u\�2�2�*�_�n��ƶ��N�n�<f���[�#�����Du��M��Q�GjS�лY�gNy�#���p�ɊWK\_2T(WJ>�eW=<�+�P��!��L�؁�t�b��<̡] ��^ud�RK����pa�Wa�j�ut�K�&�;��yiN���َʃ;-%�û�Z�"5U���#����:�'�c��!KgX�y�)�f���-d�4���Q�ǚXg:����
��s�`�:�;@H��v�c��Z��6�5����^��r�ppOy��ԹG�i1�.��붻��[��N��w��$�L��QML��y.m>P���#���E�B_���s�����ᣳ�#X(�[o4<�ӥ���A/��NA@���n��Vmk�����7�`�g!��;\�@g9R�α�r+{���iyiR���FU&�V�7���Veyu_8,ם����(֜C�9]؟��9�c2���'z;Tj��,�-[MV�g�Kv�Uc�z�#K�;z��ʆ�>�i'�~��A��Z:Iy;m覂�16�oQ�y��bl\c��%=�z�,�7�Sk��ԯj��Ns"��X�˝��s�y�d}�~�e�}Fۂ�p�n22��nܳ
�@�쁍b�/�i�pS3� 6J�2�8)�����-��n,W��y������d���Wi�P�XP-^d�P�4{�]��7��i��i�e.d�s�S�γk�R�����)�f��oƠ RHI+X�6�I�          v�^0y�%���û;�t�����w��xo7��ˆ�?{�tu2`�$]p�Ѵ1<Q�2��.�&en!�1���9�~��X	=�Cv �����D b�{@�%^©�:�c����0�H+R����V&�-t9O�O7^s�/��ӭX[n��ߢ�nH
�bǙm'y�]4]ŖM�
lO{!��/;/t�!$�0�l��|wu��NI�!)lCj��&BSh����a7z�r�=�7)F��N9k�qn�ѫj��%�x1D���3b��"�{�+����1�u�.i]��h�'LP|�3��,JQ�Z��R��ϓ�Qk
�@�i%F��fem�/Ru�`o$4�K-mM7D�AkoXZ��!��$f0A.3'`L`c2��*���D.^�̱j��P2�Z�]hl���ʤ��^H���I=�@eļF��6�Ǌ9R�oz���"�YF!�G���Ƚ5w�8?�=#�Zc5�:���;۶ҷ$�&ZES�U�X�
��&;;��f2�� m�F^t��uzo�1���lL�]�Q��3��:��F:v\q��o+),��m*�!ӑ��p(f�� C��h�����2�+��P�@��HT/q	��V��a�D&8��3wv�4�&v�ƖGBF�|�y*D��51n܀��=�� ���0\������p�MV���:
�v�QN!Ae'���)��H�&#��&�5���&���o�7��L[=�w �4M0����',H�k����ҡ�d�=%O�ai�6C2M�၀@ӊ�'�K�[f���2 ���+1$�7*ڳ$H��I�ڽ*�FFԚ[,+��wf7�j.��b�DME��e��t��bˆ!8-�(�0��iv,^$:+5���Nf̒�5	z�:������j�a����;��o�:�5�������������j��A2��sUy�f������-$�S���Z�Vz��JpNj�Pe+�Jp�5�s;;�v���#���d�̼E�K?~�+��-�PA�F��?p���~�8��L��L%�1��c˙`��j��J�s��{%7���J�J�3��qb��r��j4���6��S]�OH�s*3}n�	�pKRN�q"��*������f�3v�Ǐk@7�9�b:dr^�Ϩ�r{��s%�`�F M���fo[p�u��xnX����Tr>�a(>b�(��q��,�]�����#K�+p;�ؔ㺠�mC�ik�������,�g�
{�{5���_�0��F�$e�ŭ�yz��v+w��}����9ƛѺ�� 9V?��AD�|�ic# B�՛SX���P�:�B-�Y!7�ўw�x8)ެ�����*�+�ْRp�,U����R��|�UpgX��wӁ��;��������5�g�=��)oF�u�L�q����J�e�/�cp�����%ͦ��P�m����q�����Tn���D�/��
�:����[��7a�zh|t�'<9�}rFs[������Q����~�<��;�\��H��%���Ht�o2r�*-��P�}�\յ<Rco+$���ߎ�TMf��8�2�E?~�G-|����L��Ɯ�|m-U5& ���$���hD�%��ȳ��i:��ߵ�P��o�ﻦ}��z=��ݙe��0	�<��j��� {3D�e�����O���Cz����C��Hױ�.iv����`��gM�!���X�y#�e�X���e>n���]����8%t���
&Ú�R��L3��?{I^~�5�ث<:��s�hԠ�b�c��|^�(��}����
�]rU0I����YhO����svb���i�Wz�����C*,��.�oD?lC
���WA�ϞI��R7�2��rp��M��o�zU����f�<�����9�ɘ��=��ϕ�^F�XU�/c��3�w���J ����w�6>3�ME����+({'�zq~��)�������6��O�����?N����Uy�YFXs�4�P��W<�8���{���
[�r�����ۑ�ԪJ�x�������<�t��Ǜ`��u�L[�wwdA�gr��+*D��lYzU���U=㦂\�K������x���.�6��ϐ���~P�}/U 3#.n������T�aM`�"{7M�pq(=I���Uu9�V��}���'kg��hA��%�M�Iw* �۹r�և��\b�������C�80+T�7mB���簗������۷8��F/�9b0�U�� �HAj_	��p#�Qu�M��l�0��sݓx�̃`�N����5Rڪb����rRT}p3��`�&�H�槅��c۫�S�ݜ�&@�@e���P��/6�]�6�c�LUD�ㆀ��B��0�<�`�ⵝ���z|�X��ξ73�5D�4U��_<Q�,���V��|+�μѹp��k�d(�i�Q�7��#�>�[�m������vO֞���7����8��]c[[d�U�+X�i�)��wD:�5���ǨQ_�l�ͷ)3e]�ݓ&3���Jv3��U�vN�&kV+��֊r[����xƿS��`
��E�5����63�@�Ucsa%�!B�I�M܄�Z���"P�e����n�֊�=37Ißv�0�d��yJ�f��k�3|5�'jt�+�=Ko*n�g�\F�8��]ƹ�z�K�StT��@���U�k�}8�j�e��b�أ���;�z
t���V�}U��V��^q�Kۉ�bBI01;�u<E5��+�ي->�X��xYf��Eŋ�}�}ܨ�s�/E�t{Qح�ۍ~3���$���y*<Ўŷ^m�������2sd�T���Fr��\)`��Nl�_v�a0�Jbd%*���B8V*�߰�|�s��eJ�}���|�dv*D�
&�������
tT04"���X���c���&?��2������&���1��3x�nr⡨����n��^��,A˗���г��<�e-v�E��_�GrQ�ss�Y����='��:�q���pާ��K���h�/ksX�D�UUL����㤗m�lnB5	�6�y�9�KA��	��}����:��9�����ݔ[A�[f���ΙD�a��i��A���O��]�空�9Z�2��/�D�׉�gK�V�=�H���#w��&�_|Ά�̅�q�}�(���EAV�4��6ʍ��݋ap��k��T�߾�;	�����	X�~;l�%�]Y
�=�T�gst὾�q��
��[�>)Sn�	)��O�r�^.+2R��h\.̥٤m�$�I�s2����aE�PNA8a�Ɣ����j��k�V��=Bۘ�<w�ٚm`D�`J�cu��s(jǍ45(������Cc�#������/hּC�F*��ǖ�Eɭn�F����R�L�\���y ��t��14���$��?)�nu�F�J7����{��h�q����}~��G��ȕ��R>\���V�~=���P�����d�fo�'%��h�&X�W�gtH��������~��7���ꜛ�0$�"A�rr��]�,A�w�`^��{y�'N�
�0�:�$um�}[��o=��C���^���b,�(~�.+��چ�UQ G�,Ԯ�;8������1z/�u���	��8�7�����,R�4Ң	�&�I��ja-�Y
�#vw��M�����f�y��܄t.�Y�dؔp�s��j0Vc��v��'32���tW-�Ȩi���>��h�}��J�o�C����X�1������}�ɸ�m��E�C�k�b֩���^
gT v_I��w�82_�ԖS���(U����迳D�X�¶hbV=����F��վ�z��M�:\r��&���_�{ ¸08Ou�_{e��
=Y�Yq�k^��ђ�3���}��b>��8a)��[ҳ����ӽ=kz�b�9�4R���W�52� dE��{pKB�=��b�S��8Z���yAl	q"�����u���t�ZB셾n�u��q�&#�X����	ln�O�TtM {��1$�3�0|�'iL@L�s+.c%y��C�M���!��f �*�
Gj��ў�4�s��y9ň����sP�M� z��0ͧmWQ�C���pX��I/y�Ὦa�5T�l;���o8�2YN�;�j��B�l4R��#���j��>����j�H��Em!�뇗_(Z�F�XC�4eߖh��pG����+/�Jm�)r7s'�4�)�(i�0�h�c� 
�u�[eU	��ݿ������td��\ۡ�8���9T��?wc��a�0J�q�h5��Y+U�߱}Q: �O����F.��N��3=�̑��jje��I�/^�Z&�Pon_P;�J+Wy�-s�tP(n��2�Ol���X�ƅ����}Oύ
,��x׼���pLͽ�Ǻ]{#���Fɗ����| ��\��v~�x��N5�B����Y�A����G�	c�dViR�g�h���1��e�e�?]�Kr=��t\�y{����$Z⯳eT��6��7V��,.��=d�s9�4��Η���E*d�	�Dإ�[{q(���4�Lk�ni�� =�"'�����2;��AZ�M?<�l�5QUj���v3<Q[�h�W]�⫝>�p���dOk��
6��@���?\.��A��H�-Qvv$�#��	��2��(l�l�|��1�D�4��kDnm�p}0O�a�Y�$��j�����U�}���~�S�;P����������F��)��փ�Kblk��'�	��0�w�b+�S�Z)����ޒ>�Z�{�8�(�SE�Ț�mM�n�#o����7��+��Y�\:q@*��6���z�ؑr��V��Ch�%F4��u����9���^����Y��D1�؈η.Н���Y9 ��+/��0�9 �)gH���r�(ft�Vn�g{:��u�,��w�x�ޓ�#�0��^L���{׾0NrX���1XZ#��T���z;J1ܷ�]g�������^ʁˈ^յ=�=��1�y(�XH­�<v�N�}��7>��Z���f3�ں�}��;�:M�>�c.��������o�y@g�]���۳�P.h�?T�#�G3�\kа+�k|lQ�,g[M^z�`�b�M��j�tP���\t.�4Ҍ/.Y�^S��ǡ0�d�F��O/���|ʥ9�q6SܱWOWl�x�U�I8b8,J�6�2�k��������@�Y�Z�A�͝��kf�4�ɻ�Br�瓵P��қ�Iڛ��!8<Qd�E!uf�C#�r���mV�)x����=4���H���@T��b @��!T�6=�~�zL{���P�X2S��3Gt��I�F>�f�k��3��NRBTk#c�
aU�V�����K/�e����5�ߺxQ%]�/L�#��g�-t�d̮�5���D�#f����6~��Q��!�g�2 b���p�U�1Ԙ���FpJ�j���x��Z��^�^�f�j�f�
����B�v-������x�n
~�����%��as۩Jx����W�_�E�[�YB��4�J/P	}�tr5�es≅�\T���nPM9�*����N4�(B��p�k���~��<4��xح1J��36N��e/cwnݘ��$�wutJ[��3Y0>}!]x9��ըZj�� l��ۣ;�R/�7�Fj\���˻S���"��Pٴ1�7V�|��/��k���.W��e��P��GG��� �`Y�V� q��k(ײ��;�MAG�=5ky��P���<��sv�T��{�r%��_F�9����GC�WC��	?�ݦ$|rT������3����C�R�-�P��vZ�ܧ½ǌ��o8�A57�mk�#��3��z�Z��玲t���`]�W"9�P�s���`��:���jm�}养��]a�p��̫B�>yy�7e��w������۩�pٱ�ڗ��#��$'��ϩ毽�򫑶u�ަO0���n7{�0�1���`���LM����M��i� ŷ�@��m�C>���� -y����ae�Rδ9r���xI1%|a�]��ᆹڡ^E!G��@}�V������U���|l�a�~���H��$��,���?u��Qc^���D��?��	�K1|���̘R''Z7+G��Θb��f�;��̜����k��k�g�/(qfO�!��"�Z����fQ�_����oI�#<���.qIg��EN��JN���f4�`��=�~2U3�Ë���]�3�w�qj���,�)�O�y���Z���'�L��S��"K��n;��9�����Y�5�IU�`#
���Q��Od��K�@�<�(��}��s��m%=Z�h�Ч*�7:��,�Yn���|%N���zsZھ�����؅�i��u*;������Mz��&��+���&�$4���G$���2��ɛ�6��U��	1���[�n[m0T�nb6۠O�;�����顄P$��˰�l�	�q��S1��>8��Dh4��$h1����ͽ�wc/e�3��E�Zl~X���Yj��z�zK�G0�睭p��Z����L͋0-u�1�U6���91O��_e���(1Ʋ��Ũu}M����Ш+}@qJ!A���bh����턶W���Ӧ�J=���7�e����ro���u�b$R��P���s9-y���jB�A9�8����5��9̴9��'�Ip����b��t�o�݋ӱ���U@G�~�U���K�ʚ�p�wp!���4@i#�˜щ���jzMg�;�Z�c��#�8I(���&-������k�v	"@[Qo~�|�@Ow{�grk�7Ir��z�b$��SĹBB����Q�ح����p��0|���B%��q�)��?)��/%�J��tY��E^�(�G�]� �܉����A�����Cp��(7p�7i�]���
�����j�.xQUTȯ@���s�y����5ȅ����M	�R��u����pE�J��٩�;���x�n�:Ι��G�����̴nl�	5����=n:��*�0{��ׂ6�1��90�o�+��O�����P�Yk~y6k�욹�����\���Zrr:7F��{T5��pI���N�E�hqq;¾�߀n��;��Bm��U��� �>�u�=[����z4q"�Eo��iGM+-\g9(��ƙ���G{���d�1��c����}�K�<��T#O������[]k�ՠ�A��.;^�xE�B��t�ԓy_���kUf��1�.�R�;��`V�����w���e����:e.�˫�.
g#]��<;/����q�Ԕ�[.f^=�	����b��q��|���EE^6�S.��{�j���A� ���ңv;�sUs�8s<*�P�����=����$����v��� �ZJR$�:]˩!E6�,8���(& h���s��,�����98����+_4�J�%=k�-I �Q�}��B�L���D��7~=o����Y�����ɧ��i��)����^�3�<%o����Em�U�Tp�I�>''.��t	M�%t=s�F��Z>�N��y'��jC�m_�M��m�Y4��^;��O�ڒ�Qܣ�<��2�3|:>+׶;����#LF&����Ŵ�#�'/W�ӎ�kyzc�J�(Y�y�T�����1-`r�c)�_�{K%��~���ͺ���ϟUE�ˮ���>�uV@�퍘z�|��KLe�2��oG�e���f����2��P����PIh�<�{ܽg�-��x�2s�]����������&�])V�.�8��u�w��W�X��vU�ߚ�ѽ�]�7�iNfW���9L�C[ �.1]޾�f
�e����L�`1�gH��8�D�?�2^y�gbřvDq;����r�=X\�(Dt;N�9�n�g���jjP�b�DH������0�O���:��3'���}��UV�����8�[Dq*��HT�'k_׍��{�� �����>!z�Z����U�B�>�x`;��nY�q�;��a�J	⮒*�jH{�{%؜�1�I;��� |�ܙ$��8�I��2֮|�Z�v_A��ޅ���ӝ���|���|j�.��4oI���
'�	�yg�8ӏ&�6������W7n��%4w��_�`�9�<j
�<�Ef��4�bhMU{���Q�j�/g΁��eMC@L�7��0���H�ɗ�[��X���~>�X��p��%+��"ir\�֊�L{Lx!��(�ڑ税����ە���NN���V6adq1_�C�s,nd73���]��8�tV���װ,Ui2�1�u�=]����e�}G�6�����7uW-�vk&5)�)Q�O�����BQm���Yv�m�>Gk��j��X��u<V��W�׊$ry�@��ь:x>������;��lEm�F���^v�dd4ngZ5�ޙ���H����߇���LT�J���
��GlaU2X�v2+*�����$�̏嵙��U+���^�I{.��@�_���w
�e�C2�)�0
��!ߓ|s�N� 0uv%4��E����TI�������P(�0�������s-����v��f鳬Ƹ�'�i
�o�9hT��z�+j��"B��N�}��*7�^�=	QD��VE8��h��]�����������.�#s�r��9;�ɫ��Z#�N��j�v�G$�dgV�x��͢��1v�4��.��np�إꖩ.���tA���J��u�ԍ.B<V�u�.fWj���v��+S���M�/��;h�=��N�ڗ]��xtK�,fe�A�M�zNt��A���dtuz�b�*�͠��q澷��8��R����8�v�.���5g��d���l��yS��7�r�o�J��z�wx����XX�I~���Y�*��O-]G;B�dp�eLU'e���֯�uÁ�]�L��\��q痥ʑ��h��p�I#�s_�_R��r��^�3K�By�G^ܭ5�R*��ZNq�������7Y5�rۧL�-���NV�f��Zb�����#nbW�E�Y�A�R錐��ðI��aiw����9���3��:�P�$�R�^X��þ�<.��2],oW�I��E�:��è9�q:%�*o*Ux�)�����V�+5�n�\o���e��@�]�4�ʡ���YxS��V(�.�J��^d���U���J�7�Ne��Ɓ�%X�����͠T���=<ܳ$V�+S�����+��{E��kJ�j�)��:��ʘ�Wp��Qu�%Q�� |��U�˨kw0�v8�˾೶W	�zڟ�v%�y U���:[����vgU��}St{k�U����CH����n���www*�z⣫;k\�n��7z��iD��C[����ww�{�F^Y��\�K)�#��#D�o:��+7�쓢��PVV'����jk�����<0��@F��*.;i�s4�ۭܖ�SMH0��l��%�u��ʞ����M7�[���^l_#�GP�RwOZWi]�U��Z�d����G�YV��l�ء��F� R\y���}#5��u����Z��M`�y"�^Q�b����VSdF2J�6uh�v�:ɾruN�S5^7�ȶg�o^V�^,"]=�)dݩs\��	שل=X���Ʌ�STpM�CvD��+��J�I��D��3)�s���o70�*ѽ�m3 Z��=+��iy���&�7�ߧ�鞡^(ݧ��Q?��O(���T���U2|�3m,_�Վo�F0Sn�c���p��������
�ew'��U��|�VD�~�I1K�[ʴ�M�Uq͋�	ܹʉ;ĈpvE������[���쁫\n�s)�ȹ���Ϛ0��60`��R]{=>ȹ=G�]H���s�
�S��x?W���2:���+T=�k�N{�����-�a�x����[*8��)�/:�ٻ�hdn;;}�z\��z�}qC�_��>W�8�,m�H��r�F���j��T"Q���VBf�.�3JZC��U�t��[5Ǿ�[D�ǙK�F����IJ��N �Ȕ�u���G�/$Y��>�
I��N���7~?Z�Ll>�C�ӭCN����7@H�&��+��"�	��}��z᜺���tqS��D���'1X�&���82�CСy�Mǭ�?��轊
^!^u�%��̆�6:�]�qʢ�Gcbӡ���}g�@�ٷ��O4�,���2F�[�3�:�J6�v��bii�n,���O�/���'��0�ٷ�Ն�M��l��XW�"d��)ֈ�*�]A�ЁT�i��� �R"�I��Ի�	;q��2�m��p��ЭlvW\O.*q��,P,�GF�9Oai=��'�K*�ߢ�2���U5��QF��4�0qڭ��"�y�ű�=�\٬B��7[Vڧ�͛��1:�I�+�&�1TzlZ��wܙ�ƔCL�V՘�&(��X����
�jR�ڣ�ʥXf�Zs����%Kٵ�n)ʦ8��������u��6>��l�I�v}�M]P{7+����S��n�Gtd-ɱ����)_<���h�~�4g�
�z�梾�y�\]��G�]��W�7T��On������L���|�,:�^�+��/6��Q��;� ���{�:�kc��gTc�=iivŎ�:?�J9�s�J�i R\�v��j�[�������[��96�0��v^:�=��I���7�`�*\;ct��:P{�^!�1f��5�wﶞ�SBi87=�&A_��w��q���j,�#`Ft[�AӢN����p��������q���
�{Q'ȵ�_�+j�6*��Z0�6���5�x��s�v���K?H��V��&x����S�z��5�n�[*e^9�T*<�޸�����o���ME�����x辳�;�J_ʺl��F�r��##5�9�����b�Ӿ�z
�#*�zƱ�ML^ǶFюT���J�nz\��B&��2�{��TkT���b�z&&�n@մau^�TM�-Lq�.�B�������S̗��6��ĥ���y�f�9��^2��kb��q?�h�:�
�ɒ�J����_3���,_Xʙ3�[r�%ER���A�Y.�lTә����z5�E����,��L��4	5b{�tǭnd��<������mT�l�)J<h�Wc.�w����o�����B曀f'��黍��.w��ٵ�S;�br��D��V��(�t�s	��6�Ot�s}HT��k��^�W��~�'��/�xL]��`}�k-CFU��C�Wi��j��L]�Vvvיt��D��uΓ�4��W��o��ｅVs�ئ�r�+��ޞSŜφVn�����EJ�/�#�Dm�1�=��jTQ�4�����s�95��SBfVi������}2�|���q�mȇ�V�|r�E��h���_��hU w���ڈWV�g,-����T��q�#{O��L(����f.�/�&wb���حÕ~�(�b����u��ń��d.�1:�fY�>�ͱV�R��AQ�X^�P��t."���r-���L�l�级}���Ə�h�L	�\d�mL
�rS���� (��6��$��H��e�R�?K#}o��v=��3����N�Q��Ū���������nn%���C�a���b�v���*���4�.ɼsF-�g����ĆU���|��Է��WLfV�ל�DپF�W���ZӴ�u�ZU{;�T���IdI��V1~�~���iNa�x��������ڙA.ӗpp��٣2iQ�Rł��#݀�¼�ܱ��>��]������/��)����g�שE���V�!B��B����;��<HTl���Q|�#�����c�7�����S:���Z	�tz�܏�Ҧ�Oo���#������[���IjA�}ޡu��������V�Y���Indz&l��FȮhCH>K{(s�]�7��v�.;��C(%�Bs�_��*�穩HHt������ۊ��cl�`}\yX���>
5y�xkȥ5��;�w.\R8'�TW��������z������TU@�ކ�
f�c}�+MQ�Qf&6{��K�2Gh�b��&8��J%�r2�țt����c4l:{�0wǶ��H��b_������7�1���6��/��Wq��7��cf�$zoT'�.�4T-݀P�0�фg�G8ʼ�:2͟���?�T��#]�
пr�&�ǉ���ֽ+��������}�\�Au�vz}�����.��� 4�*c��ٿ&x��W��k�S!t��|���ꅓqG��T����p�lŚD�r���=��D=�n��n�3PڰK�MW��y�N�CxK%��b>����ۼ�u��֦����p��Ӗ��))����9�i	�͙��=B�ǩ�������������*Z�~�:G�)b=�gnvOD�~�э��+R��&2�x�GN�sf+�Q.LQ�=\y�qb���;Jb�1��ћ�u���SWݷ{h.���.���]�^;jX���ө�~���.8_�vw-���1�v�̂�F:F߅��a(c��.|м������ȳ�x�o.�Ύ1g��!�t��`̜4>̠U�|?@�\�EͫN8)_�:�7��������i"[�r�)B�:`?�#~���^|���C? ����B"�Z��	�����X�����n�p�0!��/���x����` � �{��"�Ϧhө�R��˽
z��U��t�`�\�S��K�2nxe�&zz����jiZA-^�0��W�g_��0*��ڴ�tFB����|�~�[6�z���v;5c������ឳ��߀��I�J���=b8�E;�h��(���1Y}����h�#�����^��7�g�?f:ff�;�o�g{�~�(ï���'RX<3�������D�S{5��t�C��,��M?�4��ٌ^^�E{J�=�u��*�	���s��=�T�M���� p��ob�[�a����"n?�CCR�w"x¬a>���un�u
��"773&�� �7�6�C�j�g���O[6�f8��m*B�ښ��X�k�r�n5��.�vn�\�����v���嘻H�e��;��X�	|y2A$��Q���(�@^P�F�vx��ͫE����ƴVA��\	�Θ�Uwjj�.��y��ѝu�hԢT��Q����:4(�)BW��s�9g�z�7�u1{��KZ�.�,��MߓZ�o.^�:�S�>
����J�nAk���j�`��`���yĴR��+��Y�%��}͋��(���MA�p���ךㇱ�Z�r�Ё���ZJ�X~��@�>�2��C͈�!S��V�`�����|qR)諮�:^T�>���g�>77>�3�b�3H���!���Ͻ'��"V�7'=�r����\�c��1I���[G�IYCrL�iz��v���U1�(�9���\j�0`��3��-�4`�=b�>�n���ft�m��؏�cn�A�-XiVoʾs��p�7uS�ڑ���*<�UɅ��1+}��X�d����1g�2����F�K����������=����	�ݧߕ ;ݾ��,(\���DG�y�V�V�m���w��&9{�&^��fx��=��R;����Һ����sbTo�{�J���DN�Y�b�:&yw�m��,�^��\�N%�9T�K5����{VR�c��w����^�s�n Q��o)f�3	���ʃ�ʾ}3^�x䥘u����P<޺��u"�4��{F�l��B��O�'��OM*Z�|j)S�>���Si/{E����w=��|Y�7
n�zuy_���~�J�����2�O
���B͖�@&���P���{6]�5T{n�7���m}>��ɻ7w|������6~��"N��_���������
ֶ�����4{ý�uݪ�.�Y�g�lv2���fغ͑�Z~���1sa�;ϐ��}7�^J+�U�c�)��{�u�f|3�K�Y�E��K��=���e�S�����M����CVC9�����=�|Ҧeε�J�a`X����\p�ޟF�V ��2��8}jL�iT�2ꈳMv��� m��*�mQ��=�힫��U+����1J=�/C��:���ŭ��*/*�7��!f�]�|�[�P^�e�q���t������2c� N@Pv���|x��'ezC@�5��l���T�*�t%�XY�����5����K�Mj��0!Z�1�K�;��]���"������U����;�{Ӷ��� ��J��D�����q/lt߽�3��޿|��5���%�ژ�����]��+1�h�Ja�O 7�f5+m�@����i�J��Ǻ�W-X�
����Æ�>�e*^ne>6��%%۶w�K;�nF�	�:�G�Z�}�d�V+m2DgK� sM��2���ñ���~R�7�{޺���`M�׎����<��oH�r�k�|�]��W���5W�w������T��뙽`F�߆��S��SdF���Z%���]I�0����jj�����%9td>��O/�דsރ4��z6��qy{�9��ڨb}~�ͅ��$�2]���'ػS�]H}�����d_|�T�}���8��Q�4u�tcjΕɸr(c��a�H�s��B��o�鋦r}�&�6)H���K��:�qX��n�0�4,�ꋣ�Y�m�f@��i�ٓz��V����w���9��X�WoXRj�
ys��*������9��~��<S�+5{#i���(<<�+��×Q�=]q��э1�ȥ�tq�[^9@L,K��`�0�p����od�c���uͼ��6�V���{�3a���O�rO٭*���.n⟰7s?m�����`ҫ_ަ�����o�5�!n|T�:C��nz�A��j���26RK:�a�ap�#�u�'#��{oZg��Ӧt\]��MƤ�l��2�����T�Z]c2*�"�ɺB6[���ҝ�+���i�z��`���n�t*Ѩ������+�an�n�*rz䔨:���9�o)��,�u�57�wF`�.��rZ.����S�>�b�Z��p뎎/þ9�sѪ������]�O����[՗��j��R:/ܺzs�<�-	t�	]�R�kz�.��i���C�5�?j�Sxk\��j�s��ۅ�����R),���Sa����~?
vCo����qU��B���8����i���!m��C�̜���fqm��/��jc����'�9fܠ��������9�۱�ު��~��2�ʜ�A��tk��^���"�M�CD�\spl�$;�qHb<B���������%��#����p*W������K.]]-2�/7*�}����E�k�43᭞X��~��Wq5��+	�R�y�;�����]�燯�(��U����{nZ�ȑ�d���ݜzJ-Od�k�m���<�r�I�TKs0*׺��U���{��љMz|�7��3
H~=�#�ɾ6�f���y7}�}ꇘy��wr�QՁ��+�sU5���>C/�L^@�P@�(����ufrH�0a�	����Mwۤ�AI��5���������xP�C�at��ե��XMu�Z��a��2r�V��INJ���6�Y���ʺ�~ �oUa���'�H��LC�8���'\��O��X��ϯ�J��z��lCF����X�,b�Yn-��	��IHZZ�xZ��v�����Tߺ!�ə9�,���<���",�%�@z�e��1<*��[���cnͥN8,r�Ю8g����}h��r{}���������ç⤥ڜ^Q�!k�t��ksr��
��#��2�t�뮧��1{�EL�uJ�����#��?$�w?8U���@'w�Pc�:cZV�ԼM������L����;��;�����6��������6��^I�RwGO5�h^��6�:�]aP����j��H�(5`&��j��4 Fsy���B���l��A�T�G]�˗��ڗ�}���}:Ȇ<1�����^���IlO������"(;84:��F�cw=�P=�$��^=��Ժ8��o`�_�t��\h��ۼ����m��7-㫛7�gTb�3�y}�����7�͋�l�i߳3zߏ@+�_nߌc��}�^r���=F�g��������K�c�ƫ]�/h�z��A���wu��)���UU�}�	��Y=�\x�eGK��C��=�$�T�(=t�=�QY�&.e�xӞ���>�S)��mev�琼��b�8@������{���:	^�3�a��n�����DY�QS����Qwu�0�Ф�~�y�6VֈıQ}�]x�22ġ�.�s;MTB,�e�2�
l��H��wF���{*�'m�Q^�p�x����b��k�I�u���^�΂������p�u�,kPq�wM�5����P*�e1Dp�j�,�%j�ЃU
�y�|r�E�*P"F�䏋�]���^c�+�����/���6����iV�/�E�qL&�W�Ȃ���}Zʥ�]ث���{"	�sү��e�܇�k���|�N�3�l�����t��=u���W�&:����<ד:̺G+�b�y4�S��=ʮ��<�zf��'U���C\�wⱬÓ��eڼ���WL���޿�EJ�԰���	�D�M+;W��nf��d�r�w::��+&i�>�}1�fFw�Ь��1��8�5%^R���q��F�K5��"�2��Ϛ�Z�q��܉褛��@�X�u���:R��S�u�,�����k�
ѫ�򍀯I��x2+?��u�;Xپu|�3/E�{/^�,̧����vy}����VC��B�xP8ke�Hj�/wW{�*�1�&�\�����6N%�,�;w�m%y[M����Um�Ң�c2�Xj�(zH�w��[^�V�+�U:9w�++ ����C����'9�7l+�+���*qm�{�}!�ɘx�8�v^a9���rL8�t� v*��1��]ڽ
m�FD,;����Zx����|�Fy�z�7-
���K��<Y9s�t]niFUn�T��;���k7�l� {��<D�b⁰           �ݾ�9�̤�e<���$����;v9v�ɕ��;�:�"�' 
��R��L%̒�j1��A��2][�t��;o$��2,��AV��J�b�l;��I�H"�+L�H������ڣU�Nm���H͸2��}�Z��8� ָ��1?l��_�� ��(��y��h㻆�b(��.�e�Ux��Ι|�Â?DE�b�e��ЗD�M\mظ�B !DNģ*�㋍�8@�ũ�c�Pl"�BI$|d�����\�'�Ar�r�]�N2����p�C������[v!�E�\�UܞZ�����T+8H�DGv{s[�/&q�JX��۹�y�c65�v�^�j�*�(�u7PY�-�h!]FT�N�+�8�v�N$�?��B�Ĭ�/1_���Ў�Y�m���&����`(��e�4�K�˂Ֆ)��@����M�����޷DFRG��26�
��-	�9i���Y��ƀ�8��6�͍�Nfa��]����	U�@J�h@ã@u�n�^�.�e�(A��W�ե�@�˺6b��a1�aP���u6u�a��PV���b���闙�rǒ�X�o��#j�ێۄy�u,s��ʟ� �O�c�de��$�SPh�.@jNȴ>�� \hZ��G���>����P�n�M���nc��b�H������ ��gt�&��@�M� :��>{�V%������Ɯ�ֲ��1X����dEm�6�Փ��b$�#D�y�V���='v�nPAq�-��G�Ŷ�,��K�2�!�$0�XD�4BC�m��Y,3����N����E�FV2�*��X��hQe�U�!����2��g2`�3,��m�nڥ|ˈ� ��D��J��gK�,�P��q�&z6	��l���q�3����+f���9b�DD!�I�*�!9���pN6	
�a9�A�Mgb��Ki��L���{lڭ��4��vjDn!8�QI��p�՛��JM�X�"eu�آ��N,�UD^J�b����������#0���^d�%L%�ݳS4��'ؼ:�j�&2�՗�|�H�&"��
Euf�VZ0	)!<�]D�i�iǝ�^lMz�~���Q�񫦺���U����v�Uki٫g)խ���� Ǧg#4Nω�j2��v��aD�z^x������ҟMW�~�*�I[�wx���'5���D�JT^v�3�h���N�=CIΗ`�د͉5'�XG��]؞�^����i,��c��oww�F�dbDk�Ö�E�u!��%�z�G�[�H;oM�O�UG�Ǹ6�'!�B�~W˝�i�D��E�T��۔���x��Q]ĭ`���M�7�9��-�ȎKw�#5��!ǃ�%KС'�ˮp.��H��}:��bV>�����K��s�0�:�l�T˚��;�B�a���Ǿ�����!{a��7srS���h9��.����w���ْQ�V[־���ǁ$q�E���]���j��p�H@�a��a�j����r����Ԗ�>[����/ְ@)^��%V�紮7Q���j��+j�+�a��n���=p(������x�YX���s:���rL�.�ӻ_��=4^��Ǩ�Z���;yIEG\�I���Te�g�Rr���Sڣ�4���.�fz	���
qP�=X:��̔θ�w�F,��v7����hmH���%D�>�A���`UL��~�{��}[h�����ᇞ��#{M�����*k��i��f��������Ϡ��מ�V���#6�r��fZ0���ڵbU�t��z�1��9�li��0]��`\��w�Q���u���5QCf��bq�J�㲃���y���d;�Ip�=S�wi7�����|�y�:nA�1�Ҿ�m+�8�.<�*����^�v8H��;Eg�l#�o�J�_Hv�hfY׷d�|��W�$�}p���9�h�����
)5��Nu�3r�p��|��7����pH�����V�#m0��Z�gK�F�_��j�X�$�c���a�n�'_6�SI���Њ���=β�|>�\�Mf�ͳ#3 ��>�f�=k����el��+�7�]��8��lY�ú,�|�����ćֲ��%|'D�^ ����³g�(T틕ЧվYK�!oV��l��鷰�zu�R���++3CZ�c�}n�d�r��d�7w���~�4L�G-N�ZV��
��_S�+�˝Q�R
d>����{�n�i��Rɕo�\���ý��^qk��{w��2R���T��"s�y��a�UdL�z���:�u�b�>+b�u#�.��y��N�s�h�Xa�~��i��]�/��r�{X̛�IݗhD��DMg>�n���΀��7"}Y���]��̑Ꙃ,�$�`�nz�>�U!��)My{n/�N]�z36\`Ό�]d���w��q���bjUu�(�i��S1p�t�����.��-~8�	O�g�aw�tЩv�V�ר������V�Z��(�%BAe V�:�>�M�j�����O�����W>҂\�'��Ϸ���>����G��s�m��TΊ�I��Ǘ��aL��y��x��Y�碽���}f�Wu�v����.�4|����w~�R�'�oz�.ٛ��bW����-ۼ���FEz��ՙ9p/�Xy+��*���Yh�X6��u�^���mӼ��X�({K��MSu?�����6G��}�!�/�fLn{ίfY�7�Ƒ���*��:=Q^|�&�7�y��h�v��I]ž���4a�(j�D���ik%v�|9�7w�Y�y�T���rE�m�/�G�=DXܢX��$�Mv����+ 0HJ��aػv�(7#�Ųu˽��v�m�nI�F�wμ2#(;[y&�jfO�����x��86!]��T�﷘� V��
R�����2�I���چ�n�@�k���]p��HD�rBV�<%9hWQR � �䈰Ʌ'Kn�^W��n��w�5y������_w#�y̍8-v?K���J�:x��wX, NQK$
���]l^��������o�����-�<�0��b4s]�r��;�پ�#�p1L�����z��&ѥLV��v��AT:���<H/ҧ;-���t6�����p"zJ����*��*m�A �h"�l������T��Y�6b�O�<�7����nMa�ԉ/ݿ
���X�t֥�gh�*|~�:֡k5q�<l�d�s׌|�&���Wۛ���d�aL�z�P���r�/j~w�<~Ka����	��cVz8{��Sm�2o{��.?V�vx�NI�/��������쭆�ğ��{�}'��w�1� ǻ�Uv=q�ļL���^P;���T�\�ruw���搓[AyU��S���d΢��=��w/7Uq���iүwH�F���'�`������%?���l4��l�W�:�".n��4�"|]�5sUIͷG]Q*���}:�Q}70����i<�iJ���&�a�ܨ�7㽷K^M�g8�&��ˣ�m�S�����灮����Z����y�Ogd]"0[���{�T�6D3���l���]����`oJ5y�l[���f_��ݎ�Ҕ�U��3��R7c�>��M��zpYo��N�̮4�U�CD	ke�"V�9k�BmQF�;j��J�,�ޣ�ƥK��>���ϟ�Js���]L�v�x��.���ΚΟGI%FU�J�;r�m_p4NH8Ʒ�i�+����߇�{�ؚ��cb��8�ɝ<K�����3�V�6o!���`c۹Y�:��c�)�IJA����8�B^Fev���K��yAu�W�a`���dԼ~5WU
|�׽OW�}��K���.���%}O�Ƞ�Wyr�RB>�9+c�]ݯ~�uJ�|M挳���d9�����g�\{�ۼ<@�2֣���d��T��:Ι�/��!���kX*'����S��I��)�G�dn�W��{��
�{}JQ4ƶ��笠�S}�~N�h�����d���g�(�͖��X;��m	�E�ϗ�{�x,���i5m���w���G��{�<��ZP��0�Y,�PvZݵ�dW�l�2�S������P�q'я��z���m��yf�����ϓD��7�(�ά�g��ylH��UW�0ec�Q�olnb�#m׳��[ )$��M�I&�]�]`�-�r���������x��6���ne��җ���f��x�q;p2<�^-E�v�R��y���^�}��9�krl�5�\Sܹ��ܸ���p���V��b�Q��Џ%����~midpɞ���=M�c�,�W� ��W�O�I��j9ݗY��o'W��f�NA����@ `�<���:�P)]n�p9�Gz��kS�Q��#��Q�� ��,�u1��P��p�� k>���~����S�!��T�f��֞�[�2��d�`\�|K��ZU�W���o���\|�=���
u��s�?�����O��#J.�w⻭v�)Y��+"x�������긕T�d����c��2!����.�w���ʩck��NIC���9�n+7#�R<)�pt��X��kv��vPn(Ylr�R�pP ��aC��u۹���9��錃�������2���N��zÊMӪ��tN��UO}�9�����w��@J���F�y,�ۚ�Ǫ⟆���3E�����=x���x}M�Eo+������.�f�����Oz}�j�:�
�X��c���4A��@�{@�Vޯ��hՀ�i�],�:�¯nsC(`U�^�m7�9˫C�}oZ�v�:�<���=Eq"��wf�*��ޏ��u�]f��H�6��G���_���J����!��}�O"����Ю�94/㹓)~!ì�����̻n�S�(W����P���㥸�����VX�v�8���K��R]ʆ-����"^��R\;�oq}OY��Xgs�>�W�)f�y`���B|�=��-0OM���.��+u{�ms��O��mI��ۧv���TI>�=S�T¹k�Uv́�@�;Y�Ψ½!�VL!ԍ;S.�z�|z����c�Ё#��.��Ȭ�C��߯�;��8�L�D`,0ܳ�l-�qWF�}O��C#�@HSN7��kc$ȫy�+�͇�(V����[�8�p7\>�[�"�%b9o�B�E���w|�c�Z��=/�H���,^יw{�^MGsn��,1�X�4VCCqꪼ���]�,އB�:�YG�IL�����3ր��`.����nM�X�{hd��<��^n�ъ��������AbvD.�+���w�ޯ{��e�bG�5̹{�pU�m\����"�ߟ{��ϲZ���5��V�W���{լ��[�;V6r�����Shi��J3���BkwW�5��RÀ��
�e�p���,u737�9<��륻��r�[�� �a�M�H�a�"�n��T�`�A�'�(��(������Yq�滘�Vb Jy�[T5k\��w �$QB
��曆����LS"yW"�Q��Η&!G	&M��������Rz,���K�r��V��Hգ ���a,q�٧�<=���T�虋��o�� �2�0l�/_��O�_B�~����u���K��CA� ��R�A������}epX����펗�v� �������|=�V}��L�'�v �y�g��ϧ�g�������Wq~P����>ȟ�c�b��!�bDt���~+�V���ͪ���TdMFY-T
/�ڻ�(l '�z��<��$F�L�n�lM_K����ZF�Z{����h;t.2n����>�^�����GB.	d�H��ؔ.�v�ռ)x{���-3>yT�Z��Ka�Vw�g�Tu3�'���1&���{}>�}�t<	�w:k��[���ٲ�ד��M�����d��3sR*e�v{�V@D�k|]�_b��^�C�A�����Ob��é�)�R퓎N�Z+9��J_����}YʭO�ʡ*��Uc�����s��z�m�sþ���}��n|$e
nWb��׷�߱5T����x�vG猼�~����͗��O����5W�w�`���!q�W�c�Հ�H?yU�+�ǋ��\��������U����|��.��y�Ƶ��]pJ<Gl�M�0�7�S��������<����Ѫ'��By�>Gv�$]{ ~�q��'5��Ӣǳ�NM��qvO��;!�����y�eY��at�Mڭ��%� �mrA�	�5����]�^4���{��H�ut�1����;Q�'��vF�N�G�n��@,j���@���Q�'�vz���R�����96;�>��+�xOy���슳4z�g��6g"�]E�LHgxE�ʋs(�$7&;˽�}%�ylL9g��i��'�Ƴ�;���q1�"�uo����;T��.�|g�!F�z'��@/<�I���k8��q��m�F��w�gjM�-�fw��,�>0��ò#-L���n}뗴H�h��!�T��@	�j�ͱD�F�\m2��i%��C�����^qB�9�r�1_K�l��ͩ��mwþ�֛p}��T�Dk�U�v��� ��ɽ�G}7���g���������c�~�yVu13A���R�~�j"�[�ܤlf*�4IDK+��ȁm�
ݰD��9��}Y�謿~��W��z%��g���˭����^�����{�S�w8�6�Qq��BM���׫zN9�4��������u�o)B�BLP�9�q� ~��#��]�']u�֭P
��S��l��T��Vu�=��ξ��.�wf�p� >{��@t�O�s�Jǽp=����=��J�	$oGn�����-Iҭ���a�W�w}dͳ����O+��r��@��:�4ڄ�����+���q옺F+>ov�S+�����5Օ�<����}Z����{74�U7��ó3�5�1}�	.����p������g���nZ��Iu�+��In�=3��c���WO��t������N 1K�h�ѽ:������W3>���i�|����ي���������BE�	�+�2����I�;c /��k��v��S�����Eg�tk�������c�)	J1s�v��yC���� N�%6�iaP$0�1�Q�IGj���F�z��tW'��U�3�ߦ���U�ռ^����m�ܽ9�.�ǜd�{��E���&@Q��#���l��^Si{��v�|�յu���m
��e�[|̽���gx��;u�T�4)*�sV�t퍍K�	 �G�Gx�_������͐���04S�,��[]W����엇5�#䶝��mY�]�duL�Y��b���.<D�]��ѳ9��:q��� �?����$)wI2�����OJ�Nμ����<�52���<A}�;��
�(j��W����[�9�W]��&"�ª2n�����'��Z��TU�]��Y:� A��<}8��1N[�����Wۄ>�f���xR�{�����&��v�󘦳eA2#���5� ����:���w>�ʓ���X7[��.�4��N�Ć�B[z�/*������o��WmeO1�m>q���]^Wn�A�mٕ�$L�;��Z�v	Og,�=Mv���T,lց��C���p:��0�bΫ+�R�=��fi�y哫;��K��i�DkK�ZQ��6��k9$�/+v4Wp�LS�t|������n����8��ܹD$�{@��5�g=(��*Jo��4�ށNJD`ڂng^�@�9rQl9b�^�e��j5�tU5��C�vz*<��s�Z;(i��l+.�C���(��m�k�n�����٠>�e��h�x�،3 f]h�2=���}�ԗR��vb|Bń�QG4+��+y{�x$����K��.hO��'\�Îr`�}���'t�S}��1�y�1�/tn�#��c.�Z��)�0�G��h�ԟ��
��W����P2i�V\�oe.v����c��o�=�<��T:w�`(�|���K��5KI@V��̙h�h�G~#t�N�H��`�l�!w������=�����݂��Bzc��3hKC����Aao���YwV԰F���	[e��R�]v3�R�ZT� r�7�-��9>�`J]b�-K�$�i�ܶ�%�|702 �L�C.�Nwp���ۦ�Q1d�;;`�����m�)Ω�ap�܅jt����,�R_#+=�y�[[ɼ\V���GI��M�Z��go2>1�8vp�FMC)-庨[}C\=��yC=z��uL����n��P�օ�mmc��q��ʯB�p�k�n��KOv`uc:ˮkb��ˆ-������s4�;͢�3Os;%���犇�Ko���Z��+w�}i2��h�˭���S+k�v;�fS�
�}�쏫�W.��)s�i���:������m\�]�GPr�γE-���$jb�����'r��F�z���f3�f�k�Q���~����󮔚{���3W׸�*��3}�%c�[����i�m�U	%s�j/ۻr��3�����*�4Ҙ��+ME��{NhOh\�Os�
�)���þM���-Ð��;��U�q�����-�*s|�ߧ���N�T�ө������k�L��N��F�~�1��(��b��L�����ƞ��,v���6=]�_C�7�����?|�S�TS�$EZ�G�P������~a�߂�aq#ުԯ�T�q^��Zң~���y=߉Ә�6���R�{~��eܧ�\�z\���ґuR��0��BcTc"�KiR���g�q�)_�ڼ�1U�j$�b�n�p{\��_�������C�u*~sM�;[y7���ٌ�)�;9�'��G4�OV���9C��0�S�}E*4m|��Һ�i{�v�v��~�$׻"
�,��e]��1e=�8s���m��f��:���Ng�dh:����;��9����	����,����x&e��m�$�I������ϏfF�r����h#��+��0U�}�V����%L���:��#���ה��A��k�kN6G5�@�d%l��U��ý�3$P(�d'P8�ݐM��z�����mj�'��2�t��a����ۗ"1��S�KeS��&*;���`q�R�v��.�?�R�M����5$|y�!�lW�yvh�o˘}k��6]׫��E�{)����F۶ܛ4��Q��uUW�-�;I��U>"&L���k"̬����٥�{�<��O��m����>�8���)��Y3?�q�����u�["t����$4��V���ҞBD^t˻պ�9�^��{H��
b{R���jC)l��Z;�_G�oP�+���s0�?��.Iڊ�ɟ�c��/��y�Ϲ<쁞��g
��;ןrr�kr�p(9ß��=P�cѽ��?�����K���s�#�P�35��8#����T����4������>љ�T�fI���K�4�
��z�`�
��<(_nL���sD������%:�<F��u4�r�Rx�b�x����M�
�"|k����xn=�(���gL8��ȥ�����@�@.r�\�\9�-o#��.����?ez����J�^7�;�sMg���';=z�ɛ�v�������z��nڧ�:�;�������p��N��5��]�P����S�,ޚeV�E恂M���R�B��gÇ����.*��E�Wa��^���WS[��̮�28z�CX=�F��O��i��c8����<y������5;���G�>%Z�!�ĝI	o��+�*c�����������|7}</.�{:�����#\u}�2U���ೌA�tu� Q��)f�J�p��3V�C�^��Q]���YVS�����Y��w1����:҅��Q�9xFb6�~��;�_��v��UG���z2�������]�2�&�!y"�cQpiZ�eF�|�z̗�Zּ�;_�qn;Ŵ�w޷�WU�f8 �[�׭ym�џ���:�����zߍ�G��U�:Pq;f�f��`�b2v��x@�����|(���y����馷�/�h�堨�{��e32�h��]�kg���I��)�=_;f�$r��(�6���8��[w��Wf���6�}����d�D��û4�z|ry[��z�JZy����A�m �0�c��!pdD���Y��� �[�P�+���S�>m�	����29E������3���~�
��t� �Z�43�~M�dEE`T碭'���	>���CC4��mhm��{���%./�k�����ޮ_I�������[ku��q(+�I���[�����BPEO�i�U뾃yC-���	�ˣB��Y�>ɬׅ�y����6�_V�j�(��o�_�8�}5���)ٓ��p�oWh1YxEq��k�PkB-���1)�&+_��t1x�k��ﻱzCȗ>شU��7��uئT����xOVSQ:��cy���ػ}K}냈N�����a�-���q�c���R=u�nx����K�($�榯9ړ���I,������k|Z��*��0�A��f�p��K�z%�]rǃ������=���*'C>���ӏw�j�U!u�<�kں�Bg��d\�.�s��xE�K�m�
�GL�U�s
��u�e�u�w��z8d��\,䵋ɞs�G��7���V������%_��b��޷$��0��%?]^f��>Z�"W�aG��r^�r�}B=!#vI��^���׃i��{`�M���+�	�ݧ�v{������>>�VX���)֍�>-x��4U�/ԣ�fC�>&�π���{�w�%�,t��2����<vN	���'])攋��*7��\u�A��ܙ��ƈ&\�����o�K\�Bu��y��.��,���>�kr$7y����H]ڜD�v-�psズq]f��cB�u:z|�i��>�:-�n�IM���e��s�!�UM�Yt�c'�.ѿ{�]Ֆ�
�э�Pe��K��o�3� X�9�V�]��%%��F(�NzF���Fy�򩑮��}N�tG�2K�[����4�4h�v$��3� 0����b��0�y-W{��$gq����ILW��>`
yƾ�S�T�W)i(Ƕ�m�.=�
��ڌܣer���/��q��I��U�\�QX�斘bRHT�U:�q7ln:�����(��6Q��yY����g�ʑ��u�Ƈw��S#vxtj��=ζ`FG��ȳ9Ʊ���@�п�3�Y�s�'%��^H�]�q3��7�����>o�3���1�/�cN��˽IP�2v(F��ͦ=�=���r������	��vg��q��L*�Qy��W����p�N�.U{��L���|��ss^�ӫv��S����+'#p�.�lZp`�7�+�߲��gc�S���e)�>�3ң��s$^̅�5�F����Hk��Q��2T�NY�U�_�5�wkxv�s"*�7�Z��ؔ5��}�Vb���\�����Î�I!����[C$�մ��E���ڃ���o�D�eቘ$�R��m@���}n��p�Gs�D5���!�e�
���;�� ���hcaH�,��H��3�#u�R���\��6V��5�Ϛ��R֠�Q�ڰ�
��j�����2=��=�s۵|x����Wr��`]�ۍT�y��rwa��� ����ޫѩd�	<�����$z�bWg3*81�<�%�
�~��I����:jhKF��T�z{���9#�&}39�F�wt�݊��oa.B�����ᎌ'�l�������{���df��1��e�!��t�D*�`�,Am�H�YC"rm�#Z�R��:w��z�My��{>���r.�i(���ڞ/��|0��~Ô�`j���ڧ���xL>QT�������7�ޗr߸�xe�)��4���9�nO������x��5�^Q��o=��-A]G��|�
�][�By鞲=r9J�w焰�D{�p�^wx��E�(y�&�u��n�����PO��`8�Gb��! �b�T���1��SsХ�V�:�׳S�6����l`跈>����V��s�^̋�̇�q�g}�L�;���A�'�[�*_ɟP���5X9z1��p�e=�e0�Z�O��ug7�1�??�\b��y��>n?Dsr���.^��T0XF��9- M�XS�����u��d&��L���TYWV�ۭ�j�s]z���,��uL�|w�*3�!^��e��n_^?�A�I_.ʱ�W�7��;���,ߴe�������ڙ8��T�όډ��o/G#r�+�ʠ�(�rE�D�J
�a��l/�l�^�P{_ge��E��d��t*��:�k�X��7�oo��Ke���M�FzM�-��g˙�>��}ge��B .�n��t���lΘ��3����3XI�]���V�$N�(��}���[��j��K����U��z�2p��y�ݾ�"�s���՗��e>�v�jX}�g�Qĩ
����6����ݬ=�w�'��m��Jف�0ǜ��ս;��6���U^vb�
�h]:���/�u6p��̢�f=
�2V������~�ջ�B$nGK�zG���ӑ��c�-�,�j�?a�}w���e�۞�����B�=q�3 �N�Ȇ���*�k��l:r�hj�^�Z9�"��柠��ִ��9+�O�9�����W ��~�[iJ�)Zu�n���cd�����}���=�f�������ӷ���k�W�"/����u[Bf;+�Ò�?�}���� -�r�{V�s����2LĨ�R�2�S5��e\eKN8��N����&*�oN�Ȓ��u�ggo_
4Wq6�L#������\k����͍9�0Ed�<�;��$8�}�=N��(w886�g��g'Tu��W��2*`�egـD�0w��2������.99c�r��(e�6Dy+}�lP��)Q��V9��n��b�������A�Z>�<�o���ʞz�r.���;T�@�B������������ҟ�?��KH^��ݩ>߻R<��3GՕ��/���ov�0��m�w/�1^݇��42��kWe-LF�J�A��ٲ�v𩓕BT��dH{Y(P�^6�s&
��$n�ԅ�dA���d�׭��=�L��4�nV=���f�Qpwz����Ue��XW��a�~�����4�E*����pA��j@ZH� �%��i7�]�q�E8������b7�r��@�ilY����6;�x�����兰H��?\�h���������;�a�q�ӂ%��_=�MU��y �])�����l���sq��<3~�������	'0?����t�?z9���/�Ɍ���;qV<�m�H��`�Z[zq!\�3Zt_nL��1-�u3iY�����+�y�{�`���HCWNN�4���#p3�-4ŉ������E^s,=���[QK���ǻ��&�V��j����������z_P�k��%���1�3����E�u����9�@G�������7�j+��꣯���r�iK����f��[��������>��e�c���+�������v�u���÷����k����`;��Tn<�ێ9q���P讙�y�I�)[ʭt���H{u5�x���*��X�\�b��\��R�����C�;g�y�n��v�B�Q?I��ｾ�<'Y�
�1��0�nH,y�^T!ҥL2A �o����=��h��
��b�����֍DV;�����=���F�-�h$��ǆ��i\�#k(��3N}'M_�z9^�}X�rѫ��J�[>��c���|�Nn7�)��+���4>Ɖ/
F���j�t���l�:1A���UCg��S#���1I(՜�̩�|>�x�*�p����~4Q�l��5Vi*�&��F$=��V���������+ut9jm2�m�M�賲���O�d�,��]s�|S�>�}�$S��
M�oҡ���7nN���تN��$��7F�	�:0fS��J�q�m��m�	ڼ�K��B�R��m�&#��l6�����]	( ���بbu�]) �1��r�_��pY(^�#�nvo��v�-��Da!4!mj�b���ز�`�.�+>œ�<��&���CB�bl6_
����Ŷ�WG�4h�Y���j�beCj��Ec�#���]v� ���8���s�ެ��1�Y^�Ɣe�ʜ�cf��;o}i�:ó��V7�|����1�)@�
����~ٲ7�5�C�I�v��o�>����{�l"^��w���)�F�m1ɍ	�t/�Z;s-DNM{=�<�!<�"S[�1�Eܛ\	Ր>Õ���R1�؀����UM��R�i����>��ch>o#��0�m���=��X���&� :�T�F	vs/m���B��n�YX�����&	��Q�b��3��c2��x�Mm��k���d�{W�Ջ����i\hpȨ��u擽k�Ƚ�]�í��dW��sy�}�����Tf��7�A�w��4|��_�f�������ߢ��.��tY����6��Ҡ:���� �3���� '�O�8z3>g������ʉ�U���$�w0�\�M���X^_LVFf�O�v��n���{^#�kе �g�9�^h����T�ݝ;7�2b[�+�nkhi��]��[���)�5�u�^��ߴ�mr���?u4�ѿ�Nv�k8q�����{otBE#Sjvju�{q�NJ±�7(J/����a�e,��Vp�S)���,�>u�m���|V9�*��sG�!��:&��i��G����ν�������3L��]u��V��ja��֜�<���[6#f�6Ƭ�ڵM\8�fWd��T���{���֭�8Gʆ�;K���G��m��spt$�W�n������s���X	\0��ɷh윲,4�Nzp5�9M��/�fh���fd�n�=A{�G��{8irnd��� 3lo;� ��#�������+l˻@�OvsHc�-Ҿm;<0A�[�,����'s��(�m��' �c�����j�ޯ�V�T�l��uuD���wIo]�{O��k%֓[��$F������c�ZΦv�q�i���x�Ԛ��X���ð@u�-�u�3*���ivW&�U��#h��R�j���x��d&���C�h@ZCcj%�x�R� �4T�ݭ��1��TD��q#$��,ő�������h�p�I9ɔ�7:D�7W����_����x"��^#pv��]y0�[Gz�ml�����c̩��=QVQ~G6�.zn{���"�E�xx7���y��wr4�^D��-��qb��轺Vb�I^;*��$��������k;����cH-�#������a�h��a�%�����ݤ�x��;���          M�4�[��K1r--ڹ��8��H)M9V���*�n�VP���+\qR�Y��+o	���j��-�uжB�'��tYB�P�$�
�G��5�YU0��	H�P Ȃ\v��J�ݬBt�cI8Q�M�/�. ������1�E�%�h��HЎy����!�	���"U��#�D�1���v��k�=���]ҘAīg1���o��+N����W�����ܫ#"��˾$���˲<��1�q2$�<P8�"��U5���ԛyK_�����Y�*,DK\P$0v�!�I�_�y��ڡ����j�Uac���$J�&�4�M�~#��ۺ�D��TR�oh�[��>5C�m��TE~"Rn# ��
pqxY5�o1z�^����M2�:��[z֛YP�$BF0�i��ջ,�H�
���[mp7�LaxQ�n0@��t�*��۹4oD.tI��Rq���a�����2J
[��6�Bц��>:�����;R q�w���cl@5��ip��qj�uQ�d��%X�o+�d�@�6{xi(q�P��*�R�)�;fH���X��
v��8G��g��haU���	i��rq]�&�Y!��<���pE	��پ�l2P1�(��AF�!-.�+���}���7��W�
U��H��v�a�Z�}5�2.3�2��hH�b����h����d�d+� ��� ��IM�m�P
Uu7 �}g2V!f݁��z7���H�Sn�`�z���bN�=���.�	��^m�I�I*���X�u�≦��&ʒ�M�ȇ�Wnđ(�&u�.XF��Q��T�����SDf,��1b���2
9��@�ڳ�RSV��B�M�y����Yӊ��Q_+�jb��^����r1���Fq]��Ux�.�1����hb�Woe*U%��⦕f����Yy�lX�����az���8
�j���g�gvd��欙H���h釒wŘ�� k!]��k��-yvs�U�e;j���uq �2f~���J�BێUxDf�;�9��f�Фbk�--�&�m�L� i�4Qb#'������i	�w<Ut��`����D���S�\����D����x���M�h�NA>�GnE����^�erP�۾�sI��0z�DH��>��۩!��T<{޻�0E{/��(�k�"�k�������+�ݧ��������QU�nc��35���!���`W/o��zch��o)25�Ȱ}��I媼:n��7�k~�þ�J1����5K��K�_Ҿ�|��+�ó2�en�O&㮤zi,>�!���������c�w�����x�6kaQz�k���ݯ�|=��[�ڳ�UZ^�����ڻ��]wR��o8J_m�-z�q�	�Z�P�3_�xc���Q��
` �<����)es���71�˶��KO����T��Y�U1�b
�7Ӎ`�a�@tؽ�ݸ�l�q��=�۹[��dߟV�Ք�9�j^�Fw�M������k1j��_6�Î��3qf��b[���e�ђ.������V�������M[4��&�K�獭�f{�QO�Ϟ�@����gX������Sο�g���W���ϳ���7'n�idF��3��F����(�M�X���,Z���,�o���w�woNW�"��͎�v�)�M7ay���z伭�d��9��8{]��ݭUzB��� Ѝ�^��)��f�g	1X�<��obS��ŝ�(!���z��®��G�%�^�x	�5g��D�L���H����^�.s#Ak&�����@W!���3f��3h����Uz��q�0��v�	����.nk�{g"NGF>�q'�Ϫڑ\�b:�9~�:q�V�q`��Ցk�]�}�!k�>��������Df�ը��FܡA溪��!����)k�tGg��Z�[�Q������[���xa���3��r��{e���A���o@8CZɗnY	hƟ8"
�K.ZJ�A�@9�s)en᠏����J����lk[+K�b���f��W�j߶��;EdUi��|O���ly2Is�����R��z�������/��<�W-?j�oU?C͡������DT�$�0���z��ٵ1��=�^� �0"j�zħ��:�2����,RS��=�L�E@��Ԅ��֗s7r�%�?-�;��4m�kv���(��oj�D�(�M�C�P=�3�ڟ��n��\�����cOt��f3"�c��i�s�'���+/mS�I���{t�+�B11���[VL����'���,r���_O$�4���5p�}9l"��˪����a5����ɹ�zD��`7Sm@<�/��d�U�χ*8��{���U�GR��.AJk�w��a����e܂�z�Mmz�< n�͕\i;��J��lV���z�����Y0�8ָ���Y�kf<�Á`�+S��t����;�����9KM���CȎ[b��Y`���nZ|:�)���R�������^��y�kv3�^۪ϩ��Qp#!�݆�CI�ȩS�͸~k)���{7�I�>�'�=�1Vl����K�>Z���$j�,u��OsϚ���D��ѷ�@b���d��D+�S�3=�n����b29̮�?�ԥ\�oؒ���҇C��ձ�~��AZ����\�R�i��������0���{����~W��g|����Jt[�n��~��owzv~ߙʈ@������N*�ܘ�[�{�q����ԇ��6�f��Z���%TУuaQ�����e4ʕ�w��9��n*�G���S�dR���&7�q>'�I%���Mf#O�Ť�0��Q5���ØNHa���E���b�	����5q�s�-��Ie����a%���\���	s�8�Y-U�3Qɐ+��i��L�6���,�v��.6���"� UHB,�!�OM��c�%��C*�*8�!dD�Q�u�2��~<��Ӄ37�i����?��u�Tt���%���Cݝy��j�w�r��]eǅLS-�b���n���=�^���Йr��f+s�wMV^x<
��뛀���y�b�o�W�S�L�T~��Z�z�6\Һ�Q���s�j��d'���H�\��A:��+��c�� ��P�����cILym,�Tl�w�앖�g�9��w-��,C5���v6j%��x���7��$v�6���W�;n}�^u��V�ߍ�6b��dc[~��U<�u�Gfk���a���y-�AP����� � ����T��F�.6W�m�YN{2�zFncy�F�]�����֥�V����{�m��P}�^G��V!fs���UmWp�K��Y��B�7Xp5�U�+�.na�x\,��u{�{�9j��W�\k���Z��.�]c�	�v���w�=����쀺ʞD�y-�C��h�_�#؎���~��J�ɨs�f����g��P�@����8W�Ҥb.�]�nD�RS蜀K�{ͅ0�1q���S`]֚�돺�7`��B�OR�_���)x!�[e�r`��1�ۡ:s?��ԩ�Yd�����F�6��1N��7���ۙo����cXɅ�/m��|{���J�Ǧ�Eu,���{��C��N���v���^v�W�=c�+9�4A!"B0�N1�B�#q�`UhѸ���V��~O��o���>�u9�nv�*Ζ�ַx�&��hf\g����w{�vG-���^������X�Ě�U��
�u�{S:���Wg�Z���婘bl��ro $���F}u�g��u��^[����Md�v�y��뺝!����5�� N�?;�}�;0~9�&W�u�@����F�ک�.��鶙�n}��++ޤ.�E.-��.��w ok� �2	4z}X^��	0��5g}1�8��&��7%�$�P��M��O^����q�YٕUz=��C�\\k)'�^��@�O�������2������}ND��1�i:��̄��8.��@�ʾ�ö���V��%/�1Z�g�c�ʗ^0�m0��, �2�l����Y�Znc�-��4�j֊9lm�D2 �jB���o���z�iNwz��7�'!��ʗ}U���Z���;�ǿm�4�t�`e*��ӊNˀ��*(�n�L��m(��+.y��7qT9�9�g8�(p�	Mԫ"Y%��wb��ɽ��pk�]�#� �b���M�&¾|t&�h��c%�;yw��i�i�eR�uGwP�[�͏S�r�Msܮ�S�5Y�2C�n��J��;t'*�������/�|��l�>�LWb9A�C �_N�ƌ�/��qC����7��-(T�%��~���
U�̭E�fvy�ױ���F��c��˧�Z�^��nU�PI]�)��AQwVE�߭%�׾D�`�5�t��9<^���#�jm�o��r�[�V����ey\��eX�;�4��%���l8�~G�PY�����.����s�}�������-�3���������b{&��)3�ȯ\�;���AB,w�5N��W7��7�(Ǫ��}�'V ����R`5^��@��\~��F��s����R�z+4R�CX�Le Đ#NJ��%�3��D<�#S=����O�hgLx��w��*��sU��Y7r�}r�V�n��(p�_.��%�цp�Wt���+��ܯcy��]��Y�.���%���&|߇����[�h"E��������[�[t�a{5`�> ���.���+�ښ����wT�*d7H���%Z�Ɨp2��,A�Zi�oG���C��j��Ppl�\F��r�v,In�����.N��=�X6�#z�.�]�����Yv��w'�_9�V{�O��>�����hγ}r渺\��k��Clb��Y�ڹyl�mOS;�j��uۖ��;u��)e��^�_�'N�P͙���17k�K������^��A�3/6�k�v�Gw@���`i�8�UU&g6�����3h{;7�7��]N#�%�žSʤ����7��j�s<hs�Zo=�﾿�x����繜�5Ґh�)ל����W<)Z�v������U��&(P�A�Γ�W�=���c�S��7�n��ǘ��=򫚔2d��+=����>�t{����K>���(=��.x���޿�E\|�N�"��}��F]uո;݀s���D���Vޅu��i2�b΢��̃���@��T�bĩ�οd��<Y�[���}��]e?C��<��T�x��^�F���/oa�����eO~x&G6�y��~�7��w;�!�'�����:b\��� f7�̰vK�]��@t�A��Ҿ�S�n��d�"�"�^kW�bg�>zs09����ۙP�-Y�n�^���Hl�J6�q�r�R��U�u 5q"vb�bi��\�RKE��ַ��3�Z�Tᐥ�������n�\v��&4��4_\����W��X)[��\>��+�Q咫9���Lx�P������L�9�%k��f�pGL�J1SF"�B�)f�EF�B+�I�{��ي]iV�e5'���B��sR=Pj�=�F�h������30JU����,��*�����K��/K^��=>�'C�uk�����_!�$X�'�I�}x�J�1�G���S�)b���N��-���aF$����d��ΘJ�.��m���W���q��8.[�!��1�mFV�`����W��uM��g���F��\��"�GL�i�wٌ�1*4<��6�rG(�х�2%�%Gz��]y��^�`�
�\Ϯ^�����y���wϭt�D�IU���N���x��	5С' �����q�$�1�3�G��Ӽv&�z-��T�O�<n�2�e�����:�L���c�1yr�
e~���7��|}�H�Eֈ呟�pǱ�n^N�$�5�*޶)O_}O,hi{�?xНbd\��f�_zP2zmkOP`������[��w�P"o�G�b�ߙ|�v�2/&.���B���~?{�e�t���=��W5W���.�}��t2n6���%ĻoᛱA����sv)kM+�1X`u�z�d4���C���M[d���GC#ڝ\��G5W]V`�VnG�ĸUޖ{Q,�r�ǥ{|뚥�l�`u�x��wWw��<�g���.������;��Zb�������������e�Fto���0*"I��U�d����(9��Ѿ�h�0�7��)i�Mi?{~���~�O��W<�|Uu
���I˭� Q"+�۬��	�0�}Qq(gu׬��(��z%}�Go�����&��>�}���3��)���r��s�E���ҵ1���J�5~߉�)N4�uaw/�aw�L�}�����o��L�@$��"�՞]۬�n�4u����\k��'�!��Y��5��74�S߄���,�Q�	�݉�n��c�S|�6�,�x���sb�������|O5!�+�}B��jǃ�ǲ/���C��Vq q�q��c�-8lg}��_L������{�e�z��3��_����{u0%n�Az�E^/��\�/iyZ'��~{Jwo�ߍz�������.��r^�ٸ�=�NwwէT�5(���� ��e���-usvO��G"�3enEf�n�]�^���:�z�z��p7�g;jwe����^��,%9T�.�8��nMya�d��*�Z�N)���Z������Z�f��p��nm�ic���N�r�T+$W��
Ũ�忦���Rj�G#6��Ņ�J��6{ʞ�}+[CzuJ���p�͙� ;_�kW/H��]���w��:{�{�W���|��O�z}ɀ��46�g�dQ��M�����o�U���n{`b,�62���qu$�A��8b۝=���3k��ԏ�c�iUr��,���#�|��T�*n�k��k���E�>#c�wK�\2��(��ޫ�{��l��m\���r-�#wB�(g�ui��@��{V�1��y��¾~7����f�w�gn����4ە7�,���`zz���޴!nJ��{J�Z�������4:ITfP�(Ͷ�u���W��.=0��}�~
ȗ^�{�%>���:���qO��m���~�Z��u�cb�A�� ��0Â���MmH��:�Y�(�~y���3�u{����o�ύ`w�%}��}n����u��稟ίq��T
3ꂡ[��!C���=��e��{=l.�g�H������g���w��ѳb_���b����5{�:�?~�~{�Q�Ex��,�k�+�y\��ú�~��$��ܕ7�Oǆ{!"/eP�D?l�)��~�a�"�XYP�K"T��7��s5�]R��5�V4����5�vɉPHS����h؛:�'�n��iSc�^É��{�Yku ��@���^]Dy�{�w~��&`�r�%�ᕼ˼�:���2c���n��,tl��6���*�#d'�렽ژ[I����>��E]�(SƯ��Ѽ�++�]�U
�`���o@y�f�9� }ܗ�Cl��L\�3��8-�Hv�T���ZSD��	&w����Yr����y
ܓ�GN����\��w{%^ȍ'���T�(Ǿx�}&û�T�����RcV����MJ{}�0]"��Jt �]]v�Gq��R��j���d��Ns9-8+�M�O�0�gR��/��{�砭�kp���%�ٽ��w�P��"�*���5g�>��r�WgIP_�X�/���:I�+Z��w��b���������7S6-�m��G<q����r��o����=�[^��M����*������95jI�sB1v?z>h^
��3=C����7�B�f��ʗj���r
l5tnt�<FR����.���lA��[�[��UCS+� !�P٠�E�%�;��S�r�"�c�j=��s��ۋ���/�ee���-G�X�}6�ٽY�\�h�c%���R� ��J�K���t��tܤw��Ek��em��qN�|x���\V��]�j�^�I��~�1�oz�J��+d�Mo���2N��us"���n�H�3�s���/���2p��,��ƺ	���<����}ʡ��x��v!�%#�՗���]��TӬ����g]�x��<:so_o�Q�i�A Ň�K�A�:���oo���c���mNx{�kd��jQݵ��Zq��ix`uPt8�oww����W���m�}/f�{w$=�oG	���7-j���QJև�uT�q*wNǹX�{���o�U%t�Z@���0�z���ՈNE�Ő�L�'U������K��y�ٵ3
����<o���=.?JOӖ��g�G�ܲ�.oL;��m5�O��fqމ=��W+7N�5vd��=�5~��V�\�ɉ�ɑz�OT�M��_Rn3�P,x����x���7H:_*�S��#Ǒ����y�7솠:� J�WdG��ݺ��%�ײ���~��}�K���o�g�(��Oa8���Xr������u3⁹��#z�jhjN_/Qj���32��t�W��t�ӳ��j��<r�W�%��O��������';� ^��\4=3}��ʕ�{�)�������E�=�h�Y�`��gې2�qElϞ�K]x�=JBΣ��?�HA��J_!M0���c�#b�'�D8[�H�?|I#w��~�]����xh��N�a�G�݁@:Ml�b{Z�c�_*�:|�Uӛ�c2����p�B�"W\�`z��_��ߩl��պ����D:�F}���v��i11�|&OR$lj�G����O�Q]/Ug�F������n�E:�kXa�S��8�$���?7��܏��b���.�P��c�n�;�!\�;�_=25��-V����jg��ƀ�{c�'#ˍG�]�:<Լ��S��{����v���'��P|����|J�k�f���e@ܳ�l�� 	�+����,����'1Ơ���Wu�e�YXF�B�x�b������`��)��|�a�$奥�$��i8/է�f q�{P�Ț�1��tP����1�"h��ޓy�g1�*��5!L�N�`R�tK�����PHS%�q����yr��9�Q�a`1d&��w+�q2�! �(����Q��̔*�w?F�K�@�*��DVH�Ƿ� �ms���r�ދ��f�52�Gn)���w��E��J����{I[-p��Ѻc����s��)��	���e�$X������\�s�^��l���l]�؋6��8|`��V(<z���o��8!���IWmI�g]�֠b��Э1S
�Ṫj��4�X��T�Jy,�]��L3�F���T&�D���
w��Q�|	S�m��ڬ�)�	D�a+��@��&}���ϵ��z^���O(}�����0�]k��fJ:uhѡUn���&(���a��^�R����%�XH�8Ge�2�a�.��o:�7���TX�tyгQ�LQ�R�M%;{d�p�U�o���fs����o�fE%uț����(e^2a5'�� ��?{73��]�V���{��-Qi^�_S���Y���m�X|�17:�ɝݜud�_��g�]�{�<Dj������g@�v1���!�R&��PR�ǔvb��S�p�S�}��.��/�K�cW�F��1�X�$¼�Ȕрɯ!�Mۙ�źЊ�#�J;��a_{��}I������(�Rw)�B}t{���3�]j��r�c�67ǠE�/�Z����wڬ?`ܩ�oUO�M�k!�~��u�P���C�+�u�h�{!����%V\Ů��eգ����CԶ��]\{L}3x�-vn��	�ee��Wq�ͩ{�U��Jڻ���{��1�H���s]����~���&�Z5�G��X��87՟����Ӫ�ϫ�u2�H�)��pϵ�v�@��[���2I
R ��I�H Tn��+��;�LB��Z��3�=sL����R�O)���4���*]O���(�{�efi�n�W�r7�6`�R�g\��>ح��wQ���x�yR��:;r�س�2�o-�譖���7j�4<�'����N�c����:c;ǈE��C�:k�k;�sS�/�4<��������F��IͯM]Z�T2MYuQ��ԕ����X
��/K�ʯ��h.�����a�{5Tr��8�=<�9��nJ�4��;7���*�-���eh3?R�-�{�K�F�xe��n���ʯ� ���3E�ĳ�qX��Y���o����;K��}w��/���ɗdݿX*YS�Bj$)涀䲩u�'�ӣ����wrԚ-�b��C�i?kȿ��Y�!{�m��z]�8��]��m�!�3��&�s���B���M�x��T�
�8��lG!Qm(mcm�e-P���Qᒼ�s�/W�9ǿ\ʆ
�^���
�懻W����n*���fyRu���߉�3�-߼6�F��I��T���2��A��������M��T��V���8:~��+�sM�wV����P S"�w3�X�y-��7W�/�D�)E�#JP*�乊ksY����D�ｑ)�`�Q����Y�[�����5��d�93:�{K+��j�q�B^M���f.���hW1'E�,'���x�l�?e�Ƕ��]Ivkކpq&Jr��8�}��y{�E�<7�_=o�]u<� ��<w����~��-f�4�(r�p�Χ%<�3vuX���"Oh���V��;6�4�_��2��.jB�o��Ye�=m+�-��q���#ٽ�m�HeO���{G�Q�E�C\�С@%�o�tKu�;�e������l2	�������oe:��27��S����,��������B@�<�j��1���Yf��P�����֏}Ji�ڲ=c���+,X�� �6�x��Tz�����-��z��?EjQ&�wMf �e2�}�������߭0	A�4���1Z	�2߄�P��I%	/\�RH��5�/�gtƅ&'S��\_����P����ex<f���� �{���FV��v��h�Z��'��ʎ�+\�,ͮM���,N^v)��'���Db�l�J;R͇�{�Xk|Eט��UpU��-�B�C�U����y�
�f�Q[�2f�w���c:|�����ѵ�>2�zPwC&�@ef���i�t/z����	2�͹��{�յ����RHo+zq�����!�q2C����WM�{˚�)K�Ѷ��M���θ��K/�;{O��za�~�c�C�3���)���d�����d���2�̕n�;�}���t��U��������F�L�`�ǵL}�=�
./4�}^�;�cmW��D*tߏx�F߶C�q����<��+��>V�L�ʧ���L
=~��^��"/��B���(������(V��b]�w,��j�ϣ��U���\Mt(Y�T|��ם��Ƕ˒TN�0_)�t>v�ķ�أ�����c؁�:&�,3Z8��	�,0˒�y������w��=���ǩ%
���m4
G,�H����S%c�[O�
ж/���4x�����^���4c+�OS�G���:�=<^.{��	�o]���"j
3��\^��a�3�����և�vM�z�n����{9@�w9EåS�jv�!T1�}�{f�)�'aC�G���W	�{Rۼ�Y:VV8/=J�-.��*�./�H�\��	�S`���t�P�N�co���//�fW��N�,�ZA��N����Yh�;�^�]Ifܒ��{sRף��WK�x0�V��'���oU�{s/*G ��!�A�j�k�w�!�z�s!#�88o_��&��u2���B'[����+����*Y�g���^,�!��AT#h�������ˁe���Òz"Ҡ#m�Vr�m
O[λ��lR�m�#��YR���H#_�J�3r �u�D筿۽O4qB2k"����s}����Ά������`��[5�d�,0����"���>�Z�S��і�Id��W���W�sX��I���E�TR���T(B�֠j5K�L�4�"�bem6��C9��//ߢ�(S�N�d�'n��S�n�z�*�&,l{��~���G�cN��i)��Exq�$g��V�k� !�ok�@p������r��lԌ��\�	�_��ܸ���. �DG��H��ϐ�'��������Zyq��\��@�g�4���1{���E��Ɋ�ح~��I��/�cq�$�ؤ�n47� ��q�2��6M{�ws�ظ��-$��&r�ÍT[t��a�j�S8N���^�8-�$&o���uq��<�Jz�cq��aA�Tx�F}i�З���N[w��^�[А֓�|}S,�k��L�A�\gE�����D�sg7_[�ח�2�OG��sg�0<�"��o�{M��U��8�W��y�s4�NPo���� �v8�Nz��Nn���l�'jU@7�d�\��e�1X���E��y�к�bMFl>̨\ۧ*��w\_���d[�]p�x��#y�:�o�&(=7�
�0�w��޹�<7h{�?K��Z��f��dY0,	��f�\w�ִ��M�WU=;7���9���0a�Y�6�縯
��_��7M_u��槹�h��[���:��+��M�z���T��P�y$.���{���9VeU�|̸��[J�!��;:{�u}���bZ�Җ�V��M-�x��~�g������=��c�˭g�}�ȷ2#
����gkUԺܮ���ٌ����-����w�[�7&DL�/=���}�@�دS�[[�O��E���X��ߒg F^Һ󌹧�/L憐����۬,��:�����u��$�1�Z���d��$���9�{�����&�1S�EϮً~A����	Ƃ�{u��<N[V�����݈S>�yt���Z� /zY�)�;f��i>n�%���� �����x�j��*��螷���؋����0w��2��sxP��U���CE�,7��kWv���|>��-��;Ro/���4�T�?,�B��|}���|V�N}�}�^	
��f*]�>R��y�q]��$�Ew�n��Z���?zJ�W�]]������=�f78�`Á\y<�B7-�h�Q-�u����+���b��on7r��ބ���dw�5�!�E�`���}��뻟{��NםI�nՕU�P/p�K��AG!�oh�Sz��}�ͯ��%-�BO-?/���,S���������G���\Տ6�>��O������И4%�����u"�.�ou�h4č�N]7���OǼ�c���.��8�O��يCܞt;:���+����}��}z�\�W^"�y�8�k�V]xڹ�:�N�]4�2�m���}��d���	�|�
Bq�vꦓ������A�њ�>E�u�^����;��T�0��)�r�/T�;���}Of�3��&umA�S��ۄ�"��{�.�F�\jk�0cO�`�����.���a��m�u����gP\����4���,��Dz}�.�ploGw�����
i����/�P���Z�GUuc�m_��$��_��?`N�(e�뫆L�t]�b�i�'�>�y�E'al���N �$�s�)8���4����E�`�/��3V; n��֕��5�!~��Y�<��S2(��L)^|����]����wz��6�ҫ{F)m۠H�"+qf���c�km^%7+�z���V�(�Q3�$.��l`J�K��|1�m�]_���j˽�O�P]-]x�+w�Z�0����7/�b�zGT�߅T�bUe	�F/8$��;SYV���R�׶����S7I���罦��x�}y__}ZC 8Jk�Qhנo_���k���;��Q�0�0&;�!�"u�S*�8��� OuM��/�)מ��n� �xFW9�O<��o>7�>�Wp8^��v��v�W���f1�Li�'o
�m{�W�L�r�����Zl��4�O�DYl����n�r�-��i�Α7�IT�}�_z��K��ɩ�;M�a@$�ѵm�>���"h�4+��;4��/
y��/��ߺ��h����븠m�fmMg"�q�p��C�ަ.� ��]��=������^�S��".�}��,oq��{��uLҎ�9��sz>˹ja�S�ʚ��&FQ��ž�u�
듅qG��'7�������J)ڼs��= _%ζ�+��*���s�zi���ѩ�aݼ� -�W�x��5shV�ߖ�+����l���s>��.\��dG,�}�:��f�ۅ���쀲5$�X��-l�Sr�����*r�T�o��Y��?K�moP�֬��P?zv���-�`]��A�8�m������?c�"g}$�O��Uϯc��: {��=�ڮr���،��M4�
��A2c���>��.���i�[=J��=Ja߳t����<�TLn�Ad�B���2bp[�n·zո/���9K��ԓ��c��až�Z���׼�ÉOv��K���Pp�;�{	y��Y������#ԗQ��6Tg'ge|sC�o\�	����G����z�A��QC�����`U�2�K+;���d�m��/���ו�F�ư�p�cl�8�4�d&�A�	�6T�$�[%�g�,�����?���*=�]8��-����b	1�6f��nPU��"����?Jcph�ynv��w�}�eί���N� �Z��_'�ף��Lc~���ÙW���8�]1����40���}�t��Jvj��8�\�Wѧ�deųT48�n��.J�l��V����8Y�D�Z�h�>�.H��3����i�3�*vդE��]��MԵ��V,닪Q�Bq�q�Y��3����� ��.'�ވ��+5V��?n�$R�$��,���[����.Qv��zk�G���<k'�����0D�s>9��'�*&1V;:�4�]�;����De�a�:�X�99�\�A�[��V���f�x�G��{Ӟ
�Y�V�ٙ�۵ч$�If��cEM	�"�1F�GHB�L4��%R������69]q��P�fj�=����VZ��|p;��m<�8�4?�����[��SӢ�<Jl���f�J��׉� yֵE^�S"
�P���%����D�yb�����4LK��ж��.QV�M|�}�Ǥ����x�����sR�ˮ�>vG����m�]ؼ�{_�٘~�/ه]���Сc�1x��|��;��
�b�k:;�^!S!��tS��}�)7�S�n�Q[Y�R�$���ld����s� ��
L�͉Ⱥ;�qU��2:ȐjF����7�|Y��5����g)�ZI��l�i�~��6_�e�����7/��&��212~�zq�����'Z�M�� �)�?G�_��3\p��U����ʝS�h�(&�����z?q�6;fL_��}��y�R5+�g���o}Up�����mw��y�*%-Q��r\���A?6.e죚�쏇~�+�꯹Ωv�U�>Ϛ���L�3������q�fi�?\��/j���G�t���2�#G|m����2w�-�5�U([y�>#D���M]�ە�5]�xϯBF��fiΜ�m]�:��0oL׏w�S#|�y�9�mݚ52�lvxx�ǟr����|jfvEK�W��fG5�`�O]$}�����/:F�q{��j�uN��D�ccO��j���B���]�Ԅ�z����&	���k��z�|��s�7���¦x�C7�d��"������_��A s��U5���`گ�l����F}�z�	`��Vj ��r�&�u������S}\^�]�-J����u6��[�C�X̢�n����u���yPb�&(�I[P�]!�j��d��䚾�mb�&��Ф{ݬ���^S���`J̊��CҬ>X�9'M�N�}-dř�BE֟D�n�z��筃���u����h��Ǒi�6{��!z-B%�=���X��σ����������\�z@�z�����K)�[��l}�*�=+~�NYH���z�Kr뭈1+Nv�(�ʛC�'˧u	/y\�Q�WDU��}8��o"�c8e�ݕ�Z��d�HQkq=�ɚ�����D%*̓�J�]P�6���0��|�N�W��f�~���[��.�>#Zs�^Mie�*���X�d� ���0��PH^Y��kukf��{U*w{#�Ns��������,	L����ǳ��W*_䌮wJҕgf�����K���m�ިA���f)�N�Sǻ��e�.u��I|s��YnK��)�tR�^j���\ �c�2�8�Dꭿ`󺷗Y��Y�ӯ/�`a��4\����N���aaڊ�ʹML�DrQ+�)sW5�t{����z�Х���_�oVڦ��d9w�g�q,��C��f0͊��+�2+U.W��rv�e�A��U|r��9`��!�B4(��CYx��v�
6�2c4��V��.��e-�{���ƹ~A�ʜ;V�s
����U�8
�郞18p�u
���Z^�@��A�����F`��^� Wb, ��� ,,         �i���RY��
��}:�=���b��\��tH�*�+W�����b�X7J��880"LYTh�]�˱ҵQ�Z��Y�d�{X�ܰb���w`AB ��
�j�YOb��ʚxVz������ʞE�����x��hfҾ&�Jf'g�ˆ!6�o��.
U$V*��u8l� ��v���Kj��9i�RTAT$�L����B�0�o��;h�p�e�w��/����,6��i�.J�B7�z���ta�D�%�,��۫C�X�Au���2�kX����B�WڮU	��VG0�J�+miP	F��JƄ�]07q��n.����3&�1Y��hfws257U�#��7�<[^�6�Y��ۅ��n��f���IH��%Cp���s����Ǉ,��J�חyTWVE�R����N�0{�.�<L��t�=6�n��cX(�U�;qJ*��+g2<��F4+ة5�XQH-\	FI�&EH��ICB��&NM�ˡ0�w��G���<�O���t��(�cg��ʱ�q�h���5���dn�l Y�2~�h2 �X�?���vn0́G��h��uJBPt;�pU
�X|�L�*�&�Vj��Hѩ��T�gy1o�b���#�'��A'i/^�4�B$l��ZZ��=݄`Zk!)n��h���xn]���)4�� ��oL�8�� ��U+�N�-�b�<�{���Ru3�8Ib=V�c����5���bw���L��@j,J�тBCJ�-�b"e�C�Nr�����^���:�Q�mF��Yi�ٴ,�m8�H��2��e�,��@�
'��c5D�#���1�cT!P�0\22��& S)8��k��$*r8��K�2�\���)�I� ��-DP�yҧb���nH�2h���;Mf3G�q������f��E���+�m4�_r����)�(�]�:h9��v@j��n���l�봇gX�>οW�����r�R��ˍ\�2����C�ag���N��u�+`������^u��.����N������O����̕1��_`�v�x�d	��"�F��QT喸�u [d����m~5�{i��譼wA�%��:��x�1�����u�SW����Kݑ�'����!!��=��*'�}�����i^K/���@t5����r���`���`�\�{���2�'#,�5��:��*���䮹)_�ª}m��ۃy҆�����56�sGX�G3!��%C��w����ʣ�H~�����q�i���TҭH�,7[m@px��吷�U��
�iá��]q/�ǳ�#:ꦦ���?@�ĺ�x(��	���o�pUwX��IƹtH�۪s�	[��~�'އ�nd�oS��`�Y�3-]ʮdw��s�$ŧ(X�W?i��tEˣ�<6��$��XI@���5�W�#���Yr��ءv|�W�<u�{8�A�}���U�]��U�G��G:t��1���eN�>A�cv�U���Nr9�܅��t�����Ьv���m�?J���D�8����`��D��5`�]�,^��D2��IEX�Q�U�$�_�U,�Y���G̜�7�ݶkMH�����4�)��\�.�+��S_��<��7�};�w<i%����5²��A����u�c��nu��ԅ��6�n���W�3�_wwI1ʷ]�i�͕��;ܗ�cpj����^���`ző�*@��'��']��=���nB���T]��c���u΁��ߋ�o�#���z� �'^�yt9t�s
�z4�g��pY+W�����$���X7�~��=��&������ǧ�^�6K�L�lЫה��8�;�݂@i��5x�si<)�8�Xū�f�5��}���� k��eDQBHWF;�/))xb'�s�1��Km�8��}��}��/�N�t����˛�Ӌ�Bɋ��"+�pkM(
���8����N��۸���e�k�����^׻o�W���È.���v}u�Rt�:�&��]��v����0�_-���Dړ�P2�x�a�^1'.�b�IQ��������_6:��f���)?�?����x%RI]���zt;���wP��jΜ)�^=�5}�-�~���5��	W���}�ꭙ���Mu��s"zoa��Ư'��y�����Æ�xU1:�i��5^9���R�7�s?�&�����ց�&�W��X��/��t�M,{�O�Uǈh��mr�U�%��rWf@���d���^1gO�����w����U�or�j�G�qR����N�϶�W���s���]�k�k\��x�^�Kh���yL�R+�w��H�'ܑ4�nj6�����'��{��^�r"-�A�K�xy���it���(�?e��^x`���W�ѩ̇�9$������8cq�<�М�������:�iл����F���7������
�������¼��O}s�&��N�!y��Zᴑ��7E���/�n?A�J�����ja�_��y����3��n�GV� &���i�q��ޏ}�6�%�o!�*��Mj߯��]˝,h���9G�}Y<̨�^��T%�>��w���ؿClZ��pB�	s�s'�׺���>��p���SΒ����������%����ʜs�c�U�u����*��|H1�Q�p�t��墾�Vo�y��8ݦA�$ȓ��F%ԓ�gq֤�)�Ya%�Ɏ�Y�������׻y]�_V����6Lzqے����)����LA�Ua��J8�U_ٙ�F�,%��5�',W�^t�QƩjy.˲|(-�z��L�Qk���Ä��/�w�Vn�;�m-�:|�t���)Eq6n3v�z���1n�S�g���ng��->+�p���;+�5�N�mB���y����{Ԥͯ*��H���莌�OR85�@�� ���?p<�>>�o��㪏�h�&������	k�T�Ѿ����_^0=�w,u�����;>)p�a	Y�W�*�EH>���>t���xA��%���j|�������c���<bq��a޷��n9M�W$N�����s46w�y�WС��7�um֍2dKtM�������2��M��JP���h��^��(�˴�2a���]��[�A|�8�R��m����c� h�9�,2��)#"����V��idTqz�OG`��'h����*��$�5��}&���Ƅ��pvj�GKRP�?\�v��p�yjSuճ�S�\q��
d"N��Yd�j%�SL�2�$A�)Ȭ ��j��c��E�s���7��	����֎ו(?���j���y��~~�}'��I=��=��%l�z��<��)���\V)T�I�m�&�yu�6	�����F6�׬��_(���91+��Q���O�4{#$��D)��q�|�)ѽ2W�tz��u ��굶ڽ�5~����bi���_  ��s��[u��0����������pۑ
'�ͅ��"����etV�N�X���89�h��O&TkW}W�j�5�q��1�G��OOW-�����p+gz�z��Ó/^�C���鹁W_���R�56�V7w$�C��,��jw��
!%uɣU��w7]��Tdy7v�����NQ`�I��J�Q�F�A�z�Ў��&Ӛ���V���ͻ-A��1���{8P����ӕ�J���y�a����V��s�9�\��A�"�{�e_/�����#iz���BK��(�d�2�U�B�Lw�wt������t�Z�R�����'��Џ�Į���WGq�0�{dG>|�(���1g�ӓ�
�|�Gc�;{&ęlo�df�LJ]͜���@�yML���6�\����[Sd�Z1ێ���:Ơʏɯ�I�Pg�h�)QN�#^]蟖���f��z��\�)�M��8����g����ـ���j�K���$u}Xq�5C��e�~��ʻ����F]��AK�Ú�������rt�%�돍>���+ɿ�Z�U���Jg��;�ݚn���r�Kxu�Z=�u���m��_<|�_+��-���W�..�GlY��؁�Rd��X�l��?�����%%�;�j��9���R�6}�KB1���}v�{������G��8W�*�kG�������nn2�ytw���Ln׈�[�ú����ZS�<s�u��'�/���먕F�+}�)�����6���Z츘�o<�/�@�(+)D��1�@�>t;p:ȱ�k ��N����,�Tf���yf-,�ޯn5���w�z�>�8��J���h�(��^��5Y����b��]<����+=�Q�vOk��I��`�aY�tgk�����n��A�m�;�c��~v�z�k3�D�o��(H�F��n����z�:�u�v��I�B��ME��|'�]7��Pws�a�X��)�
�	��k>S�a*g�|M���n�7��'��z��>5�8��^�bn�\�{�&�7V!��V��Ok���6U��7B�{�:����Ci�y������m,�[��W��ZQd;�YK��� �V�7v���� ��z��3�c�"ԝPM�}j��k6G�Wm�@4� Yb����<F��J���C��B�]#Ԉ��� ]+�^NP7*+���}fue�%
qH����7EL�$5#����C�$����y)w&GW�]9Y~��+I��ҹJ�H�J��{�7�w���\�+c�!9�=�.��:.|(��{�����6)�::�S;_.���~�{0OP�[�&f�䉎�u��)b7澣Dx��_c�t�'�;�g�9�5�9R�c|�t�z�Mu���olԐ�"�L�o^LM�kF�
�|M��^u*�t�$�A�:o~����q��_���{>��O��WI��P3>g�rg#�x�ul'���ɚQ1�$#M.��B)�m��l�es�/J��W��Q�{.���K����{'Ts�Rim�U�y6���=��L������<1�,M�"F{5�oˍ��.�T�3���_Vђon��\�.�|�j�mC�Ck+vl&$x�=E��w�Eg�W|���u��76;�}��1Œ|��őڶ�f>�u��dS��r#�P��_���Լ��.�9	0D�D|j�@2v�@�<����mkO���������.�u�{��̄)$]�n���o����:,����⌣H�Qy��1*_6�(Ch�Qe� -̹� 1��r��o��2��g~{ڴ�����3�{��a�(��U�}��*ޒ��m:�F��",��O�_f���ξ��N��o�{�E���5�>K.7�T�	Q��`�|k���u5FZ�G,�鞟N�򶄉X7�J�
`tR%�uq�x1N��q���:J�Y�=���~��|MK-���)Q��{�ܥkM�#w��pEYQG��R����[�4�Vw�=<�UدM�]��V�kphS�o�)8bSV1Co;�+�C���泠k���=����6�"�K�FE�*������z�]��S�d��8M�h�N���Q��7L��<���]K���p�%�9�����w=�.HB��s�i`Y�D��� ��R
ozk�z�͚U��] �?�t-!�c��Vz��{a�d�T���+ߵ.������br�t������]��a�֞O�����	ͅ�:�O4{(�-�*Sn�WA���s���5�������a���v��w@v�Y��\$l��i����'S�M=Dj��y|�+���`{d�i�&����q&�Nt���o�� �hQ�t���;p<�9��R+o��F8;ž��`����u0��@v	#�4��hB(BBL�7<5�Tr�d� ��<�o&�2W�F�8X�e�VYZ�x2'YI�~�L\m��w��c��Ww>���~�Hm�(͵��$T���a�g�׋;�[+U��NM�\�����˄������환�v��{[���E�K`6Pp�~�#:��[+$@{A;QCǺ\�f;�(��ˣS����83t��#'_��ߤ]��\��n�pj_Z�eW�y�W��%��Lz��~v6�q4��u/D��]Zs��4���"=�Y��>�([>걠�F�B��	ݧUJg=��q����(���^C�'�B|Ww�rn^Ř٬������Z)�"���ɽM��HM��7Y,vK��(��/ku+v�evz�x� L��.�MbyTy���E,��)O��p)dy!/�#�Ap�Mv:���*��SM�OJ�e�LF�$ �J.G��&c杣VH*/6]�
��$�������U�(�^u��_ek.C�֖�*��! c�jrZ�V�Tf2"[d�%غ�M�4 �5N�fV8L=����?!+���j,)�f��D_&��UEM��c�Ӣ��6�݆�w	N�t�@�^{T����Ļa�8�-l��������ۛ�Q'��H+����M�ϲs�V"�������\,���jfQ�j�w�(��e(��U�qtϝGK�;���	M��w��Y�-�^�i�Z�Ǝ�ǚÊ�9�����Fp�p�G����%�����X��������#� ���%�Mҷ:�/پ,�\e��>�M$]�5H�ȭ}���L���?@=�kY�ײ��1��%�����I��(m��U�֋����%Uo9A���r�]��i��5��µ{J�i����vʖA��M X�FL�����S��k�@�o��W�,T=�_����l�K����Zjpk��H��D[Zہ�M��p���+�[{^��x��R>$�^ȯ?屿l!�󝸔�~��@ʞPC��a#�����X��WT!��P�.͑Q��{��!��$�)�� Y.e���w�`��vk�o2w��g�kܿ��Ҹ�?��| �+ �GH��#r,^��!>*��d�Y�;!l:�{8�,3;�iT���a��s��d�LFy�c�9���m�{�{�c���L5t��N]�*]����'�J4�����ș҈���F�Ԍ�kV�/�; �z�Ա�3�:)S�~���5���j�j=�g���гi��p����OvS����Sq!�ZP��te�6c�uW������o��w�*�� F��(���#�k�56[��ݤ��ávj����B+&�it�.�︡ՓL����"&&�Q��+<�������;!U �������C�j�k��-��:H% 3�}���&�^x������c,�G�Wӎ�pD;�%����R����f-v�Q�4\'U+��]��=��d��_]U���c(POD�u��$�:�t���$ώ�����Uj��x�,���" ����R��j�E��>Q48�Ǽۤ��dE�b����s$C�x�`Y����9��7MH<��wD�j���55;�P��,CPXB�r�	UZ _%���Q�,r�ɮ��}�i������e�a�~�-�O�����K���*o�/o��w�d�ki��Uc�sI��t]s�o�W�d/yܸ����e�F1͹>�����3M%��L�W��n�⍄������1��p� l]X��O�5K��B����VY��m��벺���^e���ֈ��70�>�z�C���ʃ��q�����OWKe�L;炼�{�E�]j����r��een1��,�3)D�y��0�ʍ��0]��>��so H�FY�2)�(�Y��CD���J��D���IoL���c6\#�����������}��އv�~_�G���S�ǌ)��/|,_�rq�Ӟ�8��]�9#"4��~� �m�9���`W��w㧽٢��gK��e����^E��߷��k���6�{������+iN�k�E�mu5�U�Sl�i�������[3X��bֿ7��^�d%��0��"�uMa��<�Tyu��Fݽ�O�v��Eg�PZ������N�?���^�;�_�B3�Um*b��))�ܔ���תn��)�߇�e�$!>u|�[�h�t�8��������A�nԢ�/�\ t������t��,|G�˄/� }3���b����>XC7K�Р�ͺ>��1��l�����(�=� Q�q">���b]��r����c�y`Ę���]o���=}�����Q���9��!�G��9�u��4]���yd`u�Aŉ܍} �噫X�q���do���Ɋ>����6;������wv��l_����re~��ٔW�'1�^G3��0�mC+��է&Q���;OґQ3N�5>�qBE��Z�6\����h��(��n�e�ȵE�o{z�'�4"�ߺ;��U�a5�_1�LP�>":�̮���l+��{�h���җ�D���U ���� �� �"s�ӆ�|�q�!��%U<�XJ��e���k��
����+�6�Ė'��m��]_H�>M�ޤ�r�^>-�pv�?�h��?_50�f�����q!]�8s����A~����g5rO�EA=>����F[�t8�C!#u�:���lk�D"j�ېˈ��5�/|�`�־�z��w��v��r���M(��𛜑��[u�9A��2�v��k������H[^�P����;��:��[<^#�?�� �P�(UU��
U_���*����B� (U�*���@�j� (TT*��F�P&���EP@P��(
� ���
g�߀@P����� *��UU�UB��UU�������� UB�����_��/������ @P�� 
 P�C�5U@ ��O�� ��UWX�/W�ʪ
���G�?����UP�(UU_���T
�� UB����T
���0P*����b���k���@P���z��B�������UB��UU��T(
U_C�p��wP_玪�B���?������ *��UU��DT
�������PVI��f��H��>�` �����������V�Q*",m"*�*UH�JUJ(�*�j��J��m��V�BP[jT[j��6�֨���ERH��R6ª
J�� *"��l�تR��JJ�U/cQUR��$������QR
�*JV�JQJ���&�U�EH�6��TL�TK`4@��G-�B��5;-��뫵)Z�UDSn�;�����lj�Ϊր%�6h��wvUj��-�"vΫ�iUI
]eF��5�;v�J	+l�J!H�DBT�    �`     f��\v�V��K�s]uv��e,�k�UU�ܺ���C�U�ݧn�$��@��t��&)�*w6��v�%M�v��D)H����APP�wvf%ܮ�U��]c��ٳ�[ie]7U�Ƶ��SlF�k��d�ح��V�Wvu���t�F����u��-k��i���dj����[:]ҠH��P�5�UfRUSR�E��e.�Yngm�����ٳ��̮�W9��nZ�qR�cu����W3vu�)jM4�L����L���j���ZV�VU��IhLDB��L��b	J����:*��!��@��P�A�f��aN���K3nṍX8�h�f�FXt 2� (�SR�4+iV4T��*�	��UQ��*�m����h*����l P֮�8 A�&4�F�LӷtKY��պ����;����B��j�k:�r�B��I��R���DMj��1;l�6�Զ#Zƶ��X4��Ь �6#�MKFd��B�:S���kSXiem���X�6�6H�44
�n��J�%CM��Jhj;Y�*6͊m�V ��kl�M�f�hPm��NvR2cCm�A֖��B�h�k�vѬaA�h20�4�j��ӭTHM�� P�Zē����t� `�ҘW@�E�N���h����Q��F�;�YM(V[����k&�t�]�� t�r�m��졁Ti@��$�UH�CH ��i��QT���۳�ѩ�N����et��.u�wv��A�W'G;m����;����jj��N�G9,�9-�)D��,t ���: ��G@Pv:�w      O��*Ph�"��I)R�F �1�1F�  "�� ��Pb1�4�2  i�	)M(� x�B�����"hK VG��f �dr�A��'���9�����+�ι�4y���� ����� @���� �D@�@ ��� ��@ �b  ����������2�$��DL��V��#�*a�Yy�QZ4�]��0Ac�ad���b�ǖi-wvj�FM⥔]�Ԇ<�L�r�n�b
�h;��]�-G�0Ĥ�G��� ���LT�[F"��)n]�fe9왆<���ڼ*�v��e���������7^�
&Q�z1!2��ݏr�d.�����]	z2�r�~�jo2��Y��ʮ�� ��ٶ 1UW
�X��ga ����QY�7b��IT����jSB6����*b���	]�����7�d�Z�úh@R�Y+S�b�Ma�:"�*U�M�z���G��ѯԦ_��͛Q X�Rc�m�0n���� dղ&�5�a��/AU��5�]��Y�Ske��x+8��W(
;3�(N�MY������e���t�$�+!��-My��X��
5�!E����n��h1N%̈Qز���&����"��N�,��[B<�V��Fo5  ��rZ���E�wk4�t�iB2棬�L��yq*�jD�UA���' �/HQU�C!���O+jP�]Ź�RT�h���3hzF�`�R���hn�	��2f�G�2�u�<g�H�W0�2� VYNU�OU��bYY�Y��n��v�h� �F�ۊ�i�
�g"�_�G-�ÏFk��n��m�i�u�aH^��t�����V�f��3NZ�
yP����`��Z�8���8@9v��:tnR�P����(5��RieX�Jd�BYd�@�ˍ��v�$�D��+L�	Pt�Ǣ�QW[�h3N�(Z%j�M=�SɃ0���7:���&h�-.w:��\x.~����r��5��
t�ɪ�$T��+7(T�Mc��3��tɷ����
�����[�N��c�kj��%;�� Է
�u5�[�Yo`ec6r��x/�$��V�]��	�T.��J���P%�-p�ᎴfYU��DGu�$��D"i�kU)xA�}B����wZn��fN�(Mu�1 4� *��1E�:�`Y�RU�H���)�~�]�[2�1�xf�KZ�b`Wycwlj��M8��7R*� �ȋ@P�Xv��ձ6V#�BT21�n���Q	��Yح�[��VH���z*6om5������^�.��h��V�;Y6�9{BZ���n�[a��YS!��Qv���=�*hv��!�7$����1l9����6+Y�&�V�Y�:�m�L�PAwvF��O��km�DҜ��;�+�ڝ�U���*B��#��6�WO][��]m��F�j������*�� #.��Y�(��j'v�4f��e�usVH�`I�t��s�
�p��tj�f��.@��+m�n�M�5d�!3?����z���*eJ�j��}jR�&0��5��F���G��&�����l�E[�V���2D1�9�$�� �bB��F��&S6^�e3���1�j�o2��ʄ��R=Grl� ��u6�z�D�޹Z�{r��8��)�H���7M���K�2�����=�����t,h��V��jc�˭��.ՀCvMA�����Xd�½rk"��C�oJ	�C.��cǲ Q��/U��V�G2��x������(���g +NRf��&�H�f;�;/qG6M�j�u ��{f�mKT�X�תb����7���Nk)YP�;��Ep��'dʷ�Z��ڴ�t���l�є-��\�WU����的�8���ݱ��&:hl�ݡd�ڽu6^X4n!�4�쨦ȤD��4��2�m3�j��(7A���{M5�J�U�m�Wm���qطS%ڂ�/ƍLCяh+�Ee��o%�[K.���-E�QX	9�P��Ð�(0i����VK�X������W/#�2���B�n���,]H����LKY{6�'�Pb(�i�(�W�t�Yh^��]`Su�6�]X(���ᥢQ~U��/eM4.R��;� 5��(n��X�x��2`L��Ra�D�Sy�X)8�&����흶Xv*� 
A �=@��۬�V�,LM6l*�B�Ȟ��ܬ��f�M$�)˻���ni��lt&�gM]IF�[ki�7Sh�D((RR^7�Qԩ֧�Bh�3i�{��r[Xsk2�nFfC�f��n�Q���ct��L���oHݓe,��v I��![QSc*ōA^j�F��0V2�F��Q��z�o%�:�*�t��ŚB��I�㩁���ʻH�,��W����l���e�ڂ�q�.n��1�d�J�縄��;Wa��ֈ�$� 6�Ԣbo噫 #�,�����0#����h�;ڂ�Odя.���ԗ��j��l䳚ݬP������њ)�#H�-S�"�ԻՏNSͩt�t�&�OF^Zi�uZ�ݧ=L��dݏ�&�L8��l����9�1%�N˱�rK��m�V$Z�8�u]GI��-K 2���c���"
�}3r^����4pA�����.')�`yGr�on[���Opޱ�:��R�f'NErԧKY��]Ӏ����ͭ����36쇪TV���j4����#�g ;*d|�r�:�9����g䯍<`���i��+[�d�$;)�o1\uu��An[;��63w['��.�U�«.�b���u97w�5V�T��N�1��d�@  r�X�Y��Hw:��N�A���a���E��9x�R�Ŗ�K��PgwUT��|���c��ͩ[&�[�^˳j*tf�ő�Ul"�[Q@����I��{t�"=S17k�na.;*f�n��f��(��ѥ��F�Z��Y�i#���-�Ǐo7�c���	5V�1cQX��3�� �r��T�v�7W�[��F�jejy(��oE�Z�l,��nK̟�2+[SN�Aܑ;{�*��y�+[����6+�Yz�t�{���(m�@\/�D��hĔ�x�uh�÷5�2�I���4���W�᭶ ����t6��8��-K�fm��86�"qB>�tv�Φl<țw�nB1��&D
�s5�rދ2�[jC& Bi![�(;�I@ݭ�����)�]�iM���m�u%��2�m��-1��q#��[��L�54���;������Mrݪ<�۽́�[%���K1�J�rnXz���+`ɶ��u�Ij�fˎd
M�&c׻�OՋ�i�1N��3&���jɳ.1�T5"a�a�o?]Ʉn�����՚hL;H@Y5x��6� �����jM'bTU���.�7��^�\�Q?���Hͷ4fn�ȦTn� Rhn�^Ŧ)��L��i踎Ė�#�T���h6[6�̢�I�iw�����%��i�w6R�k�(aIջۼ�7N�4O�/�J?�hkF$�ٺ�q]#	� Xķ��ʊ��8��"��V�!��Z�2!_�2��"惐�,T�0��f��,kM���ZMKEmmcn�⼼i�v�4(���ۡ�	��Ų+p��mG%m^˳R�;�5֝�l�&�d~��K,b���1�N;��V��M�&i�̭��o@ʚ�ʎP�r�\Q��c.V���T0�`��6�+e4n�]k��P�1��K��@��1�3�[N ӝ�Z������ٶ����N���WO&f�C5Z��C��t0�8(5��N�wX��ûF[P�5Q�"��e=xXtՒ�N��x��a�X7+ �-֌�b����WZ	l�9�5c�� V��,d��+�2 QD���2�J�i1�Ot^�r�ެ��#��!Fo^� �P�4�Ũ��Ec�n$�mV8��ù�K��̔�Z���!��NÊ�:4�2~z.��0�4;�dĴ���:k0���ՠ��&;�[�5��s!�V?8�ԼDœf�a���Ú��f�%f%6�\ذ�N�
��������\'
��h5O	%�BK���l�+%�3h���M�^,4�Gv� 6��#aG�ha�o��ہZ�X�36�1f���T��V�Xh$��]mʺA� � �2Uf��%m�����dlY���B
21�ճo
%�� ��� +#���4]��%Tɸ�9�aT���))Fė���:�e�[f�w^`̤�ѻ�^Fj���I'�g� ��Տ�������(*P�7���$�Ă����h�ᰡ���8Ŵ#$�F�%�Y�[ݵ�P�pY�Zf���Fp2�2�8�3uz�fh�FAUK�2�ƍX�`V4ɡ��u��n���(?
t�w�n�/�:H9��Bwe�8�<u,��ۼ�A=&�bF]3H�� ����P�dh�,"�̂
%�ڡ�⎢OQK�Tխ���)f�P�)�n����4j����⥉83j�;1jz7;�q�OU�"�: �	�K9�I�j�hbJb��E$,J�F1*b�*m�f�eٻaB������Kݩj�Rf����dB�ku`f�*$5-�
�*�.l���M���:SRLn3��N�a�&�,���������c�I��3o4���MȮ�n�h�!U������6�7&��^���Yo)*����2��o��	\��M��,��;^�	B��� ʗ��D�j�Ր=��i���i�M�3a2�l�Y���/EiuS��-ͫz�!bZ�e^��Ƀ�L��&�voU;���5�h5,.�J��dX��H�;����[e�6��͸��D2op�ݥb��\p��&�Gn�u��b���,(0J֮X�R8&�`��V�H�ёT.��E�d�YR�k�@�g2��b�h���[(~��1V�م[ulӣ�۷��[�n1Q����BeJ���U�u%m�SeͧX�v��Ҡ�`2��X.�#'�+7���ؖ<�ZaH�w�
P��Fe ڇ(������O�
��Cf�Dof(��F��X����@2����m<6�-��k �Wt��	�/ ]�����f�-�wX�@�x��\������^�٦E�p�Û2w0���8�b��[�o�Bؖ/ws����i�w�wsr�@%F��Д���<tM�6��OfR,�����%:	[iM �a��cBɹSNP�!0Y$ލ;YP��nֆ�X� mZq�r���ӬUlʒ�˷0GVA�z&����F��ik�gD�����TY`&T��̬h�0�vM�R�今I�z�+��^��Siބ����?,�7K1Sbh�@5�a�1�a�Rm'@�wrk�˴�+B��e(r�Чt�Q�;2�n�ei��YN�^���Ͱv,i�Ma�����P���(��$"����,cFV��t��!&n�]ˑZU5n�֑�)�Ǐٷ���fhf����KL�B)j^���M�3)4��-V�I]�kM�{g4~3Mx�\��7�S��d�����S�H9;�G�s�Ћ �P�W'�R�^	�a"E�me���U˫���!���i�9o0=��0�=�:���:"������O����m(e�2�ڻ��`V�I���2�ŋ���j�g�����M����F�Aod/mV�
���j��ٿ�7�AWX�*4��r�Ȼ�gk#�V�u��Mn8�5���fA��z�\f~Z�O�T涵��5	R<�c/3j�]n�mB�k!�M6l˚4�BP�K�
�t���vmd�eA��۫�R[�ź��k %�[ȿ,xYL�kcx�Wn�㡅�-]�H]��N��˴��S��t"i���cw-��!�ȯn~ԂD���KpL���+^݅G���(��sq�N���+v5��<+��qec��kM��t�:�����:���`��l��_�!���B �Q[
��� ���(�/�A�rG� ��e��{C]!�Y���p�H��:�-�O%��s�4�]��$����/[���(�Z�k83V���J��2a���/m�)[E@��K��srZ6D�2�ͬ���a�18�M{����c1��ѵ�����P[Xaӎ��Z�r� �e�{�Kjd�2��*^��i���H1��ysl�^MNݝ@��t��p�������Qr���:7�e3R��������Yx��X޶i�ŋ�y��̻�>�rf������x͚��ZZ[��iWb��j�D*W�B�`�i� Ն�B��[���
AfeB�ؐ6�U��w�pإI�4ʷ�j�A�.J+fU�Qm�6Ԑm����r��ʜ���n��1���O]`�M$��0����35�w���U��2Ԁ�i�z-RS?,� ݱJ��弔+p� �x� �Hb5�j�W!�u6�7WP�+s7�A������5ghK�\�2K)�W&Yj�m��V��ӹ��#?KX���~W6�u4���)�B�G@%��&L7�e�Q��[�׎\�X,�a�D�{2��T�X51ͩ�eމa�ԙ��ǒ�=2@����w���f5b���Q:����ܶ/o$c�Uj�o�X6�
�-V��ve��4��uأr�f+����sXݭ-�h
a�t�,ۥ���e�� 'N�*~B�[�9�.��E��,RZ�%X�7)�X0�v���EGS�Q��Mj��R�4���q��B�;t�10�ku�~EMd,���s"4`��h����[����uk��T0a�I��WF�f��wu���D;[L��xͭٮ�h����a� -��尋T.���0^��KRĻ�	x���Y4v� ��ު��[�5e���N�7� w.
+�
(iw�ս ��m���u�:{~j��͗1Ţ����rOڛ�����{��J��a�i�FV8�v�T�#�z5�@��B҅Z���? ���-
��n����YR�`������Lj!�u�?m]��O$��L���[�7/o(c����'�d����#}v�o��;������67�t�̛9�$\�k�H�I�#}�p��oz8�\�nI����K/�J$��KZ��p�mvv���F�H�I#�$����\�1��Ѿ�7�F�IF���aS'��(�Fҙ����1v����,����|�]�����䑾,2n��I:7���;�}ӻ�г{^��ʎ���5�MczC�JM#8�����̚��6bC#.8ww/jgQ��eGoVb�M��i���Ô�sU�#��kZ��]^�S�˭�����GE�hd��8neo+�֍�	����]�j X-�F�.K!��-��{@���@�*ޤ_���8Hr0"����[��;!��:k[d-�9м����ݴf�n�v��ޑ���Ю��a�X���jt⁔�4�#:����K��� [�C�T������qˎb�sD�D=%cyU�7�]����;W^rڑst�<&�Q�8��0��6��д���5}AXVNL��G���u|�j���u���2��R�,J��=�I�B�b] Β���
�x��z���i�B���F�u�Du�;tcA��n��]��ZK�ߕԣs�
E2�e���a��Y�����G�aM�S�u9�m���ʛ[�,��v�w� ��۬6��3.���Ç9�iD�0]�y]���㈀�*M�ւ���_X7p+P�34�Ӽ���*}�R� |��l*xxD��	��
ݱf`�KҲQ��Cv_� �c�b�{	�3�䷗rג�O6�2v!��\�b�IK���;aŖ��皱V>&��=$4�p��e�����W����X�U)�m�Y:����9���rʭ��ꥎoB��/WsKH���f���:��G���^�SK�����TC�wV�;:�������dA�V�z�gl-q��,5%L���D�swm݇��c�����0*�wj�ظĔe��n�Z��_�E-	��~u�l,{֬���%)2o��LT����∼fփD~��o��M�aV���j��n��\Z*:����a�-�J��F밋��C;��ޤ�f[cx(�v��E����s7YN��B[��dJ��ܗ��wC�%v��cb-'x�X�qܫ��
KBt��4�Y�m؉�ݛai*e�

w�"G_d�����Ǜ����C]+B4�5
���̶ZG��	2���ri��!��U�r���(���;ӫwz��},���vH�[�|v]m�G|��r!ԑ�j�C���a�tV�fK��i,��)0N^ڛ�E��&�Օ���9�0>�.��JG�D"7��4�Lu�[�fp�e�c�v=ɡP�H�7X�,���=.\�z�ciڬ#�QC3Z�p6��1T[LfV�[��S1�qZ۪�-'����1e;5�=RܖFqx�6��z��K�����p>��L<�� л��u�;
ܴ����
���6U��DX���V�iIvU�G#t)]B�̍�� {�+��]�;��k�q�3/7R<�),S�
ٛ\K�W�"�d��փRG|e�èlLJ�k)4.�h���+73ky�3�zD�"�/)~�l
���8��X��7�����/rŹB��.f�y��w}��it'�n=ͧ���V�PR?�F�]���g[ͭ�|X2����@�Ӕ����{��{4u-�Js,((J��c!sS]��S��^*�KW��c��lxXLxz�'��Wb�����w�Dd�K�Xnh��r�K���['r�:B���R���X��c+��| �y.4�m���v�5{ʮ;�2�M��X�D�EawVJ
�-Ŝg~�qG�˽/I�������v
��Š��ȲmИbȲ��>K��=�׫4���� �fM������]�޳+,���{��։Re֗\erwB�o��0-���j�6��o��Y��S�_]���� �5�Dg���I��e\�Ιԍn�1�s@k�I���g*Sj��vW
�:�J�hÑ�����D�,_k�����E���THbz�~�����V��f@f!�*���&���v�(��l^�3�-��v
}�%�ka.��S�aU.�t%���=z��<��p>��Ƣ�q��e�](�(l ��W���0Sp˛�Z�ԁ@l��bP[�xs��5
��x]��A��F
�(K�TU��=2�`�Q�E�XT�B��r4�������uȞ�Ɓ�Y����� ����kv��=+fSΧ�PpS5����Bܼ	��떹�o�CG���Ƿ/�N�s6Σ#c4�=��t!����������u1�3�tպ������Ue��g9����c����M��Sn�Y�f8�4d�3�;g6�t�Ⱆv�t�g%�^�8���]3�0��7KP��ԣ[�fn��V�Ds�F=��u�����&췳6�2�]We����Pu,�jMs2���Qe�S+7Xh��p��Ʀ澭M�{�m;�rB�O3.�_U�P
�U�iҴ��
��ibhʒ���9t�o��[ٜ������NeuF��1bIi ؼ�Z��Ƌ)ĝ��'�z�P�E�\�ݰ#8�f��啚�Nn��*Y�w�G��.�y$���j�S8�:���p]#ͫ���p�q��v��`�`���1d�&˄R"j�U���7lke)U�o�ܸ��,��U���u6!�#���E8�{�Y�=ћ�a�,|Z�J�W�(��.�`k��:DP�:�:����`��͝c3��*>ۭ{W[�۵���c�\�b��'��6���;c�X�J3$p�$F��;��]����;��#�|k%8J��2K�>^�X�3�'����ך
�6M�W8jQ�k6R4��/�N�W�D��/C�[7���4N�01����r���</#��
�p����:��Z����d��Zvw��c[fm��[L0C2���)��ż��#o�Ú��2.e����gkaⲴPHe]A������ZtѶ̊͟Z�cY�p��@��ZwE�J��AIqS��T�o�u�h���GI�]�E�*�<k��L�C�>[��bgR����7��������B�C}F�n�ֈ6��;U����;���	i�Wc�TJ�.������kC� �IqG�Y�f'gk�*W��2�t�)���c��G�?З���EL��%]C���d�e��B�v�%2�U�x35��L�![OY�̱p��5����c8n�lg�<���+��a���;,j҃�zLT�C�t��]����RVh�-oC�y�<��ڼ@7�A�HQ'��w8��6���&NPU����<�]R�[�!�f�3&���+�O�T�"ɷ˶��d�xD����c�q�[�O ���2������������-��BJ6w�ڭ�F�a���2�c%=���W��i�ē�=iN5��;����TXf��<%AY��/6�c�'�R84KV�F*��0����n�Vl����}�n���U�w���Jdg��a�Y��b�>��]���8]m�P���ã��CkЦ��-�km9'GQ�wq5kX�������9Qe
a�Tc3}�2����A6z� ǫ �j�md��t�2������]K���D�(�l���V#��uZ����^��y��0�&>:��ް�����R�Ҥl�w.�N]_%4�R4e7�g�8�,'5۬n�D��ZN���P����iV�p�=St%W���R��3&��0
�Uak��*�#K3�ˏ��tD捊��Ӈ�H��pS�S�������5����|M����q��mَS^�V����Jn'�c��r�g󧌃J�7ɽ��0c�L���k.:ÌR�N��:�Z� �twIl���Q>�f:7a�] �B��	Jۢ���������wp۹	�s�E��9j�r���k�70J+�ܓ8>G��@z��ɒ�=]�%Rb��n���>:S��G�f�7��Ky�Y,p�9�ٹ�-g��f˘��	A�t{�t�SwÂ�#C�uu��u��@;H3qMR���t��LL$����D,�N#�&5,�nﺹP����+/�̻ʇ*��JC��革��d�"�e��3�Ҿ�ظ�ڪ�B"�x�u�7�-Qn�.�H�䣻¯�;����G��.� E"&;ԯin]���9�B9�T3��~]_t�כ�3b9N��,��m+=b�ڒu��qa\v��E����R��LQ�Ν��i	��r���k�w�\�\P�B���0���@�$�'�nے�8�`��}����`�GG.�[.��ζ��U��Խ�(�/3e�V�l�{�=��y�T� A,�Y|r+Fd���2�J�'X	rש]��#�}6WU�b�q&K�
�ޢ����wjy]�ӊGj�F�As�G<�X��nA�f���Aͅ#��1|V�9V.���=��	=/n���G�F��Q���`�u�}lѾº�A��h��8Tr�'v�\Fr�'Wk���x�����d��!�v�_T���}b�;�����t�[t:��X�H)��1]�� ���,'��Ѵ�挔ܳ(�6-e��]�&sі:$��V�̎6�&�ѳ��V�̵E�B���p���'[�:����R�3y�i��hm�{7Fz�h=���5o��0��{��H�E���g[�}Y���Us��6�i޽\���Y�l�V�9&����v:��!۶f��|5�����2�c(�=7
�� ۘt	Օ��i]a5̻����PR�+��]��J:�R��]��B�ɩ��N�\�7�M�G9.n:2��ӧ�'E�;o9���Pn�8&��S&.Y�rW~��T��}D�tbT�,��J�30�*("�ܗ�V���>V]��Ռ����W,�2�]�zlA���OhL.
2*O�ٱ1�2��ހ�̹bB�;@�!y�,�L��nh�T!Oj凵�=�t �I{������xl��zb��,f���́��*0x���"��w[���BN	u�;�9[%�B5bKsB��C�^�@�p���7CX�P�Od�R\o��]f��ݤz��*�al8����z��f���]߶1�KVb;��ܩZ�D��zYӆ���ya�G�;�4��$<��\ܕ������Փr��;&���)�*�i���&AG��q[W3 eҵ�d�Gv��(��Q�&��c+�re=wM�6��\��yvs�M�K�v���q��Җ`xFq'Z)���4:�L���E{�-f�EJ��a�]��ʧM�j�;�)qg`g���t�CG�oPЙ����������i�Ǟf�2���z��zl
�a�t�s<��	�
T֮"-EFV�_��n;/��y:X�R:ӎ��û;��눨�z��0۫|�F�les�3��A����%�5�Q{/ii�ὔ�;PT}RA%���C�2I��uں$���*^��aZ��N�[ ~$�:%��o�$8�\��/�o.p��BWBI�w4���]���/nL��i��v�P��1T�*Gz���}�r[�����+O��p�7��(s�x��Y�WMUƶ��هa�RS�������Fz=���Y[���+;�	bs"�`�a:�k��pI�t��v٥sK��Uɔa��G[�z��􆲱I{� �B,���Nto/{n�_n��#��a-IN�/�uw@&ˮ.�Vg{UKB��Y�S�A��GZ�_�#��D^��S#6�y�Ƚ�7M�~tK��R��#�ӹE[���[�,㓎�}Tn��:�p�l�3d�b��p���}f����
v�`��=|�]�nֈ��b���T�a�aF� 9ًr�@��*�F�!YI�>�z�e_\�7l1ۢ���SmZ\.!���N��H�ң*֞��I�'2��ճ��M��qb_��̭V�8�� ���k��K;ٗ'�AL�ɝ�p�-Xdm����h�뎲%B��[#�Ys7l��*s&�9g[�,[VkV�S8�2��y{1R2<hZ��W)[0+jAF�����٢^�VJ�1\�̏�J��������{����d��^8=���W���)
�
Gju��䷞��G� s�+ݝ@̺��)��}����J��f��yW|�i^�.�T��4E�X� l���
XF�n$�v �;�2lb�29�ڞ�t&��ӻge˛�����Wq\2Bns�Ώ
u�g��/�r��iN���[nPgPGp��͚�vwq<�����3�#�7+:��f=�L�8:��B;���X!����C�*t8r���N}�6��ir������� ��h�5t��[J�X=݃Q�z�L����Z���_�>�B�jt=BVKY<`�v+w����m�Gm�%��E*gu���c ���mth�7�U+�q�[�181��N�L�p�.�.�vZ�4��;-`���V���ȻK�[�M�8�0����K�N�ۼ ���0�m�xx�c�سA#�T�[��e�&�ӏ+w �����#ޚ'2!���+/9&@�딛�?��S�ߏ�٢�$����#���+:<�� u�YOEqX6�9��b9��ԥ��%�{RŒ6�U���&� �|gLs�i�B,�snh�b����̣]5~����l����C���Z�%�wOnK��n�/��nK�7�^G5�hL4�T�*�z6�j����Щv���������VMv���F$*MCn�٫�	d�m%�&�븣�����m�.v���#��v��}�vǙ&���M����t]�̣h��3|i�gS�3��68��J*��x�̄f��Έ���9]RX�u!5g�9SCXS�;���ue����̮���$15|TiL����]֫�Ş�f�k,'�;�u.��{Gf9����"ܴ��&ӾNr�7s�EB�+���R$Ve�a��7{����krQ$����ː���q�z��woy�@���A:�2��#h�'!x+.Tт��Xb��}�Uh�ٶoiGO��pes#+lJ�����*�r�a���w�8+�j�����6��N=+l�ּ�P�q^p��B�]�3vmbK	��V�zʓrp�z;p�M��d.w~�շj���  ��� D"?x ""�� �����3�f^f
�	,��幗3Gc߉s/�e�� ��NB!h�s��h=p�N�փ�v�g\κ�.�i�#��� ��I`��7�p�	���ݬ��Gu���TZW��Hm�aw*5+��E��Վp]���ƑGy�9�voF�G	�w����%0�2���,v,bK�U6"��4�E�	aΧ}f��ݮ�+;F�U;'j�q�Ħ������8�oaqG�]�Ђ��շwy�:'ki��E�F��}&s㇦���Ʀ9]w��3[�gm�m�]JG���6Gsɺ���h�3`���6zfʮ���swne��S�ks�c�䓺�Wa�b]J�6��i�����'/_^abZ�S�1���:Z@��Xxζ:*��۬w}�8I�qY�V:�$<���A��+��ٱ``=�Q���B�b[��꧛aǻ�ŝ��Y����-��Z��f���p��#	���^�ȍ$�v�mWL�֫��Z����̷B��䰭M�^-|���Y87igg赪]�r��Jj���(f���q]$#�u�ۑevE.V�����8w���_��#�˞�s�<���mJ�U��giU�֒���ͼΙ)��(.t)��'� �/&��B}�xI�m�[����~�f-�{��v�]4+ZF�z�z�]��h}���mU�=���]e��<�l<�{�P33#�_P���۷*{��ײo�u��s����ǖ1��[]{���5���B�����p[��/����q����[	� ��a�����U#SL]8ڠє�!�6m[4��;���}�F<V�J��[��+�|v�呢�'Nz냲,���nFd������b�U�`Ӳ���G80���{�݃x�h
s�@�#C��Z�Pe�B�e�y3@y��<�@h�9W��UlQ��(�i����8B{�e������=F��)+޳w)�(�Ď�e:{��$m��m�\jcgk��n}��e ��h�4�ѥ�yt�b���-\x�-4i֗�竌ͻ�oM�O�Yc.4��5��N����z.��=y=ك��<�ء3�t�9�׊�	ؽ�l���=�X,~�M��������?s^��4�wG/���9�u��\�[����B�N[O�c]���4��;fa�"Z���	�y�g���u(�p�d�~�`��u�:�>��V��(�t��4��+|����)��Ͷ�p���c���]/�b�;�t
�e��r�}�x���<���6�m���6|i�̟+�5�&��2���*��b��8��4[ێ=X���Z.����ʷX n�FB����u�m�
YӖdPY**�,ݛn�o�T���F{��A��Ք���Pu�t�4p��;�:Xb�����ʷx�&�z:�шhK�f���ek��,u^�tco��_ ?hT���נ�dlj�������1nE<Z�.��/�<��TƙX���s��V��x�K�c��rf`���N�y��\|������P�N�{����W��6(��y�j�{�៽�����������:�b�T�Ec�ח��+ْΣK���M\J�b�[��i�_��u)��6���L�K��rl�ov�D�ƥ
Q`��C��9y��Z/yg�u��@�$}
�ى;��B�5ڿ'Y7�
��:t��4��<eDi�,��V���y9�᜷򽩮^�x�rRu����|����Y#<`�<4r����
V���z����gb��e�ئ�h�f��C�X�%k����9�s&7��.w�M_wu�s��Yڤ���ztf�,C���'�y���N�`�^jX���,�E������Q(ͯw�����ܸ���z<�,!��
q��.^%Om��q�k8����+����˝Q�R�E���c�D�(K�n�cc�si'm��9�6�{/�5)[*jY|�+���X���'v�K���Xһ].�%��u3�Nݞ�;X.;�������+J*FoLh�)�>�G�o_U�Z��M��Q�,��J(�5֮[�bL׃5�4pЮk��9���V�e�8��F� ����O{;����KgSB���f��㣀�/]L���Ub�t����v��h��N��7�@B�cu��R�Q�6T���T�����y��G���q��~�[��0oVZ�T���3ޠ�Wv�`e��F/8��%G��
54��z�70��,[+r�Qt.Ւ{���n��N$+'覨E�԰�G���F>1S�̾l��n���ȭ�AY�)�[�'9�dp��d�q�!�HR�Yv�
��X�=a�|ⰺ�p1ٕ��q�\��v���Q�b����取���>��l��ʧ{h/��[|+�y��\)�^Y�b�s������=�����2�g����Z��斤	+)�Aa����c�4�
����o=�C˲�8}�?wOk55̒O	�%vW0���Ӣ\8w<i�S���3�s��.�
绸�58l��}��:Ǜ�ck�ݨ�
 wM^�u ����n�4���N�/2`�E��v�P5���o�Kɶe��|ulE�.�y�'B�ۮLk���ُ�4�U�T���};��X�F*��M9��v 1����p�qQ�M�[}�8�m�C��2�x
�S�6j�%��{�������.�=R��Վ�{�uq�̋f��i�Ab���4w�m��9<Y=o6��;-ђ�X��4K/F�'ӻ&�h�P7�x�I=����?m
�>-��pi:�炖�/��3�1n��5wg8:�����R]{�L�PI����w�����B谦¶L{�Cyy�"���"�NZ��kO��3�J��p�#&�x΅9(v����Zq�M�0�*�c�%l��<�ͼ������"E�ka��Z:6��HѾ�׵�.��ăBo(�T����Ŝ];�����,F���ګ4���Bݛ�w��d�xwrʼ�;9�ζ��B�uz���+w��0��=�3k�&s��P��$M0��P��{�滂�x�'�E�f]�w�8�$6�dn�K�<�U���.��+E:G3�K��xJ���f&�&�a����t������mw���[P�^��mG���}K!��i�e��=���.u|���v?=�������pc��d�0�;�[m�e�;��=���^����؎��T��Zn̠U��RDLO!��;�U�YՅd}̕r�O��kj*�k��壢� �9���K�C}ۛh�j6�gHb���B�)��}�j,��O������ ���8wf�υK���\H=$s>��+D����j��<tt��+}�x���VSQ�b���U竀S��������Z�@:���)'����3�u�e���-�8Ef��D��9�t�u��B�q:t�#�m��Cm���:u������t�I��]����t���t@&�|��?`��+RGxJa2�y�S�2�Db���0<��{�ŃPo3��&�;���㲖�W�q���.[�1@6��lq�gvG
�r��*�hmN�[As�|�W��m�e�]���b�����']�_�7t�������۳�v�l@����6��Z4����Yzh+�:6����B,�#f^x�آD�5*�Ś�Wd�L+R�c�U��5�`{4s�dy�6�4ˬ DhwL�Y�#}Z�t�z^vY���9��^�*��_�xq�����V�1m����D�����6g5�\�]��Jw�,�6�1f���z���^eG�6L��
�Ka��I\oFl�s*r��w*��w��A�H�H�e\H��YQA3m`��k ��N;�8vqA7��d!�/[�Zs�I�\���5�!Z:��	�;�(cеa;�tT���[`+�ܺ�z���E��o@��qq� 4���i��_T2�"Z��f�Q��{�%���� .E��[���k׌�����i�=r�u�?��5Qt�h��Y
��-��ś2���&e=��<=��C�6�f��IY��*���}�x�
�S�\�1���A�S�o+s�hث^f���?rq޲�/�_(�q��e�|q]�ť���(1�����U� �g��!�q"��
���oP��ѻgm����T�`�k��A�]��Џ.&����np�B����G��+:6
�*X�]*�*.���C��U��E�!�G�v+��s������^��b�n������2o{{v8d�Z�tX5	n��
��L�0h���	8���{�J`s�][��]٧W�m��7#Y0J��'�y�ג�z%��4���G2��(��8��ˉn�Ǣ0$��x��Y�'S�{��u{܈�}���g�-�t:s�3����~ΑNU{�������Ѵ:����F�|nZ$C0��9Cض�FC��K����G�q#%�$�=�\�2eĆ�ݓ���^�u�tf*=���3�9N��ȡ���oM�4;\��N��TѹN��������}I)�o	ۼ�o)�EÕ��
Y�����n�w�Sp̎�Dt�A\eu�Bu����~ۓ�2&�󛑣�¡�
}�D{�W�X7��yl.�ň,M���=���ef>y;O���u�w}��
�g��ٝ�:����ݙ���8^/)� C���ˡ]�o%>�t� PW�T;z�/�Vk�z&�U��y�\^]-��x~V��5����l�K����	}	x:��-��k~h�Z�3^rw��l�8�p̛�S?��,�d�@�Ҍ��N˵r���׼�TI�%��aL�k�%���Z�@HGP���x��Z�Â��o%�:�4myG�$e��@�ó3�y�����Q��̱�d.��#gt}��eMs�z�\���~��c�6����]�R#�Mo�f#��I· =�i�غ� R�~��ʝ�1����m�ofx�zWinH��䉽�f\s\kIݮu���V��7j[����j  ֽ��N�b��0�ȍN�j��E��Þr�P��a]	���?<��J�*7a�i���ة�����/�������E�Tn�oa�q�>YFH��=ul�N;�-�+�J!��ڳc��r�ͬ&�k�\�#%��Ռz� J(�)�6�z�[�6ܕ߮�]ew��]�=�T�b��]�)=��ң�+�Y4/���R�<�y���	�!X��	���RaVM�23{���U����L�'`ګ5��Z2� ���ba@��5:.p�軇T$Ĵ�Vq�\۫�:�&����NNN����pV#�����L��*��X�S���&��U�f�f�����w�"�}��s)�wHjؤjjĖQ��d�O���olNs0v����6n��U\3���ݟ0`G��<+��U��֒�����Ƨו�	ܗ�����/��Pt�l"t��7��Tf����#��6��
w	�:t]�Y����B�Vs��ܬ<Q�tA�/u���q��{ЯC�Wu��GPŪ��K4�SL\{a�n�vE��6����'�>L��k�sC�i�"�PwN�n����xS�.��������U����l�Ӟ��_�̶��^��a�ݑ�{05%[�ϵ$FD^�k0����%�c�T��׈C�q�9�s�`>O�����`\N��ZWLG�y4`��]9��B�	��7��en�"��uȿ�A�.��!�*:
��L����X�s�A�zlkZ�~D� ^���FR����s;8~���:�{!�k�������������P�R���L���'z+�)p9����۬-�lr�z���P�_hh�`�}�m��<�I�|�����qs���.�9.=m�~�����9���ʾ���N�{@���9vY�,f����T��^�"?<f�a���E�Gz<PN�eth������=ا�����n�[�婨]����tޙ3
=�kwR���oV=pa�h\B�͘$X�<5�l���U>�3=���p�L������%�W.����{]zI����7�$�2�κ���N;]�7;^��?��/z�9�����yf�^�Hv�R�tH�(R�u �׋����M������7��u��th��玬� r��؏��J�T:ۖ� ��ﶖ��:c�U����6;�h;�6ߕ��<�֛|�_��&�Z�q�6:{�u\-eoou�7W��Z�X�6 �*+X�r&J��g�w��G�]�C҃�]�[�EP�Þ\�s��<���vq��=�S�p.�yグV�o�)U�����܇�N'��.^���������s��
��߼ύ0�Gwc���2d�jł����d]A�-�MưutM偋N�Ӳ
�z��C�6kX躰�[�.�Z��y��}a�unn�ws�c��Ұ���PY�z��z9�=&�X'��ۋ9�V��&�,a�`2f\a<��Ԇ#�ﳩ���s��a���נmҵ,��]y���r��9��#p�)���}u���i�1�ܬ$�q��4�}/�3W�y��(���r�ow`}�mƪh�-�u��Ʀ��`�m��ĭ���[^��rBb<gUs�� ����uz.ʼ
Z���i��� ��Ύ�����J0`�t�#��x����W����Z�LeM�Rpᎏ��L����l�F�@+�[y	�r�PHLԔ=���C�N6��`ET�H���@Qd�G�#S�i� ]��t�*�&+I)�����b��VZ�j-dviO��ڍpc�C{SC�.uo����e�x�2(Ä�����^�^���,S/7�D�"7�\B�p3k�o�\
��㲞�7A�����-��J���|F����-ի���LF�o1�p�|��~y\��v��R]�Gctث�R���^�g]�L�3y?X����F3?jG_g��^��j�M�E�I�/�i ��^ݜ��[1��΍S��=�.�rY#�B<���o������=D��V�#m�&��b����c���&�����!]��K!�4�C�"�fm��EF�6�]��F�}��ѣ]buAD9C�cMmNt����x8u��<&gS��+��h�DÅíl�r���,�v%^V�KM�XC�.`�W�'T��U߷4q�^^Z�r�op��	u�B[t�;��]�F�=�ò� �:��H�U�+���JE���Ҧ:�ɜ�N<��k�V$x�u��@�]����-C �ȡESSn>;YN�@+���iea�;\�v�4q�&(ю�� ��r�6|;o1Т��hҼҫRXm���:5e�\3'Zv�u՞�8�C.�j$�O�p�2
�P�.��+,��gt�j-����ۚ�(�1���J���N9�"c�F��c!��o3V2��!��q��7��1���6��m�]�g�bYDv�<�T���k,Æ�ޜ�n�[|�:�v�D��<���
��M�	Z���'z�Pk�nS��,Nw��7E>�S L����-� �������%����Y��t'�=ڏ,��i�ӭp��ء�oAlE,�5�R��y:!e�������ηr�hM���Db��W��=Z��1�6��yD�9}"��5�Ʋ�D�7u�s���l2�[�lnp2KS��d���9��E��"2㼇�j7Y��.LN�ȱ~�1��Hp�|3Z�ur j�C�ZS{p��)�3�a60�u٢�[��Ȭ(B��Μx��Rj��:p(ؐ\[��ޫ���2�ps,%e�b�pf����墷#5��`��;-�Ԭ����F��n�s���)��Nv]�!&m�f�s��������-�:`����En"�J�}V�\�T�e�3ˎ�VvU�딍���\9R�4>�R:��곽���4ǝP+⫠;3�]j��c�ó �u��0��9B���čW?^����h2�n��l�t뱸;�x]]�f6���d�t�ȃۀ	eݑ�hC� ������$��n)�Cxq�+B7B �Z!<A\P�W��Ki.�D[��k��事j�P/p�ܔ#��}�W2�_Һ��GZ��Y]��n�h���Ѕ]bc�`ɼ�����x;�t��.y���@�s�.����Z�̒���b4�iVd�7&7Z���FkƔx�h��o&�k����λ^�jQG_u}{����ؔ`64��*J�wί���u�CȢ� K��O|'T�{k��Q)�u0w-Y�6U/��zT��k(�.=L�V�"�w`��
�҂�/0�K�I���8��na��|��Wsw�g�η� �(��Ȑ*˳v��}v�[�c��Ǎ�Â���'��wA�ŀ�:p�����[=�\	�����rC�w;���*��d���u��4��!�"�k���zV�f��6�!��9�};1c��)f��v�E՝�Ǎ�Gs�����N���������Sh1�!����fS�.�偖�ӧݭ�\�s\}��#e��e!L9�yDNU�����OE�s;�u�`1��}n��m!��nK˛F�� ujj7YSF�E<x뉆�Ų���{q�W�qc�73�J�O�zkI�w]��n�N~�V`i��N x���t��<}(�L���(��2(�dl�˗��$�ь����Q���p0�
#�
�>!�$�`���J�� �F>#H�ʺ���uj/76��؄.T@b�f!`{�HEy@G�&>�7�F�%K��$�1�"$��#H�5Ff0��B$�Ђ`�J �0�g]"
��UY���z��1�f왰�bNf�rbH�@7�C1�@��,�f��t�x�^܈��c���b����&8ƑT�i�@��Y�&���1�1�$����5~�����`��I JC�"$�G�4�U������x����E�3�!�0	Y�$���O��G�'�qa��cH��"L H�a�@& 7�}n��Y����W���X� i���iq�`2��� � #��D|9�IL�lI�\b߮l�df�b��q��b*]VܑJ	�"�@2�D"0����Q�dl�X�Z���woe�4`|a$��`|�2 �DŘ��`�0$�#�4�J IE�	��C���@�1�&0��f%��0=�I�a�� �3���G��0�֝��3��~��U���ŝ04�cLV�`D"�L��$��1M�H��(�dI��Y���1f"�D	(�Y3>1� F���
<DQc�T1�%Dv�& $Y��Ӿ���z������S۪|  x��1j�����g��� ԉ�҈�4B��"	�A+�D�H�D��#�<@����ő9�q�D2!��&y@�\�}e�y9�_g���~Df���^ʐ?�����"( ����0������bL��B1֨�2p�`3�!� <�8d���1�ǯ&bȉhF�\p$�@q�����]}a�}B�w۞b<`Q>�7��0�Q��n�G�D #%�s<E�`g��2Y����$	 x� �#J��DI �?� Da��2��,�HD,����& �e\�u_�����;O4Mm��LW��Ϧ1�kdVU�y���k����4�O�C��x�&P�L���E�����r��]���c�?^�n��4�v�^�H9k2��V�"�\��s�[�����D��ދ�'a�?l)>�P���qA.�.�&w*���,�6����S�UWDIf1����p���0���!D�#�J���:`i�$�3��Q�	҆@���T���"� �08�hɋ#�!����� B�q��/�3���߷vgX�$@\�u!` "#H�0#Hcb"�O��P4�`3�r��#��"�X@��� 
ܧd`��.���K��Y�0�#�7��⅐4�DG�I�`Q�"@��	��فF���$
��F>"�9n8��D L'�ԇ�!��f>���B��#��������W�+Eiܭ��]�� o- Q���,�	�>��$q�V`q}�� #�5f�F�0,����@DQ�bLB!>1��d ��wדa:@�7)�1F> ie���`�N{�W�z��T�n��da��HDK� I@&��cH� %�Ę��D�1(�Z�}� I���C�4`De�GH�E0�E���ND`Ԉ�@�
�S�Y�qԽ���ݓ��0LG�Fܸ��Q��> ?`Q �`i�G��"LI ��	#�!G��@���#�E�4~�q@���<�"<B(�<p(�D�nO�]!J2E��J���)v�����O�p�@�F/D%���T��)�Ȏ(��#�fD|`I����I���0���Da��H����1񀍑ib(�� ��d�B��NMOsά>�|w��y��Ř �8E�:��1�Y3|�� NK� �1�%&H�!��k��I�����0�� �N��`a���G�"��R��ŝ��&S�A���w�gx��^J",�b<FH�,��H@Ӥ�<Ia�f�"�:�L|D#��3�	�/��wK#�@(�'Pf$Ɵ�`z�|-SB�0.���	�	��XBT�,�E��m�����7���#��"�Z�	4_!�8���E�G�( �-��!� @���"p� 4�0�����>">��FK��e����$�`=�g�q��괎�nkJ��6�n1��ș;4��Cj��q[��������nBx_~��S�Y5H�kU���� ��VN��s�[w�K2��'+W�}B�����dW��=pA�)�n�2�����DG�ʺaR�ޱ�M/v��	*��l�R�cN��]ά\@�0	�����؋08�!F�wT0	 �J	�8��P,��"`Q�3��DQ�����"�#�9�H� ��#�<@��SDG�ҁj<@f���Wz�d���q��7������8`C0b鈣$"�����cht�ϣ�n�"���!"�W���+�4���zVv�E�!me����"�{���:�or�Igzh�G�}�^]���+�P
I�w��N����$�q�#eՖ����Q�UXs��
��bm��]e�7dzq戯���MO�ʡf����"<�3��U�ν8����Uz��q�<#^�8TGP�S��'���*���� ��ƽ]Ũ�R+۬P�o��^3�_gs{j�P�psA�W�F,�$�W��֊�8�6}���N/����[����ָ��p����s8�Â"nQ,�[�h"hǦ�󯵰�>��ogYiqkF>��Cբ�	 9q��Чò̮���ᮜQo2Wkx�u��(\��|,7�J�gc��=���O 6]��މ��˪j�V�'En�4FT��i���<�������X���p+릢g������ϕ����bn|�8��Y��$ή���r��#�j���m��oD��K2]�ٻw%g�]��qY�������4_jӣ��K��@q�j��ʚ)��dy��Z�\{��*�]Y^<�������G3��ޞ����J�c,iw��/A��ǳ?N�R�̰�K���#�9��?+*W�-L`�3�ŒB����k~õ3�`Wg���/3M���-�0���}K�gMA��:�^������m��J�}��v�>���z��OiG�η9���N�I��M������N�?Dk]����Xf��I�s�W��߇����%�ܪ��U�����>�8�����WeV���ҟc8�,�8Hۅ/c�:�\*�V�ϭ]���b�o]��G���PIeu��.q�s/Dc���g����0�6Z�͔�v��lu�>Kٜ*Y��{O���1���y.��c�{�R�T����BA���ȐQ��C�o<���e����̰O�G�i�j��,)1��R�t�`{~��4��������"�v+�n&=������e2+��]+�������Z�A�o^��ː���X�2�����~��ĜԱ�7��3,{����>Y���#�&�^8�Z�J*7�Xv;��g׊s��sB^[�+�Lv��C���c��������z��w!׾�J���Ps�A�w��_�&�����=vu��$m�Ԩ���2�JBP:�]�W^���mo��jrՔ�,F�!�,C���U���:9����L�u���c�&%:r�\'�SJ�d۝v_4w@�:��[�!��M���Ƽ����5u���
�k��b�����<���*,�
(��z�i7��lE�o ����2�
UD��L��Yz�IL��#u�
�x������qW��~��i�*!�<�hT&�t�Tr�so�+y_� ��>��^�c����$��o/� �����H�.yo�j:��
y\K�B�>Z�*{^zd>ë�� ������c�ّ���;{8�'Y��e)p�=�Ǖ�,{ƺ�<ď)2�#�J�S�k}�I�jN�åZ��ܽb��Yޜ�;Mga��K�[V���6�u�Z5�lӧ��C��Z���N��v
3ń��6m� -z�{pه?Qݘe�o��~n�o��m�E�"\�WC>B���'�Y�s�dg�x[�jw�&m��K4������ڝ���i�+��&�ì�I�����1"4�5�-㌦<�*Q��[ς��ga�����R캾#j��D�w�_����/��r"ײ:�Trw?#�z�t展�;3m��y�2i�m>oev�����p�
F�]̻y9�ă���blgp���#t���;B^��:H�[с��j����c�p�1�+QjεN�zԶ9DyM�N�S������!/�P�n���GѢn�
TWs瓪�v;?��E�oT�|�������P*�G��:xi#�04�mS�99�
��{h���sᛷ�`^:G�{�8^����'ڟ���S&���:ɩ�e�i�=D9^�)�{֪z��=k�P��A/l��vr�ë�]f;[̏S��w��׉��t_q��>���IE$�:�k�rb��bB1��ƥ"��٘(y;��X��򮞯X�k��re�%��t�f�U��h�nl�coZw(��SDy�R�}��ܵ�=}5@����N��RJ\gv��h�)�,xW���vI���	�CU)Ħt,'��p��20Xj��
����5�%-��\u74+]��F=�,_��&�<w�ޑx�ͯO��hh���o"�u���)n���j�@�H(�S{�,y��.f��a��Wj��t��מԲ�ְS�Rdv���z"���΁N����¸>��=�1׬F�M�r�\F_��qB'��X�uf���I,�qaZ/�HǸ���4�gS�=��\*�~��K��Y{1�xL��S���EL�O4�s��>#`���*��ж�]��s+(0t9Ӧ�[tG:tARө�qq�|d<4Qew�«�u	}�N���$؊�^����w�z�ŹZ��w]\2��9�s�t��#��]�����67:�Ĭ)˽��F��1��'e�2�6|'wC��J�H��zk�^�r�ٗB�`Մ�����9�������ߪ�g�O
�ZD��_��IR�RʛN-޺�=���u`W������R�vc\e�w�	����,:��n�1�	�*ί/Mk���Jt��js<%�]����=9Z���`�X�0���CQ X����;Х4�5�QyB}�*A�1vOzm�]7�7��]{
���R�^��������?8�&O���rʍf�K��c�8��r������t*�`맕�U����ޯg����iS&mZH��+ke*�0��ݎ�u���!�k��ϰh,83+KE�CŽ���3>��"�SV��҅w{߄A3X�5���U�
L�K��'͌�8�A�]ީ<ԃ��>껧~��7o���SJ]�!d���ٍa��� ����/*���^]�`ץb�~��Z�Hr���4�FoMi�����X����w\9+�L~���7�nNq)���[��A�og�4��r�����K(i��X��N�>�r�N�ٚ���q٘4.�4ee�S�W�a8kC��TY�7h<Γ��S����
V���=�%r��ːm	���k���B} ����;�v��AjPH�����թݫ:��� �Q��@A�d��Ǝn�{�o�V��-�K�-�;/|;��/�XC�f<�3����<�_N�[Oɽ�q�������;�����ew�ӥ��'	��%{��!�n1�fr�|�V+/)��|�V�n��u�1k� �jhg������I~���L��&����{�}���~2l����VC�-mwH����ǻ^�l�k�k�����ͿZ)Vn��Y�dupU�S��꣋��lu��fo](ěs��Ǉ���*���5h䯧����}JE�P���ߐεW+��*����^(�4{9�><�L�i{9�w��b��j��HeܹȔ¶j�ք�(����?,/˽��:R���Vq)�AB^kg�Q����@S�9��_�~m��n�C�z���E�*oY|6'h9��v�<r]n@����eN$#@��d:�-�YͭL����U����\:bI����љ�2�f�̀0 [N���z����̋��+�kg�gC�7Ecvy9Fz�2�qiZĔB^kQ��K�)���ҥ�3
�J<�R��r�[��Xq�V��z�(jc�c��UC{v��1�Ru,�w�[�����T:mi�*�r9��#	�2r�u}�����[0�����.)J-z;@��yBhg�+ܧ�ٝ� �{؇L7EbuϧS��Z�r�X�7t�W���rؗb"_-�?9|�TsY��@�ߛW�%kY�k�Z�&�߂^T�(��13�稪���ܶ�un�S=^���ހ��s�-�Nڃɻ��iK�l�O.�ZR~|�_�q�E��}CA��t0r�@M�5�j��+��u~ٛg�L��3����- �.g&�bʈVO�F\�S���k� ]�܉���Vw��?Xǻ?L�s�#"ځ�n��:2ޫMߝ�q����[�kvM�:Ғ��E�-��zա�O�TPI���MH�s�|,slV�EܰV�o
�7��c+���~Emz��FX5
jɶ�wU ������l�+�#�te�G�����WG�+ix�z�C��DN���B�ѳ�,ҝ��
����i<��P)�P�8�}i����kx�;���<MzҶ-J�ƛ`v0جk���g��Oz�����s5;odgx
��>"����:zw�S�!�ْ+pvm�"������ҡ����8=9��͐�Y� ������Vc�n���	�w�He�i�f/	�RSc�Q|F��;KѠV�7V|�{��8���}��:ѕ�c�g6R�ٔ��6�$�[����*�=ٝg�G�*��|+�Xr|����=E%�ɻ����\,vowuA�M���EH�t�F�q�Φ�qԴ�ET]�e��}�`d]�ߑ�k�l:pV�����GZ��tG�Y����&v�=r�]O�F�^��B�ٛWWƂ��~�^]�=�z�Zy�����]�RH^4���'l�߯��"\G��1=�=���6t��b�XU�s�}1Vz��E����i!�l�����_/M$�G�N���_�2]��a��>E���#{~���,^%�����k�mԿgD+�9�h��o��˽��R�y����S�U��W���o��Ѻ�%�Һ^�E��������8�TEb�J�	݋U��,���~]:w{��>�M]_x.��^ތ�Z�z6�������D<od+}4�t4���| �z�����͙�f��1`���E���D��x�ˋG����W�|q�'�)�y̓�����~{k'��<�scSI�h��E�vM[ݜ.2<s�^_��;��񠷵
��F2�F�
f;������|�&���f�vC���\x���{Sʝ��kx_v��=;�'� x�-N:�;�噳�֚C��O�]�y���1$7�]]gtO̘���ߨ
�MNy�{yݸ)�F ��eJ�U���Yo����^p�.�*�70b��;c��XS��GQN��e��ȫN�q,y��Vnt9wl�6���Ӂ2����Q �bV�R��D'8�BΊ(��t��t�n�A�!��cuʸ�� ��4^Aֻt���<rq#���!t2�Jw�u8��!��ú����Д����Xq\"�x%[Q85
�F�wp��}�8�@�Q�\�?*�u�{� �)1m*��r��p�'7�sf�6��S�d�{v�ʋ{�J���S��N�leM�a<�"��ɕ}W��F���h��W��W!+9_
G��7?�2�T�Ԯt
���l�c�8F�����Y�ˣ�9iE�n�a�6F!�����,��ں� ��\�9�i%h=X�cf���R���w�Y�'�*�m��r������\�"9��a����ʷ�X=ܨ�ޠ��Y��+d��ю�b����Y�K��&.�JoMb�X�;f��y3�a&0=��[A]*ݓ����zoA��\�e��!�6潵B۫G���4&��1MK��	.l7�V��Zi��5�4�t�i�R���Y�h�Tn�.\���p�T�v�?m�͝6����@؀4G��FV#�7�W+��.�R�:hR`I�pA��iol��{|H�q�jgz��ph�z�N�Zđ&¬3��k���v��	�Z�����b�v��1��9��5(i�� ���;��l�����"��-w��Jĭ|_u�|؇�=�����3o7'W.C��bm	�8���
�wS������p��+]�3D[�R�^t��,��[��B�_]���Te!�y~<"zw[Ң��~5���,�ٕ�P&�B2�̠x3�f��nR0��Q��vI`�umP�ڻ��I�XH��OM]j����{�G�6���w�����Fhu�'.a	��a�M����[qU�K����v�hU����x�ʎ>�y���lh �3�2a,`J�|ԏ��_n$.���ڳ�G�����5�[u��i�j}J�pub�U�ι���ͭEբ��o:�Lu���Jr�����V����Ř����=0i�p�c���&�w�y�ub�sy�~��.X��c���0�bOZ�Y5֎�` r�<�����*^�S�2jV��]��l�͐Ω���R�����<f��4��u�L���]��e2���ʍ,#f�$�����t��3�?���Չw���TRh��Z�աj��gV���ֹn��8��{�\��<���c��~��n�32ó�������{�(
�2Niժ�Wg�ֿ`���l�&���N6撚ζ�#t�Ъc�;l�(uV� !��gnEW���iv�F�V��w�]�]in�iy�k.�C�Ʊ����ɗz�M\�[-Elqk4[�;���$%�d@ξ��_;[�X��F��5�~z�'>���X����Oqp�Ҕ7;9��8ք��*K�u����jov[�w:�МuϚ���qu�����Jj&�B��6nV���[Y��b���w-��Xb����z%Y�Ǳ�~㷖��@��#VD{B���i�ݿMt�5~�]��kr�n&��YO���k�j�
c��i&�	�������ΦȬ]����w�Ygg$^`����S9IK0L�e<�{^3�<ݙ�Z�<�f�o�u���� ,�bz$�,U;>>[�)k�&vf��<��yY� Qa�/<�.�����^��9�fS�A��-_�H��}��֫m��U�-��{��r^��|.R
x*�Q�[�[������k�����s�����>�:j�/k�,� )�"�.�ߩ�|Nr���j�yZ�J��/N;�r�L��w=~Ԣ�R?G9a�7���@mZ��Lk5f�c"�����i���]��ҭ�a�o����5^�#���+�7��Q�a��q�<�h�u6B"�6x�tJ'g�Q.z>������W�=��9�mi���ΐ�k0�����<�h�0�͡��'<��ҝ䞺F��Z&�#~���sF%Ľ����-�Adp�f\{���Uҗ���/�y���p��������W=z��N�`�Ƃ�t�cCVk��Е`P�=BdT�։�QRiodN�tZ��O�s�г�չɼ5\9��Y ��,��3&t�GA���M�ΆX�W9���Lu��Ys��Nގ�����Q:U#3��ѷB��T8�/{��*��^kBv�r����`l�>�H,;���L~��n���z=\^�Ӯx��@�7�����\���RS����C��ӝV����C.���CJ��`�~=��a��$�R�4&���g7�S��4�D�d�G^�;:���'��(O':���{Ba�櫡����h���w�����ܜ&������Ŵ��u^�|��髣���w�؝4W?G�������^Y�IN��~r��j��5�k�>f=�__�W���݂������S]��H{k1$�d@�iM�n����Nm�X�-E_�ҥ�W��A��4D�^{�Ӂ����;Si��u^"����׻�-w��D��(�x�������OB����z���~�+�Ŗ罁��mL�ЩSy�o��md�ۍy<+`�3o>��n��B��<��o��]�|!�.�\ˣ�׷)�������M�2 �tͻ(ue������q�N�э"swkN��=���s� ��ُ��L��7	/��X<�ɋ�����:�9^�.Ԭ���\]�Ǆ��<��^;�z�<l�}-]�\�W8Ηg�c;g��S_U�T������!�k{Z]6��q���Q�B��n��ֶ)�䫱�e&;0f�s���uޫ���{d܊��5 �⥗�[j$.�ڎ���tMgK�%k�E֯�S0��qɷ�����|���
7��R;P6G>0w�xV�:;�^�E՝!�ߵ��njq�2�`V�X�cqҪq��a��Y���^[hg�=�s|T� �	oB�
��+�I<)gN�U��t�C��(��l��q��|{^-�á�]��Kr�׈�i�<�}H���zVE��nǠ�܇t�:2���L�w�Å��c����E��/v��W�cכ����4�k<$d�7��P�~��
Npv����[V5�ܺ��+c�[�l?-��0|��1��N�A�j� �ϥ�{$�q����n|Ǥn=��hO���dtru?r��e>䤞9S�g?/m^���%l���q�X��K�ko�ɓV�h6��jv�����kU	�3���Y���X�'�E���>���I�n�[0�EKj��%�uez��;�:��ro�%�c��{M�&��3S�7`U�ِ��x���������o�FWM���P��S��Op��8�b�tDHmfbp�=�{C�=;:[�l {N���F���I������?��C##���;SO=��]����-n��ü���YK�7b�;M��Ӵ8�f���E�s��4ص%1U�@���1��yEzC����]u�ˍه�I�X��ݑ0�
��)�Ԛ������/1�^`�g"�������+1��V�+r#+~N�CgwH܉x��/*�y�ت�U�h�B����^`�T�i������ G��]�uhk�4��Pk�G*���k����d�S�-��\�ܻ������.�VC�^E�����N���O��~�c���yZ��K����Q�ѷ�.�P�f{�QA�1��C�<F��o�r��W���w~��nU�YW��ܑ���x��]���l����6'{<s˯^Ux� W�*�[0�����^�!'lzf���C�[��ԡx;�V��3_U.�H��>����s1��	��:�?�J2�s��y^��m�g�}k�S9gvWl��۞w�B�{T6�M׍�3���^K?@:a�m��{(e�=Q�����;��?�/ˈ{S^���6��n4����Η��$Vo�k�C��b�~	@��̓kZW������{�E�Oj�sn(!�7I�=OY��l��Hv �*��xϳ7��lNVֲ����ӂ'% 撇o3J�O�u|��Vd��Rp���X�ͺQ��H%�ͱt*�L��L`���Bu���߆*U�ޤ3�}*��Νϲ.�L�ƫ�9lT���}�ݮ���k.�W*�f���vuܛ��N�(c3;x78���kU�@��l�cPc[��H���{�YH&O���:e�ц���8��������i�X�ƏX�ɘ�9o�2%ۮ��NWO{0s�o=���k
�;I�m�=�6��.v%J�W��_�.g�o9C�g��۲�4k��+Y�x9�&��X��w|�TV��j̷�_0X�Խ3��U��I�_����Kv���I�V�蹀�.�ֱ>�X�F�g.{S��^i�_#'�g��
/V�w���*^7xJl��$}��w'ʼ����T�����*nT��l���2Beܬ�重[4�je�7�NE��"�O,�5���9��}S5��ǜ9[��/FJ@{^�QP�<��m�w6e�W��Ǐ����[5)^���l�b��!^V3C}�(Ǐ_9;�a{ϗ�7�,�m3b`n�YrК�f����t�0{�a�(y=��3��M��{��#�+�{c
���c^��i��3�G��
W�I��Ե��|�o_
[�3'l!`cG���l�6w�T�LU}�=��y6��j���Eދx���ײ͉)��ǅ�kF����DBĲm\p�Z1L�N��8;2�4���ڬ�7e>h��v�ޣO��/;� gGл��#J,�ʟ�P������.�;��b���6�&��w_���v�d�Y�Ǜ�VfҾ�>N�4(�[�4�fR�1�.��wO+�Uq���{������
��[�ֺN%�gc����\X�/o{)?ڶT����Z^U�L�@-y��5�!�z��S�׎��eb�Y�N�^��&�
��{��Z*	+��]{��vdZx�}�(��/ȧ��jx��]4m��=��u�\��M�.D�Hu��t�j-"F�L�K�~~�rð7�I�U����6Lno�=��G�������TڄIZ�z�7e�O�F�h�+�z%Uפ�]2뀮Ƿ�S���]C���)����z�"�� =�j���=I=�1��ѥ��!�Mz�_�FF��ќ�#s{��23@�,_d��v��� �K�ҲO'�]:TX뫕�0��:�k�o��cYٸ��~� $3��@ܻ��>�b��<�������"]�����=���`�x��Y<j���.^�Q���u���[UEM�˻��xv��38�/j_U�x]e�x��ǦZ�T��E�Wu3Y�eA�n���;۳ͥ�)Jp6(�CF�B��`ڽ�Y,)HLX4\�uʗ��pP=*��v�%yf�ZS9�u˫b�a«��;��3/ٮ+��˔ԙ��xN��kZ�9m���%��cc���;A���4�o�#�aOL��k�쫪�:�F�j/*Ů�p����+�.��/wלj*@UEa�k�y�q�#��D�I�w�R��$�ն|�z���s�#��y]a�6e|�VR�P.~��j��YT��8�`��&�P��q����]G3�^ћ=�~8z��x�;����*�J��L����~'�OK��1O3�����Ӯgz���J9���#���;��ۚ�̍���6k�f�}���Vxx!��ߤ�ݿ?	�@�4��m�*����*{����Z�!<����g)�c��G]�J�z
���X�)�@nx.��zϩ��ϩӟX�i׀��0�~q���ܵ^�S��D��{��hR;��N�݇j�/ujUF�f�����N�X��x_���dT��7u{����*Γk?~�P����7�h�营�a�|�ێZ}�g�'��O�/nb��Dj�z^���H���ɋ�������H �{��+o��R�|���^(�������D�~gF�*}�]@62�Jfp���{G%7��Z�8���V�n�⩃��4:���s{���i�Ô)�Nl�ed�'�f�Z#Y�ݪ����8�@�����pӥ��]�9�V��ئ���b�w*)]Ƅ�����[�cXM�(���J����	�)a�i�v��؅@uڡ]#��/�4���I��sO�[{	��JY1;`�D�s��k���̛#&_J9��0�~��մ���m/T�jo{2	�{�ܽ�t�[�	��gAi
"D���䥢Ƨkc�S�o��X����Pp�G�ۜ���u:=Bx�|)����݇�;���d�R��r�;GmK�o�7+*I��:�y:���])R�� =/��w6u��~�z��ļ�n���3�=�7���F��j�
�Š����4;�]ۑ��z}�[͜x`W`D1��N�6�"(L�X�~-Y��+e.��=�ɻ��]~�SW�q��g��*Ʉw7K�P	�v	sY{�j۬�c��b���f�NW�+�ǛĺO^��z�����r�H�ׂ#^B���+��=���r��0�ֽ��vp��l[g[fMl�LW �>o׼Q~ ��cڇ�yny�V�S||g�{1�b=�aH_�@@@���툦��7g�z�%G���]E�+}}^����V�p�v�~�/�T	��]zyS��]�"��R���H}�j��D:��u��Z�P]�C1u>���Wc��\�;�K���J�Q����
F�[�r�t���g�:��wx��R���7Op����;{9�e�ޮ��V-���w���Y�b�mM�TVY��l��e���^p,�Q�ʗ��2����R��6�ԷzŨX�u��? {���潓��2�����.rK�:=��5���K���.?�kµp\�r�x�ɑ�Ws������jK��k6a�&}�l]�d����F�|eV%��|�mO�3���h�]96|���`����U�=�.V���xEoF��-Xd11�^��=T�����������q3N��yLb�S����W5/�f�T��z6��ƌp������ u�;pǱ"��ɊFlE��	�R��<�����]aq'E��2�s��s���[8=l��>L���eæ��v�j��f�Z�/�r}P�Vj�w'|�s��#�}�Y����=�io�]�k��{ݙT�w��^��=q�T�o��uL���x�uw�̛�4el ��g���.Wj�J�nS��Y����8gm��ǽ�T�f���/���~iw
A���[��Iᷧ��45	ο����3o2-Z�Bj�jF��b��?��0���.W=;3����!���6e_!����1a]�P9j��Ȏ�+�ǝѕ�ԑ�V�	��!���b��]w�~�\����!5����r����Ӫc�%��й9+:����O:�w,"�:��mF�F闡j��"���]� �E���mowC}H1�{3yڧ.U��]9��U7X=�H`nrez׋�[6 z��3�q;-?9;OP�����k�]y��>��%{ �گ�ժ�'t��"dÜ���ά��]���<7�1,L���z�|���*�31�ȶ�«�T��ov�˗5�����L/C��6~Gr��MKN�"<n������ҷ��ǿu��˪����m��>1�J�=H&���x��.$i^��w���ˍ-e'���޾^�MM����ڝ�8�
�2��m^����6J�>�<����P���KQ��7o�V͗^xh��{�c���Q+޾^l��ܤ0r����3����ߟ�fMו��`�Ք� �U��v��֯>�k�{n����*�+}+ŧ�$=^�.��ۜ�bwa���W�Y��Z�g��̟-{I΋�+'��y/jZ��K���(йb&p�ַ�B��F�-�;^r��n0�ȿo��ORG4>�Rf��#�x�VA�G��I���e"�:�$��a��[�r�!M���Ő~55��/8���[�F�^jg�yu�]K���!K0Wgc�8D���]�[�������L���f�XF`H;Z5
����
�fouc�q�r��P��
�QT�?�	#'�&t�}Ńsoh�T9��B��椩�2��WU�Ɲ����� ��O ��=@_;�iʼ��bv�{�r����0�����qD	�d��O�%�X�Up���|uF:w�iۛS�Z�N���u+�ŗ�j�Y�Xv^��p����&hqF���������42c�_[r+���*v�%�{���VT����S1��pC_=�qīmu�"Gke��F��;\�:�>ֺ��6�E�i�׫�ے��Ѵ�m���vr׷B�v*Y�ɷV�8�p��u����'좶7K�4�v�9n��ҕ�L���4�,�����/�㳝�j0]5@�3D��j���923V��R���wa�hV�e�;fa�]�#լ7��&���e��'�5�����͗ZL�2��e���P�hy�깎�W�Dte���fK�x�4��n��YѤL���=zuЗP��W"�����+m����%~U�+j@z^~���.y�b4���9i��F_6if,���c�s���U�_[0SHX���.s�_0o/WZ#kzt�g�]�>�]k���{ݾw���݀���A�6,��4�ܱJ��/qs�G)�fʵb���+sz��%�kl�d5���/j%���Uހ�pېAm�{���٠7�c�\j+Y�fB��b9ô�)��p�l!�³dʕo�����Ӳ0�4L���%d��YC��e<�ԛx�gU���J�4\{+R� ��m; �b�^�M�����Wdĕӱ2�F���Q{v�]G�#uxj.T&�T�muel��o�N�u��o5x��<S��S�յ���N��d`�!�ps�%ee��v7��D��p�̝֭�����scx(�rѩ�}k�˽���r�q0(��B��ge_0s:��ӽ����]v�����0�-�Xs��`7���|��ݔ_���R���72��r�:���Em��Iu�5��4t:�g�-mJ3�r�]h(j��;���C��{#T[ǌsx���Tn���,]���\�Y��r�h���b*�V�Gt�K�_#�{V���aC��9� ��:��<0;�d��Z�I:�hk����fN��tO����f/IJ�~�V�M�{7���!C%s��3�ȁ�d47��;L�h��Ԥ;/�;�*���,T�=�-} !Xg_����M=(���L����e0��:�)���WvN��{_F�Y�1u�LY���[a�Ai�:=qsS��<}��ː8q�.�i`��%�C��<����h����U�+����q��d��Vq�Ҙ���Do��V�]�\hC��b��<��V��Ұ��N�*l���pa�m�H;�����t�^����b�Bh���%FSr���v���gk|��op%1l�ͳ�u[�����s��d��W��7\�f[|��/]h�_3��7�?{|E�n�g�a^E$�gud8tv��vb)+���+o0��`�?�Acɇi���G]�<�O�E3`)�]b/ӻ��6�k>,]V��?xB��P�e,͊P5"�^�Id��<�ۤ���o ��8��U^�ʂly��hc�#@��Ϗ���Uȷj�}ý�0NYY��x>�ﳹX�TG��ПQ��C��R;w��Ibp*�1�FN�5�K�=���u[���*7�s�m�hN ����� c����<���~Q��9X��Y�3>�4jT��9˘���ڿ�Q�pY�L�**����a��y��M����ϫ��mC��kٳ�(#��eb�R�)d{��� �y�m�z��n��\��i�tR�Z��gES8膣�=��W�����#��mΉ����EꋢE9�|�Y�Wn��UҦ��#^E�hrw[��z�h���ؚ�D�7���q�)�<{٨y�W0P��;��^}����7�ڜ���v�F������ߥڇIf���c�zˁ
��T�M�ʨ���U���kW�����\$�<��ջ���R���-15��1������@�^�8]j���%X�[Z�Q�K���N�S�\�6�p��a�^�CNKk��r�W7]ML�i����䤻[z)b��1cE��ebwi�مn�T.j�;f�C�iu%�8G8�#pl���N�ۭ_^�~�^s�A ��3���	�-��*�>Cβ�ޓ�?
f,��=��-��Gܡ�����ͺ���vVz���~�@�\�2h>�Cn.���5��oH�{V�珥�����ٮ:���?t��~e1�B�{NU���P��ZH�R`R��s�oܽF.�hu�jz����zt��}�pk��zr�s$vh�P����Z�>��}�CV�3H&��!N��u�48�r�?F����S	���&H	���爫����}0A4qH�~��'F{�q��͞C��_z�����}�9�-�Q��j����0ׯ�X�?��/��r�Fw
z�5~��������VI[��m��-�T�<Ų���=��r�X�V��;ی�����
���x�c��j����U���'�!>�h�ȉ��zϬ7���L9�z��}�*_{�P��e廑
��T|�n�SטV,�Ȫnלޫ�M\=�Z~�ӽ>:�~�6�X*M�l]y��������4D:������KC�!�Y-��X*����]YǷ�\��b�\OB����)̠����;�T�lu�Ѕlƾ2�{�4�;���tȷB��r�`n�0`�=Ym�f��HN�:f�,uq�.H��D����,�&b���Y7+�mҙԑ���9�e��=@�/��^qY5�(��nJ���W��=~{ӽ .(�T`)�m���K̯Μ�_���=����7+�.���k�
�=XJp�$ѯC��3�t����J�s^/��BǙ)qV���R��!�xn�
����m�lUP0P�� �TN�O���y��E�_�ͤ5ԡR��J���pmw~龭S-�o�,U�C���DI��������<+s�z�A��*Q<�j��:z(�������	�1�Hϐ�\��C���A��ęM�|8��#8�g��z���.��\��zke;�u�г�f�ى�j�t<j�i��=�U�}�I�̷?��]�~�2py�y.y�]:���5/n��e��=~��fP��r�
�D`��t,A��۽�9^���zM3�-��������e�cه͹2�M�͆ Jw~�+|�V���:����Q%�Cۣ�=����sz�Ym��y�������[NJ����$�QX�]�ڢ�P��վsK�^P����)�H6A^���`:ʾ�M����}z<&��Xx����^�9����qyt���bQ�ܶl&Zf�cJ��T�2�Cu��u\j��wY����F��`�$�ۚĒ��Ϋ��NI�p,�y�{&�/�nJ}��u����7����׌����iPuf��:��@��
g�_Up0-�Vc��A;����o��h����fnֆ#�IB��"�p��R�b��!�)W}���#��A'yr�K��w�m\�p>�<ן���HV��'$������k1�N��<���y��-J{���+������i$mj1q)�w�R墆��㌊ld��tO��	�]+N�1d3bO�ȟ@���%��w^�&�u�1����R������zsWY��t5��;.��V�~��5��)�RG�&����=^&�����化��p�A]Q��׈5)��ϧ}�G�a7�;9�I��p��E(X�^����@Д��Aߴi��+5;ԁ��
p���rV�ټrn�RQ�ϓ8��9��a�� В��e�G�3]��8l���v�=���V��Y��~���y���y�+�#�= ���{�ZC��.��J�k&,>�x�����fq���רb�54&�~�uqc�Ȉ���\�_��k��w&�v��9��� ��j]|+�,x֪V��ŧA�n��;4a� ��^3�,����!���bWE�V��"e�lhْ����O"�eٙ ,��><�b锱+\=\��w���\��ޥV^L���N��m#!Rm&�gϔͼ�>�wj��	�G[A>���*���;!�ⵯ����4��+ǭ�Q����oc���^�� fWM�Q�V�]�����.��S���Q^�X9�֠�b��ֽ�������/P 8=�hk�?Mڽ5�ɊJ|]SM�E��p�)wg���FE���if�	ޔm�?\��g�K+r�.xxEo:W�;Ր�)���@�����)N��bXV��q+"�6�;��G����n|�.'�:����j(=�;{s���"�7�x$�����8޹s�����ue%Ի���<*|�#]Ʋ��y��s3V��}q���y����/�0�~�t_�f�W^�>��c��,^P
����+����~�/G�:¬w��D����osE�[�H{ز� �׭�3�~�黹���<��A�y���/2�P��F:��}�P���"�x`�4|/#[�PܘZš�Z֡��k�X��i�l���fM}S�.di�0���h�V�EY��Oi�i��ETɻ�s��`˓7԰����ER�UːT|A�F��bˬ<���������Z0c�<hU�g���<;�,�֥�f��NU�
�6(_SV��s�(K݄�-�݃ns�GyR�C���!����h45��9[�-��UW�/GX�+:�
}ϨlBIN�*�n��k�U�V���"d����[�-^�8X����u�j������s�k�Ԭq��T
�#��G��o�K��Լ�{K�9�I�kU�%M���R6��p:����� ^UQ��ǚ�������;���ӽ��YU���e����\3jy߰xD��ۺ<��a�)�S��r����޶�hn�G���+���QLB{��m�?'�	{!��_5԰�K׹���j��������ْ��]�Gh��n�Z㽜�Uϋ��#	k�]��/�}���[+��9��N�ٟ�_i����`%oLǈ~���=��{��%Ѯ#�����¹y����ּ0�cpuDzr|���~gu���G6�F=��'SS6*W�uvCF�U~�g�{����4�m��i��<'��ۈ'fh�)��)X������P��7B}^�Ɲ�����G�q�u���n�x'|k�����Ŗ*���{�L�8= c��)+Ľ��D�Q먦ۡv�1:����1��5:�8�T�p��b����3ό�
��h���ӺST�r�/ی ��}�(F�\����h�����]-r1�oAp���^��K�wed��X�6�|����z(���ݱ�Y��4�N�o&�݋�fkS��"U��x��jf�s��{�*j]B�Աq�	�О�B*������ʔ��gئg�4R�q�ۍd�w}Z�M������E)x��+t.#7���*�S�|�V�[���^���0;�OfC%��\����^<U���w��;�p�M��b�`��_��4Nn�t�i�I�ӌ@��b� ��Ҁ4����m`ʾJćӢU ~��8��I{r�m�쭍�tlKn]�t}���5�%���5)(������x�j8��<���\�7N��D����*"=��~�:�qܴ��u�6U�[��'֭YX�g�7����P�V� �t&e/r����]n���^�vx�j���C�p�g�+�Z!�B�^�Ւb�ӹ�*�p=�Q�~�/!/UW�Z�=�����U�[��,��r�ޞ���1�2D<��h��b��5�1ݯ+�>��lk�S.We&�g�sށ�������:�'~�55�I��=N(�x�}�qxH��(�E�9.Se�R�Mn�\�O��۷�
�y��i�P	�
ڻ��:8�H���o^�ܜIz9�g��nV9ݒ�2V� ���B���_SlZǵ?Kh�v�vugN-�Z8-����cGYz͖x13J�0R��d=�,��j� 9�ݓ���Ց]x�ʥ�;��V��/�-�n�ftz����p�`�N��=yN�{��\�o_���G�s�h�R�M}���i�b��b��lf\�3��]�K�Y�t��U�n+ 5ca���r[���]z�>�@g?^�˺��!��|�w��1E�|�Vz�Ć#\]�.����=9q����v��~ĦI+D���]�L��l_U\����1p3#������ܡ{�����/�U���Mh�ٵ3�o) f�{S��y;���Fǽ�r(���84b��ub
x`%�ᒅ����Ӷwgr��x�9���ڽA���J�:ίcq��
�7���`��7�&<�G�re�4���_��l��;�*�=N0.�7��ˤ �k[���ꕛ�3GO�n�T�^��������%H�;��0Ϟ�w^�L b�w\�£�fݯ-0��'��œ�w���j���vs�ri��;���K�M�,�6&����$��4�BE칝Aᕂa~3c�<��:Ւ���<�h�#����xac0~��^@#����ڍ^g;�u4�T�c+,eõ���&��oI�I�*!�J�6D�Zu���X9)�K��tN�^wT��KFò^5R�_#�logt޽UfS�T:��qJ�W\{z͸��fm����knܒ+-�xW�Y�^�4�=1#H�[��B��5�eN�jY��~��OK8��mK{�Lf�@�7�G76א�ڀ���՜�I�vr9ᴳ5�I�of�ŏR���,��zG��{{��i�%da�^Z�kd+���e��1*P�pX���s�ӕ���ƪv�s�R��y��ǵ�hc�����&n�YS6�\��iV��@Z���������J�L���ƞ��T�z���t�Ų�Q�~�C��j��w����v�*�v��u-m�USR~g7͹ ������w���"����=(�o��c���m]ǒ��,��hu�Ky��cj-�sS��v��m�~�7���z�6�uOU� c�+�s$�wqo�H8����N�p��^ܭq�zc�<�d7M��6������Z�П=��둂��y���Y���ˇN0c�Z��/�&d�+�}�F�T:�od�Yzq!�1�MV���;'٨7�\���̾�Tcӭ_+4oo*bx��(e�K����|���3��<Y��mu\�K�N!��%BZE�msv{�%t�fݦ.
�N�X����-�Sz�]��w��,n��G)�"ɽ8.�%mfe��]P?�Q��K���#v
5���g㹵<O�&(W�%���x��YN�����R�R���voٝ�~9P�2��+(��@�Y��G��bsn�[�saV��:+7q�h#�H���S���6�lf5ܻ��7C�V�	���'�����3:D�re׺7���0fq��Ä�055�3oz���b��sƜC�sUCʣ�23�3e��e��o�g9� $�;���oD����s��_mi�}��0g�b: '���j��Tո�ȼ=�X�W|YD��b�&}���h�J��n�x����(HP}u�C�):���Ǯ{s�u�ss��/�7;�W �21W��霾��X��Y�;37�3�?c=�s�. ��U>�:�=W�o��8>�o�-޽���Ϯ���.n�csE��Oy��н$�bz�B�iwLY#1�]�g���h���z�,�O���6��m_�d��=P!��G�N���뗂�s�׀b�z%�E?�����/z��t7�_u��t�Z���՚�Gw���3lFw�(��w� ��d���JȾ�����:^��~�2pQ�$�ª��-u��.�97��k��'�Ǵ掭ZiI��\���V	OVR޸%.ȰA�%�q;-�o4�4S�FWl��F:���=g�Y�WV-Z��8��v@��C7�jI�S�L��s�Ve����G��y���9��>��<�,���ՏΓ|�lT���Jǁќ��..`�κ���ݖRwy���:n��u�g4���3,��4�	�c��e�L)��Zڵۅ�T(����ԣ���d�RE�V����+��l�]^��m��&��k���M?��#�%�^��teM�3�l��Y�ei7i��5f����ܵ��:ʕ�pw��n�A�\���1c��Ƃ!��Os9Ι�>n��/G�t0@��Ǜ�{VvT(�Ò.R�*:��M�_<�YN�P��v�CD��6�u�|�����mQ�W{R�y�vt4��x-�Eme꠲-U�����t4s�O�ؚ��c.gB��֒�WJ����="���QP�� �	n��l�F�
�,�L�X+k�{RN��=#{m
�v��H�{�+v1Q�J�%��:�=���Pe�r�'"��(f�Gs6ޖ�Q=u��b�Q�V䕇.�_86��k4I��1|�=�*&�b ��-�uYĭ^T�x��}a;���5B�-|.���i!o4m=��v���{&��r��{W�|���m\���rV[�{[rpKv�r�׋��X�.Uʥ<8���W��-���V�wj�<n�^�ч
"0tsک'q�y�'� ݽ$��d�['7z�/�����uҎ��%�I�H�=[���	3N��;�]C��+9#4	��Y-�姅֝�|�r귗:PYS�@��宫̔�1wJ�uh���/.m�lХ�q[�I*�K"�Ev���t���d���$��*T(s��܂����xN�=�-BV�]np0�˝��u�c��B��Uv��Sx�tYZ�5�K�if��h�3��v;F!6md�']#Ǜ�sc9P���~U���6�_Vu�\9�V���[	첚t��l��1����4�:��kh��ʺ����
�ܠ�@r��d��n����Nw0�����^���S�u�z��#zo9��r���XBX3Z�j�bL��Q�&�Pq�
yoڼ�tLP���'kmva�����rgY��8
NۼQ؟�$�{RȔ�]�7C8�w���s�>M���es�W�o�l�	N�gc�s�jG��]�~��Q�0su¶�3ө^Y�gZK@��
�	Y���w71m��~\_	f��b�n�e��II�
�_M�:�cEe!��ܓ�.�9����~Q9Ν@���u��.�&¹�����zv�VЫ
�݈�X��[���_ t�6s���Й�Nf�U�i�}͚zM#���1��8N�"���<���֦t��	�rk�yt��T�;}�lP�گ
��a���!��c�gc�hmv��;E~Y��z8V���Ǝ-꣮��R�KX+:ن�u�A8��:�3�Z;3p�qu��mɢ��j�PK]\��Z� �̆�TJ�v&o\f�����5����t��N�`��f�G�8��o'V��.��D�9�B5R"F��K��ܻ�fj�T�%�0v��!�z{���o�������=� m�~��Ik�r�!��혲B��Ew"��/�>[�g�я�����E��������s�ꨘ��\���:�>�n;�Y�%ƭ����'���A���&�#���洵]����W*��7�9��Ɵ[ˑ�K��pׇ���f�K�q�O<	��V&�s7b�s�0��f5:�/��F�.Dg��=݂ku߹N��=����?$���L8���>]�����8ݣ�Y7�9b#���>W�բf���i�Z�M�N�����ϊ��L�>�.'�F�;6�L{d��uN�x"p�`��^�u��j�l˻4V��3���k:rju%��O̳&�_0"�'W��}��J��o��v��0�+$�u=&�j��<.�z�uE`3n��{�>�� �1{�O� �/��O²*�����_�vdӻ�wg�S+<�9c�'��;�x����f�lfϵ迾�a�m����%�7�]o�~�=1t"<��@�G<���]]Ls':�b�H�^V�M֕{���l�c��D��ȅ9L��� ��Y��mM� +���EŇ�ء��J�p��ݝ���]ur�E�`ryh4{xb5��9o��Grj;h+w}88���z]ۮ��NTYlp�92�H:βt�1]&v�^���ds�L6$�)l�55��d����͡���!}x�~�js�:���	���J��=Id�{�͟UZ<2O�^އ�1x�,��ւ��#S��T;����#KxB<K쩃���4�T<f@+���ɵ���>���vyו͡��b�(Ϡ�c~�u���ƊG��d!����.�c�˫�	�6@->>c�I�w�w���\Z��A5Ϊ=4t��{��
���XM1��㒜�vK��}Z73�Y����{�=�u��7�Sb��3:���@0:�� Ùk�K�3ȹ�3���u��T$z��xo(�7�I1���ګ~�W�؝��^��L�x�����=�d�G���|i��ǆ-�j]rgt�s3��5o@�kj"o�*wyj����`�*�`V��J'���}����>dW�et����렧7�{��F��i+a9�e��i߆u>wȎ��/�Dɟ+�8|l����X�T�(��3�R��=�tLzɾ�����(z�2Du���.s#6/�(!�]�f�z��>���5C�+ʹ� �-���R�3���z��ҽU��B�{��{��R��%<���1?�6�+ʗ+W��晟'>�5���p�D7���I�ҭ���F4��D1c�M�e�%u!+iv��Q^�v����f~�e�\'i�Q� �r{7�q�����Ji�
�:�&�����3�t����R��&��o5]�����)��v����:������}%(�2��d߶gՐ�<J54��31��{=�Sr��f�^��3G}��W6�>N��>��ЌO PC�����խ��^GJ�NNR��
�҄��j�"І�4�+�!�9O�Qo;TO� {��n�����P��C�ߺ����u{�론�u�e �'j���/�펊�7�5�s'u�#����w=�b7�J�j蝎�����z�o2hu�������%/<��ϯ����T�֌g�'���Y8�m��7/DO�y��ю�캮�ѳU~�T֍ׂmf��\�0���v�v|㫧��F}i��5�7=|7T����T���hw8�(ׯ��tm��'�WE�~7��wdD3�Rf얻*%GZ��EQ��Ԩ�.���t��e���������Sh����Uc��x���M���n����U	�/��_�G�?D���%����!��ע��f�
������+,��7��_�V�^��'ea6:;��_�p���J݊�Kv�P��T"�u������������m�[�־���9T����{��~���*2$Wb��)�до��=�r���g;�%�v��ѝj�Δ�&���Qʚ%�E��^1�v����T�<�Vh<Z���f�O p|;�a�M��lZ�u�yN�U 7V�r6"q^k�W[�����$��(]i��vm,7\:���].wW�(b+�)E�\���v��ޣ���zSCNv�A	�6R����{%���[������:sv;�;+xYņc�'R;D\��1����ma^�P�*e�O��v��C�yVJAa�1O>�ۇl��qӓ�C0lf��+2+��{�浓�}�{�g	�
���� ��F����r خ��3�n�}����/�L8�����R�����]��M*u}=��7��r7s[�˫�4싛�W�����6{:G��nq��1��oyF��������P*S��^����
��wv:�Ϣ���0����o=�1�,\td�ʪ;9�/�#�ug�����"rx��r�B�w���p�h9C�׶��{�к�>�~u�LK���ު���j��Z�ze�I��'���o��{�ѿ>�'��*#c��L��Q�HqS?�L��~��,{�~~���?��3�V��#�~���{�~�%}�� '0{"%Kʾ%-���g�ҕM\VN��"};�>!b��:������b�c� ڍ���߮�|wbxaɴp��v� $Gzu+Kwo�b�.�#��*GJ>6�����a��Og�z JF�������R;W��{���h��vh�2��<��ĥ�P���l�>�t+G���G�L.��UW���m�1z��T��'C�O��¢4�t���7�J��C����$j�M�ɅB�6F����܀�^��N��{8��199��c󌋘�y��BƠwx��
�g�����qν��7U+u��U=�;m��vtU�͹�Y����靽3b�M�ܹH��
�ԭqϔM;�&����NA=һ���-e_L�K��\��u	l�񈿵.��7}S���b_,��R��n"�g4Wj��C�s�>߲I�w��-c��R�~c0�����v����z�R�;#}5�|�Rث�c�f�{e�T�� v�:r���v�G��T-���aWy��j}�Sn�G9���g"�{=ܳ!D�G�ۘ�`^��Hw�j$��~�*�c�Ǿ'ҁ�!�#����[�-3�8�v�{%���,��V|ϑ�E�~=�x��1�Ί�<��̱�G6�+0J��T��=�����D�}Q�W�ms3%�qz�
��ѝ֙�9�Y�ưvv��WV��o�&��BR��S���ݝ�:�s�n:������'G��n苍���b.�X ̳Pe�Z�Bz��=�!�;���BT?mO��/���h��yFx�����Z-XJsb�C]�Ztq��>�z��@[9�/�5��}o�>X�Om;�}���ٟE�N`k}����^^_o6j�q>cw���G��ӱ�o�����t���(W���Ȧ���(Wީ$��W̟��u+x�]<�:+�W1�j�D'w畋m)���۝�_k�@�zdY�AI�J��vH�̧��<��i��їõ��j�U�ކ/1p}J�IG:dB��Z���Պv�w=�Gk�UC�N��⹱�n'��U�ǻ#��q�Ƨq,�ߗ¾ɜ�d����3ʪ�o{����+���<]�l,���=��A�Wp�]Ɲ����S5��X��0֬���1S>��ߊv�𭈼�R8�S�a��5�C����#�#�4��M�?=�s����.'�������?v!ls7'���GP���Ժ���<�&�橞�����<;Ƚ���|A��Dϕ����=5��Ԯ\��t�tc�%���up5Y�-�)��o&���#R�ޱ��K��^Tkv���Da�ѻ}���b�ɸ��Lp��l��?7���O?OP_5�^�����}dfl����wg�q7}3���t�z+Mg�pV~������/��ds�'�S*��������s�xD���MľC[���Oy�k���������Y�!�ˈz�p[��xl�U���DE-R:�sZ��>�C�l}=,j�+��^�=��p�F���MB�T+�+�������b��J�|Ѿ�]Ь���=����,�{O�/�ڽ#â;��Ru�߹Z�(*�x̣C��s68��>=�M:���%ui�бTI�s��K�s;�~����21�ԶpT��r�t�Իq[�ű��]�;�i��.zz���:�rYD0��-]���â����J���cb��]n�?7��;V�2�� �c;&t�ɨ�V7�֕�ط���|�����Op����|D�C{�8�Ք.X��|�����v�2���jۘ�)�;}��М��r5��@3��N�wWLm���S���q^��g��]1A���3"�[�sm$&��wN:ژv+2�h�}�ՖO��wX�R�s-�c�X��3�&~Ӌ���\��D}{�����Avf��y�ŎNȞ�U"D���+�2;K� �w���uwm�eX�[ gl��ӻ4w��������H+�*�}?uT/t6����v�ǳ�;ɱ\P�F}���p�܃�roh��^�h�h�9�ۈ�n�U�Q錒1�]f��:��[Z"C�Ɏ3��X��wCª��`Ғ��]�Qr��J!���;�l��qz
�0���D��q�.�EuVj�[J4�iå�D+��֜v"��f���;I�RR�6,�ʾ,	��d����:���Nc��gg�)��Uo@�t���a9�|�'�X�
��E�h{>-L�߇�7����wN�T�Ɵ�{[R���ݮ�[�Ju��XD\s�f'9{�lFc顃3�cL�q.tǖ^
$�g�^	n=���,�p�T���VX��]��U�t�;K���3��OX��nf4|66��:��]o���Wݹ��qb��8n*�T=
�w�&����Z+T�k]��S��_�x,d������T�u��J��&�t�![B���9�ղ�(��}*󄓱L0u)�^=�$EF_��NLŖ���+�Ҧ�Mfm�fNe�#�v]>=��BU��H�`n	�c�ħ4�Ew\]:y)�W��mU<qB��f+�^�R�{f�R?.��g�7W��o��=�C�OF�/*~�}Ud�d�'��""��t�l�P^C�Fe��ýأb�R�;g�ۋ[�T5Cx�q{��aW_�8��T��PٯDv<4�O�ӿ*ۿ�!��ϖ��=�G����C�t�qkj`ק�e)�@p�\��漯vTz�A�[��ͽ^ϔ!1�ߪ��-��wa�q��5m}E�I�L���h�7f+����z�uE�2<���˂b1x//k����F�����42��צ9z�w,�B�	]Lmt��W%�h��yONw�E#�7�\��>�����x]���������5�"��OQ�Q�Wr�!]\缨�c��#�I}�,Y}t �;��?{c��3�5�f�\��0��ǹ�8J��k*�J�Tn׫
���^UI�o)�NB��=S��3Wݱ<<:�֠s�<|s���̕���X���{)�&���-�ފ��o��U�%&����|�c6ڽ�)��D�8�wb���E���1"����¬@����Q���N�Q+���!X�xa�h6�G�2����WFj�a��[Ԅw�'nԬ_�s3-���6�_�{q-m��	έ�א�yM-����х֑u�-���X�1�""�f�뵕,ou��L���5b�� �w��a)$� ���
:�6F4es9.���\A޹WZ��������{�d��ؗ�����\���+��E��O��)V�6f#��-���{ K$��ޤ�I�c�!F�"�T�y�b�gwmb4|n�d�w�\>���?��ۃ&:��׹����r�S0L,w�p����s��9��%(�9��z�z�+���/�ߧ�nn��س�n$ϑ����S�����¸r��}���Nϣ��Ln�𞮑e,�E���?����΃��� �>��ɂ9�L���3/��K��mz�)ZO]�N"}��X�{�n���V��Q��g��鍨g��>z}��Q�7=�s�k�W���#|��\��ͼ�sW�+:C)���U��ǣ�#g9a�$Ɨ9�k��'����~6�Y�gR_h�6��2�pNߧʊ�������"�Gr��D3���>��qҫ7��3��{ Fug�(I6s��BIH�A
��H�ݝk�}j��縚�K,$�=��H�8c�.�u(z|G��)ɤ=�C��s��eEَ�$>�Axf�Vzwb={4CW��v�^&��щ�V��#�M���K�?�����G4*�k�tb�Y�Л�+G��U��r�=EP�ח�A���D�Cr�Px�5��]"˷\�r���x�l�6��2�g]�uΚ[�q[��v8o�.���d�e��?oH�}�&a�&�Y'XMۼ�vލ�o'�q�
<r�w��4�	F�Y~��U}Ku��Qg�������o1���UI��,/�_��U�O�O�a��
��3:t��xz/��R�t�&**��K�u�Ȏ���t�W��S��ws�Ҭ7�̉���8(��R�JU��������=g�ɭ�;�\7��&��Gܭ�|��h�;+��wNgdz"z������咼����:�t�/�,<��w��Ƞ�"(�"�O��.���w֫��VW��"74����T��<�Ip��oE���W��p��|E����qMRQ]��w�f���Q[a�ˏ+6��z�s�2yC�bp�C��U;�+��*���˽����s=]�:�?aYAm�N�;�c_�*TksU���Ff6���	�����b�g:���K8������9N{�^���$�U]�7��)���Զ$���EZ��k?+�2�~�Ŷ�G��޷Aq���h8�V�Χ׭x�m���n�<�����Zu���.�ʨa7F�D��{��(��\r|^������f��o�����^����8�ь��B��r���E��J.�����A1����`֡�8G���?��Tβli]��{�Ҷ��4��7�G$l��S�V�[�xc��1�܈�u���W+0`�t��c�9i��u�N��{�ȫ=�Ŕ��]�<L���[d�hl��d]j5���s�ɒ	p�0��uoz�0jm_V.����V�gj�X+i���,�J���T�O���n�V�mk��ܛ��
P��|�p\�2�JêX�ZX�\��מ�h�Yչjl���-��L9�������n*Y0�V����Q|�g5g"�yʽ����rKY�*�*]��e�]K7v�A���'�1S3(�M�MVuL�3k0�o1"�� ��wLq��=W�;8ՁH{Ћ�Y��j��	��(�cXF�U�#򩮆�\���C
�A�3;I�S��sq�y�l]Y��q�V���wF��u�<OR6�rȀ�)]�U���L_V�Et>�"�:��*=H-cmT˸�sL|�k�uc@����N����,��׽ӷq౹oj�O�l�u�+�p���R����0�8ܲt��6ۤ:Wr��@`Hr�Sɉ�'f8r��;w���ZSD[c�p���EN��(�/�z�\����O�mI��YQu+�o�&���Й���&ř|O# mm�D��$�yi�㷲�J�>�s8-�<t[v-�ߦ�1S<(�rc�xk+��X�+{�_
��[h��}�jy�w�j�v�ס1Ly�C���T_�r��fa�g>8*avTv���G���M�tg%��$����wC�����	�9�����	��XN���v��W��yN��k��lDn��xU�d~�w�:v�F���vT�gl7�iVfN�
\:<]�%�:�j�l[[�ގJ���v�>!T��ލ�}��Ք�Jޢ��*��u"���g.���#�Y;̍m�R/dt���W閳���wq	�����Vᮢ7+�:��Db�S�E�<�Z���ePw[a1�:��m5��䏃v���yej��T��t����]��)t��Tű�.[f���@8��2��jem��2�BV��Yæe١b��˴븬��W�Sj�ѶE&n�N��i{�u��7��Բe�h_�M�{���Q3����PO(�4������O�X(�׏Y����sko�^��Nw<+�/N;�cf
��ǽO��Ic wn[���62�c��B|��.a��I�ˊ�]�u�]��)��2��nf�z���1���C�XԳ��ieen�Mo&��6�h�1�T-�R:�y�"u=ו@f��՛��X]ms�$S.#v�vaGQ�v��&"��u]�^�I^q�`�)�8����5X�rB=:�k��a�.���C.[L�u�5(	r�&�8��2ѾV=�K��w�����7�Px������U�|ϖ�� 7fh�{3;����NV��j���6d}�I)��L��no6kJr�6[ɳ�u�ݕ��]���12���f�[K��ޜ��ϸZ�������j�������[�ޡ-[�{��N��(�e`�u�RD�=��b��9�tR��$�?V�;�5
^t�ޖ��л�7��p!�,����/W����O&��x��E�>rfFlr�{�@�yߢ}���%�}�'��.��g՜:k�^d���#��`ma�:'����p��ZSR1z�����V]t��>����#�*�`�S���؎vf}7��kyoR��{կ���}N�}k+�~�t���K~Eg��N_�Ē�����p��.6����v�ڿ��Uw)��[E}Xͷ�Hl{b���Һ��~�b����Ns&��5q���)2N�yi��\>:&T�Q��{�,T	�q�qXDv?�/�JO�$�ǩ�3^���4��!�ɯ��/~�cqNN@�^B�])�K��L�)dpBա�{[�۟m���tK���R��\Oin򇪨���ΤZ���i񘗇ǲ\K|�o4�+;j�B=�c��L��A��qb�V�zC�>�/;F��-]o�L��@�����)����ޘ�<9j��u���Fp&�V���W�����{�4�ϟr�ux߮6��'|uXʟ`5/K�[ק&�e�߹F��쎜.{�O��+"!���b�`C��3Cv�����o��ZS�`�+.��/UD�Z���Z3�d�I����ht(�n���e����<���]#[�4�L���-�d�v�i�2S�Noz�g����P=�Vv�oD{[uE�T���7��I�l��m����t�ӗ��m9�o{zqEn��WT����!H�����4�
frrpFp�٫��7��d���~'҉��⵵��Lp1@wN��Ӻ�BW�����'�<��uh�m�;{<MT��~��|b��.e-�;�k�<�(�S}��q� ~���Rz�na��1�5����'ގ&f5�TL��𕛛�f��n3�D{j��
����z���#���o�t��:��,��ѧ*F�K߅,��f,���_zM� �u�N��ׯ�ɘ�;U���C�6%d7������e���q��~�#�.J���⫟g���I��N��OmP�|j�ۊTB��A�]F28���T�מ=B.v��8ۓ�:#�;K�T:��$��'6��/y�Pn��`��R�Nf�W�:�>�;4v�e=FV�i�.nq�vub�7L����R�7;�EP��������'W��РS�s ڳk�G�2��ǚy�*�����B����;Π�5�uSɐ��wGn\��F��Hxq���M]�M0&�ّ�ga�{����'��r�k&KQ���G�Q<ӌ��2k炠��ٕ	Mp�^������m�9T�S�`PBŉ�N�����D̲:e�s��_0��2�Op:�¯�R:2m,5:�Z�Bt�Z��sU�6���u; �[Ī���X���]	�wwK���E�Jɮ�
j��9��Sٽ@5�{���{�y��[7:W��^��,�!'x��?}�ܖ �t��*d���ף�Z���6Zr�]�M���Ve�6�/�Y[���;��V��O"��>
cJ�W��IW�v��<.4�.eɳ��".g��!�}D�VDs���_Ɖ�1�r�8&%��ՂRe���jM�Ya5���O�|�7�V�'�������͚��ٕT}=�uN6D���=Y���d�I�6�s�t6�Tj�V�v3�T�*���8=���+��ok:�����[�=�a"= _w�zP@ǣ��Xe�Z�'B����L��}@���t/���y&�O�9�kSz��v+��̇��W�]*ǉ���z;�_�3���m x|k�_t$����o�1�1��{�;OO��ٗ$ˮxr�.]dw]/�g�:W\�=����VO�2eA���W�w�*Sp�o��<4wg]f��5��B6X���G�;ѝKg�!S��&}_	���ܺ��&�r���}��w1૾�\g�!�~�s��Q��Ʒ�mk��h��-UA����	:=�)�˫5�~�g眞~�8y�����ۮ��2��F����#�t3�6�R�\�nw��	�+�Ѽ��N�#�0��D#hN����ou_r�^S{��w�5�phk�;k,=4:�W���;�)�,��v⣽nb6��R�v~H ����`86�e�ꎠ�"o�ޭ2�Yk�*V����Y��+`7���>f�I����{��<Nzcוp�f��&�\�N⭚�s�	�q8n;.ؼ�Oa�](gv�z"���4ky��z��i��uXcë�A�!�]W&pC���ёh�ܴn2���FR��{���ၙ��='s�O�;:�wܗeP�Z5����P���Rg�A�g���ӷ�/}JC�z-73������T���:��ܠ�yq�����.�j�~!��P��6���j�ɫ�)���]C}�wi$�{'�d�j'��;m- a�q�rDE��m�HP�%
��{Q>kG�����w�㎎��<��;��G.��~����Q�E�}s'�x50�~�\pH��>�����{_��Êr�yj2�8�1?g2r��>�}ÿ�נ�:ؙ�(H�f��; Wg_CP�$_^��wyae���9L�Nhf�c�t��yB�W��㞭��#fGzT��Ժ蠤����~a�ND��^�YV�H/GX��X6���蘺}ٞ'h��5ǉ~�Q��]��{��^��uI�=�Ѻ��mu��Ə���J.���ti��S�fݴBi TvD����{C�H�UZo��:��k�U�5K�)�X�w��gݕ�$Y���o�3�I}�vӷԠ���Y�VU��jتs��^(�8�ܦ.Y�=�ô��/2W���	�K2��oA��w]�"��nP��ɔz��R9�>�����gX}-]�/��cA���
G��[[����Ϙ�֭�XXk>�q.�/5}��́�9>����]�H��������(�o{<&�/��s�{-�z���>2|-*��>���I����;\V_����3�H�_x���8�ύ��@���^e���\U�>�+՜(Ϻ8iqZ�Tm^W��� �/�}�i���eR�����y$�ί}�����.~W"�}�%���3���z�s���d��uX!w�����m����_��M��D�z�@�sT�⺿t�͏F%Q���j7��T�s����X���W��4����m��{�k�&�/)�Hx/OL��G�r07�z�\'�}�z�c��u7��J#f�Xā��S�Z���#�����K��PK뽊 >�WӾ���G���h\{R����)m�7�5��IL�Yt��=���Tt��<�pℝ��h��/�y:-JЍI�UY�s볶�4?��[���ԃ����L��>��HQ���f�!+��Q�",��r ��w����}:��e|��MO��������ٜ9��t7��ZpW2^\0�GH�M3)IB����ܦ�P�d�v�%�o,KM�rVo�v&g�˹"sf)B��r�ѥ�`6�Ub&��7t0��V�|B���{uזA�d�*�j�%�;Xjۖ�9:����>y��	����E��j=v�����L�Ļ�L����;�)dS�?D`5�s_\哮�!����W���9��#h��芲��W�J��%'>�>����!l�d,��������V�z��7�����^�K�KUG����c�]6�o<v{�ub����<��I~���٫�B�{�����0c�����Q|1@'�W��L��߽���05G<��h�Cuo'Fxn���aX�
_`�L���>r������?Y��Q3X��xM�C�ׯ�;M�T���zxe�j��T�~�0e��|3�.u�S���E����'rbE@�IϦ`������@��w����բ����Gf v��RH*�֊�������^�Ѻg��r����JT[��ӽ�1�u���3�v�fo����[������0�.qt6Dt�m�c^Fg�[f8G�M��3ї���JΓƹ�4c3��q�"r�U�YqucԮ����u����&Vx�\)>!�!n��E�s+��γ�~���d���Dw���*k����q�����S�;^���r��s����E��=�D��)��Q��gf���;�E�N��a�8C�"���#,����ȱ[�_sfZ�luf�خ���A]ԟs��*����p�9Z;��w�����c ż�����Soc�}���J�ph}�͔�ڝ����"��+�k�(h�E�eKmNZ�5��;]<��h�����2m{�6M'H�Og�Hq\b�6"=�[�ĺ �ۣ�t�>�\./�5s�l��5��FCs�V�d�A�b,���u��ybI�ט��"�-梗>�O%Z�zx�3�`�J�{6��ͣ�7��i�,��F�u�X���I\�D�O�z:�������Ҁ��l��I��3(�.���W{�����%;���K�vA�-��*����k��w��M�!�"���iE<>�
:���9�ᝋ~޷��9j�s�t��Y�Y��ʝ���6܎;Ȉٵ�X�3ΌPzS��=���YM8ss׻�1��y�ū�7�#�'Ӿ��z�a�VoW@�+\m�"��	Χ�W�ߴ�>��㯳��|�|�DC�X��*�1Zr�(N4�=�6�;U�/B��Ц"��e<�x��'�*<9���aX��r�F+�E�7���ӕ�H
�q�t��F^��rdI�~E������ȷJ{��8��9�𻩏����6{T{�z0��L�W+�݊<hʳ�_B��qa3��^�Θ��4{��]7�Q�ݟ4�)=ή�Ǜ!CQnw^U-�p�-qt���xP;(>�'9���i�vb��7���f��|�b�ݪ��S:�G�&��ޱ�?����,���%�:_m�[��j��+$n����*:�/o� a+���7�6�Y@Ѯ�tT嗩❜�BcY�r�o@�a�Y�~Ak��[�o��܁9�� /U_m�Q����qI���k� �ޟ+��{�`���b�n��m��z�q�7)��5Ns�PuJgý�钆ٹ���$�c�]I��m�X._����}Ӿy��d��t��ݟ��*�����%�$F5ۿ1���x�^#>���vY�1�޽BG���d���Z���z8C�w��W���f�m��h127L�sts�������Mz�p��?�.����1}�KӲ�a�~�T�O��c��+6�G]{>���7��u?�^�#�J�l��Z��ŋJ��R�1w���eF:�bT�u�O�g����M��meS�/hbx_��6P>^M:�VV�D��3�<.��|��q{�Q���{~�N��w@�薵s�D"�1gp�{�׬��I��#��:��5?H�qnZ6�������_��3����3�\��42&�"�U%PYM�E�ա�����sC���^��+ܯ��u>�;�ތ��|�sѾ4�Z�v\�(8�����ZTM,A[󭬧G�q�g�}It�&�7n��/�҂��6&�gs3+\W
��~��[T��J'H�(���J�l�s�*&%�� �U.�I[��᳗Վ��S}������<��fʐڍ"ʾ,�������.d�{�ٻ�d����
�uw>�]%���﷫q:��P=N5�6����T�8_�c�����\�14��o"�Ί�,ӷ����!��SQ3p��\O���~߉hߡ�q�����0_+�Z-��")�W��ް�37o���S��Aދ{ٚZ5�S��Wd0��6q3�Xà=7����sR�����^i�S`�>�u[Tz�b;[�Զ��|EwtW>7_sc�R�\��P�?����Of���M^G���o*m�:�{��*Y��J�w��ؓ�u�I2�7��W+���漌[�e��J��_i�v�ѭ���+������U�$6��h_��>Qߎ7;��c�R��]��z�Ĺ�Ӳ�����;7���=P��>�u6;ë3.��0�꺘�~����� zm�˯@�9]�CJ�6�{�c����6�J��]�uɰ��/Te(�e��_[�<,�zd�# ��yeZ�.0��ks)E�ۻ�i���%=��P�i�_~�;:��k��몞5��7���tN�c�^�}K��62XӴ�<��t1�|���5"�N�oq7���Q��
�c�m:۩Q�ui��>Gi�Y�/^9{��<�[�e��:LE���@���S�Z�/����� ˜Ht��
A�X[�����f����F�����4lps�歘���Oo<z0�&54����%�'���Z���5��1ȯ�
��˶�׫WQ��P��|�՛аA���l��H_�=t ��k�Nnd�@�[w6(ճdG6�����L�^t��ǳd�%׷���B��r/j��F#���q�>-����o;ReƏ��#�;�D��	��O���7�Ag���mv��������D8�$8��h,��yܖg���~[����b2:�yr��E^\w����=���=����7��ak���>�f�B+᏾j��{}�v흍П3��տ
L�$�����:��z�����*��mɊ+TH�V��*#��U{�[�Ml�gZ��������J���_�-�v%�΀Z��Ex���<#���Llה�l��������<��`��X���7l7��Z��U�(NW˪3�n�p�5J�5��{��=�K���mZ���Q�3��ͫ�3�yߍhH�T�\����/�����}���U3<�F�}#q����H0����~y�$��=�f��GLw8���\n�+�;W=�ӹ01?mx��))=ݹh��&���Za���MO���sc���d���9��_R�v{��l}��4����r�]�y�7��p�R�z�����34�B�Gu:vqM�qښ��B���>C�}�t'�����H4��S�B;���e��1�ΓOL�K��>�{��Ǩ�麸��d�k�o����Y�����'/X���h���0�!�͞���&��Q�H�,��pk���Gj�K������~W�/-��z
�'ه���˪ �,GU�u�b��c,���b���i�����sΛ��$@�5��(l7������1�}��\�v��ٲc{7�o:/^�-�Sept2tbV>&핹uy��M��N�
�,��ȝ����v�n�&�5q>�6��\�V�X��!��懬V���T�$�^Bpc�=�r��%���(��ܗ�Ө����ƺA[A�CxCo8	Ic�����ۻ��-����z�M�a��V�}D�2��ї�][�6; �0�2�N^En��zr謊]�Wq��YD����э�L�����N���#ۺw14�u\�{��i�w:�U�����+���	�\�X.�sf~i'E2�d�:�MZl���oc����[�:/�g9c� փ�F�N}��y���=��eu��#N����l�U��+�u�b˩v�g��,Kܷ@�)k:����f+3�*�T�h��n��r$�;�G�4��ݼ��������L�Ԉ�n�Ӈ�����U��,������j��Ŧ(���"���M�or5}�@]��J����q@1�v�X�NM���~J��n&wËy��Ӻ yhƥ��F?��V�D=���oV�Y�)��h��u�۠o,
Nz�%�3FfM��"]	�f#sy�}�/MJV.�e��
<d�f�$
QC(CԆ&W"1
��ܭ��z�m6���L]et���gz��_X���`��sD�����5�����Uf������7算�`�.yT*��Z��K'U��yY�ȷ�����CEԤ�}\��k�n�ɝkc����+���';����_4�9*Z7h��C�U��&G�]�.�kN��[�,F���w:�Qd�9VM<�YA�\��)����ݝiYA�ep�ʾ[�V�2j���ά�Ŕ�U��ﳜը��*H�� W黎v#�H��a���˔Ͷ�	�A1�f��u�R��Is�Nd�S��i[�hɆ��LZ���x+����٭�v:�ܣ,t;)�q��^L����ʌhx1+ԥ5����e:8E�Ի��چ��ػ�ݞ�iQZ�yX̏�"X�w\��Cg#�\&U�/3d�bΗ7C���7^��7��hnV#�:�ڥ
�8^f���}z|�	�u���ם���)|N�a�4v��!����������:�c/c.�g��w.P&4�$���7���9v-�W�Y4���/��k�zi8�#r�֢��(dO.�_d�)������$(����8�1���3�ӎ���y�W�ɜ�D�^��#8J�8i�=ʺ�9�ٝvv���6^h��8�q��cӹ�V�;5�쪝��V��u����d��&�&�����x�7hl�t��z`�4zk�������dR� ��/�q��`��Pwl
�^m��H���C�ʾ���Td>-�oHWζ!��~��9�;2/�}��*�B���������B|�7���U�z�S�����dg�|P�A����Lߜ�O��9��\Pz�r`�*�:�d�k�+����&=��)�&aJdwBə���,����C*�{��gr���	{L-܇���yQu#'����Ma؎'�m��|;��`�Q3��]͎��aH�����ƫV��*x�[E�9\q^숂�DH˷��;���t,w�4��rrҋ��&��{���9�xp*G�+Q�ו5���w��A���ޭ�y��2���'u����C����˟8�ed��Y�&p�,E6�w)DX��
��h�}���:3���8��U#�ǣcFk3� ��zȕ�T����̍~X(���Y�u�t�_n�K�
��5�]�3sY���t���nW�.�9;����%=[~���w����/}��1k���wP���`���o3��[�b.���׹ i�=���tt�{����g,�D[�	��T�6��j�|�#�����g��	?L�|tyZ���f���|����Y��5�����G��\���ێF�.��v�F;S�%�e�����L�\�5H���s��;d����o���Nʒ��6�����z�n�	����K�ȹ^�Û->xn�M��*��;g.1��f�}�^J�����,�x���dg�2f�v��`;���߭���`��n�\���A)�<��ӌ�r���|E�&���Õs�Py��+�]΢�d;�^��}|	�`L�s�x�C�{+:�iWg�\��{k�&��0���D�p��w�欼��Ta��Ǚ�%_a�N	��&{Qn*��ݜ/󻱭y���z���Z��s%ͳ��4�>�w`o�5t6?�A�������w�SǱq���3�7k&t⊔ɌRut�]J%Q����?���Z����rj�C��w��	����1�	���`u�'�v��}��`�����@`�n��Iy�\�t>�y���c�M}��L�e#��q��iV��ē�)��9�����~�/Ȗ(~C �U.��S�	�m��8�y3]�UB>��{�jٲ��'P���Q87K�co�38�u�S��;IX�U����.�L�uS��yٺ-q���-W��8T��9�n�3C+�*�=��+�E����U�'̒u���҉yq�o ��Q�%N�
��C[�H�9L_��/���+7d�n��|r���$W��t����ǲ��Dfm����o��YmX��j�ItSd�D�Fv��7�Rv�COna�R�U{]�܌wu�6�7��f��
 ��cS���wpܢ���	�[�,�ްKtC-_�
�|�X,�o����߼���a�9Ƕ$���W��_od5��c��)ȶ�_d�t*�����D�38+z�)��wI(�EίUL��0Q����I��<�ϸ�p̞U��4'���
����)��#���
ߟ�Z5LرU��k�P6qn>؇3������r(�9�ٛ����ja�W[���p�c�V��E�\�7�ܞw�0����=���z�}k&�lT�<z=}��\�6���{����D�WZ�)�+�%\&C�h怕#[�$ɪ�3B��M+È�Dt���ԴM���'��QX�����»�^�>�u�mU;��yR{NV��:�q�G�>����xEN��B9p5�>WN����>�1������+�T��y+t9{��q5Oj�:���j���͉� W�̚�Ԏ�ڽ1"{�1���r�"Lfd�K�h���&b|��}��u��̀O�Ǻ���ܲ�o��w{��=��%j�cj�Q���S=����n_C��Y���g��7߉���؅�R�a��/+�ZRw����^�0�6�"|ɞ�SQ;YsXj�=��{n5�#p�ê&`>C��<g��b�~[{���ɖ!34�k6�L�N���wݮ@JO��Q���r�q�V7z��eǱ,���F��E&By�@��kT�$�{��w�-��#n>2�Ӵ�m�vm&�T�m�nv�O���(+�5m���/��sK���nPD�b�fw)�֧�u�u�|�3P�B��
|B�����i����k�7���'�fJ_!f�}�o�����s�UKؔ.�s�30)	���~�`�g\��q��wC^�O �IJF�j���:N�b����.�t���t�l-3A�^!;$ֽ��uQ�kz��Wa3pOhr�>c/���� A<%�gZ��>�Z}�!��s��s�)s��r�'@y���"k�3���S�A.�U)�6`�n�Ȃ�3kZ��Z&�-fr3�@���!���f!����b�l!�N��x2���;�:U�i�r���+l\f�:��)�~����;THC�L�/���|B�}����:�-�T��/2�B=Y���b�����a{�m��a����\�r:�e�)�]��t���Ř.-T �{�>�3.�;a��g'-�E�Z����W3xCT��{]�ڣ޾�D�t�~P�L�T��=#���"���d���;1Cm�t@�N��jS�j�b�Z��y�}�F����>�"��<��*�'e���������{���\cu�R�a��C��*v���a�s�Y��aY󚐵�Ҭ1>�ao�Ы�j�r�g.�����d��ۗƏ�[$���O�㮢q"{�L����HM�u8�8�0����S�ym�P�+W������E���t�e���bv��LoYzj�Wv���EwzZ��r�S�\��sX��Ti����{�n࿤���@���'lmK�K=~�})���䪨�z�yA;Gh/�]2|�x�췺��	�34q�t�kj��,��fm�'n'o,LBU�/����H��a
��q;~�}�-cx�����⭼��9�����j®����!�O��(�ٽ���:�g�Jr\�ŕn��E�������@�ѹ�Ea���>�{�>�t�¢�<�vgf<��~o����G�6�0W��T��y��/�}��`L;}`_�$
!���_U��s��~�r@z��:������9<����W��"3��*�Y�Ѿ�����r���1n&<Vrg�Tw�������5���sR�^��Lߖ�%�p��}+��K��
��>����	�*�:u̢��xB��M�̧ڃ��Eo�$C=��1<�3����5_�:]�j�{�e�����P�\�ؘ�wM����;�ĉ���W�����(>ʳ瞖;I���P��6e(��a"�u	��������+��D����Eͩ�ECK.�����8}���^uWdQ9��-=�a:���Pښ,Ӏ��ї0Y^�3���!C�ƞ#+9�J�hˮ	T����z�wh�P(���ۓL6���_ob[F�8�N��1�M�M&�B-L���;jCZ�e+yD�d^��0$�hB6��n�g�ME+#8�OyX�3��	�H�!n�qKoh�7�Ud1�&:�LWG�]�	���cǻ{���T���tx�?�ʏ��\�vb�Y^ 4�����Z��L�ݔ+�t)��
�.]�Zj�`��C2���%����v���.� ��'�:7�=&N��)��g�ŌEn�|����;�Rh�������9�mȋ�����5��X��*v�"�ٳ�aF)ױn��t��ϡ�����Ke�Y�׌כ}�����ӊȀ3�WE�1�0f2�2x�g}�(��Op�DL��go��]��S��;�
�l���w�0����}.yxTM�Y.�ky���˺�|����G��
j��)m�+4�=܇p�h;���D:P��̢MN�j,_G�%yR;��8+;�GH��!���P��+g{`��0�K�Z�Î���v#���uf3�����N����p�n�5>j�H]��U]xx�m���b�VU�e���:D�9�c��vzex��K����B�ۭ�V�w���pj������w�,̽P��8��t��Aܨ�m�t�i=�B]*�4�~�<�{��dP.��~��v�l1���R�ݝ�h���À�0�EPW<�a`�M�=J�Mݻ��������81e7�y�wհ���̆�k
Ja��v��gtuq��J��Ȇj��B.�]�	��x�y&R���M����Pj$��u�f=�o�b�kPu����4wixt!�o%���,���~��By8vY�s|��o�yf�Z�kqvo��ǆ�j�Ϸ�J�L�L�fO����i-eoײ�,?K5����5ڗ�Or՗q��-R;@����C�{sE�pe���t޹*�X��^#�W���`*�4�_�:^dv�.9�^�j���}K] :�u�@2�j;�k$��[�P�B��� u����vk�Z�Ԅ%�j~Vu*��π2T���!��6n<�0.Xq=��M�Ό�*^��o�dk���T��Ù{��O�LwZE�O}=t."y�6`x>�0�>�}o��U|c+������p�z:����rL�~�:�ʷ�`�̽�d�>���s���C{ɬDZ}�z�<���m��g��>��ى�+�C�VP�c�18�8=��t�%��Ӯ>�@Y����f���Q,�n��}Ɲ�mφ�7�Y>[��wpU���z[�*�%r�$�(L�9>��{�=\�=��W���U������n��`'�
��Z�Mu���OGi�D�|e��ȺO.ny�g�1Aޡ1pܓ���W�kM���Bz��f�8Ю�-F�ӵ����L&ձ,��;��$Ѫ�2)��c�W����1u@1�Fҹ41���[ѧO��ی,���Zq��Rg��I�ǀl��a^X�]�[�ʣ���4e��m�%b���N�u�m�k�ط��-h��x�⣕|�G�X�Ss&lJ�����\K؋��M=sWœ����-�}�+���Q D˼�3��A�c��V��j
���h��>�>�{�%e<S]NwF�l��?�����Ͻ8>�:p*�K\W��ϯ\k��@~ք���p\����N]��T��u��1��nF����7�c�D�ߠ����rW�
�����8{2���ך��0�8�I����"Dz}UVR嗘�9{U%���cW��K�<����97��ƛ�d�SD뿡��^�����F_,S���{��I؎�zFLB3��)��܌�|d�z"�I��]�S����$)��禽�^c1_�{�o-y�T��3�KG:���Y��ؾ���[�����|J��>�}=5��$NULO���j9��&��!b�y9��Y�zdun�p@>.�'���s�x�Tɽ�d먏I�����w��N�����n���XQ(l�x���<;Ll��V��j��8�_���!�hu$cnR���g&�Q�����2���#�`���U8ν�����\.�+�;6��=��z�Q6�'{(RU��$�&=ϩ�(00JĪ���WJ�X��4&*�ՠ�����W��rI��*�2�>�riN�Mz%~7x��P�]�vv��R��]�i�j�Y�Q�s]���wh|�%e��aef�Hg����(Z��)`ҫ�|�ql�`^�Dw�u�P�N��Dh]q|���g�L�N�������6�n^hYf�;y����7�eA��!#Y�x�6����u+�;�V]G]j����%��f�
Y��؈A7�G�K��
�>�91��e��py�
9J �����Q����x}�jf)���*��<U�G�WT�6�_��緣<�0�>�'��5/|�w�{���֝������&(����ی;��u[}� 鲞��7�qW�]a�٧S��-�����:ju����}I�7�M#&�N�嚔*��R7�3�f��Ϲ�r����ӥD�P�Ӫ��>�������v$�/wIs�K5��2OT�w���+�6���p�}�e��4�G7?�<�ܮ�}ٹ��CV�������T;��l����Tc��/8���L��z^���v*)��:�+�6��{��ܝ��}܊�{���]
�����G�d7c+��C���
��%��8)�={>Tw��ʌ�ސ���W��K���?��S�u|���x�G�~?h�?_�x��YXFB^��tM�^O�o]�o@t�LI{Dl��ү��X�O�^�tqh�z�HV��U�"�JU�0�u��Ҭ��G�QM����ӫ'���L�����\�C���������^`��t.��R�6�Œr���m��v�o]��θ+����"�w���g�j!�.v����h��m��.'���E�\�8��`&rO��X���N��Di����=������T�Mun�uh��Ol��XqqSUl�o�*v��٩C��$|,�;V���t��ڪt$剸�퀯K�8߯�9��+�[6-�7��ð����C^?���9��N��G~Zh���������<�*�A����w�x�𙈞E���}˥a����B�nw��$��!��&1(ڝᴷ�D*Yv*Q�At�����/}�6�Yx�Xb|��׍,�a�+,I�Kwd^���4bH��t�>��u�{1�bMD��K4����G��`���OW�����J��F���у��Y�^s'�^���J-�ą��3�S�SC=dA5~�3��s���.�j�%T��I�*_H�m�G�'�xd�ß��@�:g)\�b��x��b>��C�Q�<������"2O\���9����^�x%��T���G�>��s�2�=��͊��됩�i�*�]��TK�7~>��'�����ׅ����!Y~��vH��7����_}&J}��U�s��q�K�t����Ү�ዖ��)u{3�=�H�[Y�m�=�c�١ s�5BP���+b�٣�J�+M���ù]�\��XK76�p��Ш��F��I�YSV1ңMX�h����۳](�Q�ͥ�(M�Ӓ�.m�]����ar�ø����&����k�:�ʦ����W<gA�d�6�9N� T��Ab��Ix�k%�a�v������q,�R���Z����N��n�.�]yu(���`�Rs�7�C(�17,'ϖΖ��s9�C��]�k7���Wf~�
"j���;Y�lUu+��A��=�n�\��<r�Wj����a�u�Gg�`�z�Qa��u�|��6��ݷ��aw)��{]�z4�Tw��u��a�=�*�og'*v�q-��o@�?�'b7p�{+���ziӛX������m.��/5��z��͇�⍹���H8[h�b�T(�C5�ʥ�nlI�z�֐:�c��w��H=��u�y;4�
�����qb�{��p���9�&;��!�W��b�Ƴu��@�M�"M��^;gJ���ahۢ�-Ԭ�+�Qa��HT५���靔&����6TL�i���n�mg+��t�/P�heb+8'7[�h�p��g;�I��s=bR��S�;���ge
�d�H1�Ɣ�W��I����!$r}v��T�B��w2��lq��`|��.�K��9�)ƈ��d;X5�h+���f��wt�MwE���-\\��#2��!l*,��d�fp3Yͼ�۵�OG&�Jz��b̘K�N)̓�x	'��$h˂���:����t���Ρr�3%��!�fY���f-��:EQԆеy���.�M��|Ԯ��k���W���Gހ"a�9��#*'����ݤ�JV�J�3 }R�(r
��{\�B����TC��(dꊠ0��L��:�Z\x�b����x�ڮ�c*��-��y��G7���[�.���WN˽<���鈳�eQ��wlfn�����NWB�����f�L�c���/���4le�D��3X�/s�\�pR�C6�Yҫ��H�hj������V��([�~�n*�֪(+C�<�漙�(+���m�:�;�aŻ)S���ḻ��*��3�e�',�me����%�0��N��6cVr��:�'PV<ǯ.C�>�:�c�x�v���!�f!��������^6p�}+�1�nѹnv
�s�qZ�����O���Ճ�����2���d�B��ȯ+'<��LL����*�ɾ�)i�P�9�;��pk��@ib6xFR�O��R|�xJ�;h�}2n�������=�H��{Z{K�݁�=}�O$�j�v^�=�MGi��>x!V����&�}t��V�$5w������6����7D�h��xĀ;�RWZ�M�P��U�!B��ٯ�+L;6[��f�/�m<"��\��w�	�%=��Drstv3@ ��5t���,��w9F�'nX�Q'N�2�+j��;¸��V����
v�ɱA��.;��\�^q��������ڧ# ��K{*:��Pt��7�R	����e%1����ܡ΂����[7��/�n�g�(7������fA���x��ϐ��2����J��g���iB�r��ҕpv�~���O�3׾�73���g��M�*���x�;���e�<�c��%2���%��� ��^}c����P�,�Z���}`�p#��v���)�Fr+U�3�&�s6c�&�������(�C�����AŴ~����C~T~�-MM���Y���%g���{�:; D�Ҕ����3-�܍�̢�~멟�?GkC\���?u&���Y:��}�Ezf�p�_L�w�e�]�P<�׵�Ό�ua�v�Ѓg6�S��t�R��8�=|#h j���c]T�M���}4�hs���lu�][J=��꿚���j��+�ź:���n?�=�N��~bw;!�!g��w�#�l��Ը����Bs�+�A�S5|<���O���%r�UU��4c���Bkz7�8�fU�=(B@=�A�Mj�^�#�R������(]%�}�e�9yK�P�v���u��nv���3R���R��Q'����}fxR���\R��t�DDB���z��oDý���m���V���H���I��,�h.l:v"�.vˑh顗%���oM]\u�g_i3pK��N��<��.��p��y��E%��=2X��j{�o��,>#kH��輶����aeZ�ˏ�ެ��T�D��y�n��� �k�}_}S��2=���,q�[�M�������^��9�&6~S�K�<��M|��+�l��W�1\g��<�$������lVP��,S�J($Qnv	^c$uc����f��7."�pڰ�%y�v�_C�6T98
��`߁]т����sځN�ӻ�#��5��U�]�P=�WU{y�p%NN�8�0�f��R���p�0�{vK�#��d:�mfE��f�|�g��my��xNg`�˫S��7�擊[&L:��p����V�"Ϯ�c]뛘LL���_�-��
w�R?%����Ά��q{4��y?�0����6�jՃU�z�Ao%?};����a}���c�nz��}�z������{���u�[���M�3�`o�d��Đ�n~�MV�D�^�����֊��[6��.��1�KzL��V��[5ϲv}�瓊��/L`���Ց�����J#�Wc��<��Gg�r�p?\�{�T�ø>��
��d{z$����e9�6'jv��~u�7���9:�)f��Nk�{Ne�Yqs��4��zaK�w��Vq�7k�4�[��B�w�i}ӯ�O$J�(��)PW��N�J�v��:8�*��9Њ�s?tͨ�	؎q��.rh��f����󮗠�v䥠lwҰb�B��\�N\������(��t�PôJ�,�_!3 �wܣ��o�3��n�U�c��n���9od�������q�g�9-��UZ�����4���q�w�\r���{�f���ێ4���9"`ʶ'�/\/*��Gg:��zxj&k���_[����Rp��~ϢOI�o�Osʗ[���ݝMBɈ�;�d����:y�����R��3�g���!p���P��Gn�f����$�Y_\����h���'�Sے�u��F��-�P�ˮ��IJϢ8��k���w���K��;�?Hz�)C��񛕵�a��%"�NC���2K�΃$��+�/[h����N���a
�B\�����@ћ�K�ؽ�'Fdʵ�[m�o�}%��y�z�o��q5�zM[��P�f��j����^~ <f�'���'Ζ��z`df:zo���Cd��9�r~�{_ {me��m�dST|3%�J�s£�C�J[��t�=�����C�����T�?q�>��3�X뉾��ؽjQ��;ʦ�/�z)_��lW?��&�������5��"���ܝ���""����n�k�6�y_�oIݼ��qw<n����{2/���ˮ`_��W������&����j��\�!k�E4�p;�֨�����o��nPn���hZ�R.�B�Âci�֮�ln��=�2�N�d�u]Xu�T�Ǣ{�X0���v�Wǖ��nʳ��vN���y{�`x�V��j��]��/y�p���F�[���YN�N�{[Ք��t��!��мks޸y�&�F�[xiU߄�7�hs�4��.����z#㹇"}��84�QQd)��{z��m�"gVt��B|������Ň��f����{tz��0�Ǯ�վf�Jm��Uj7����9�W1����pU��Iz:�7�k���UL���s%�����'��*x������E�"����	k�!�Ey� ߐ]]�o@E�� ��gv�J���zo8�-��LXYF3��r��m������K�3�:�%u\�a���]n���|�:��W�ϳ=���j�,��~Q\j,5��L�꜃��7���?I�Q�r4�Q�Wv��ؿ%뉚;n�þT��u�;4�L3�z���f�360���4�Jߡ���d��Wx̜y+,�5�US�f��z�S�GuuL����O�lgLŦ'��Yu�G�n�5��zmk}��b�V�Xƕ�{���g���oٝ��ϱΣ���=�4r�8�ت�F�����1�y]ֲڃ���^yE⬘-t�Os�k־P	?{����{8-W���1"wo�f]��� ;��MdOlF�OK'
'(SDm󚌹v��*�NV�,Ǧ�"�Y�4e�-b�׵�[�k�}%���m���+��I ��S��f_jep��[���(�5�^���;�_,6u��D������w\��]lf���@H�^�<�o���y^[�ʼ�d9R�#7_
��L�\��᷂�Tv9^���#9N�ҭ�a6��#�s��'�'{��r@W�ʬ�릶��w�=�;�9�/m�>���^����IED����.��9�j��n��^�2K�s��w���1i�YPm x��yh�c��u�-^ޙĒ�:���d�7��e��s�i���8�OO�����Ϗ}m�+��V���.�J�����ӻ˗}l�
53r�cߧ��lH3�+�e3�m�tfyA�����O�[k��ւ�_���f}Jܛ��������dϪ�-�X�Ƚ�*��<wn�8�|���%�O�o�d�O�[c��ٗ����Aj��Ē�6��Ζ�U���v}L����-o����W:ڻp0�DBf" ���za��R5�x"�f�C wf.{5\���Y���Ɯ�|�:�l�l4�<a:#U}�S�����6�����ށQ�k�r|7���?3Uç��<�eƧ�R�oU:"G��ts�QĘ�]��A�կō�y���m�:���md~!h�4����.�+z|�L:3[�Qܹߗ�u	�o���{U�3���k.t��M��-��y�B�!s��0^Wb��7X�ѭK�+�`h�aVh��6�����z�>ph�G\܏x^�����T�0ܬwR���/�[OUX�]��e��֮0$��#m���ͧyɌu���]��u�]շ�k�xk�w@Vεo{w��6�|{����AcϠ�~+�{�î�v)�c؊Sï���1�8W|:f����yߖ�c-��{��J���b<�=8U��#G@��qy̮3~S�%�������u˟G_]'��9�g�x��Z�����QU�k#{X�Y�ƻ�=�Ƕw��]��Z�ۏ9��}퇪i�Y�l$��}F��^^�OS����TO���P��sq:K��/�!}s�x���O�W
�����k>�>�Wl��L�^��ʙ�\�N�Kٻт�wm��"}N�!�S��k��ں_J��;0.��z�����9�C`=����&�u>9Q�����k�k{����>��[W��� T'"k=�}u�u�|S���iO���t6o�b4'�v��l�H��޺��ϻv�K�6e*��d�.�����~�w�|	~�ӑ�93ق�-<�㽓3��ji�A_Ɔ���u[={f������"���U�}�	�x��i�-i\�j�2Mˠ�-��_%�j։��5��>��sʌ�#���l���{twU�g!ٚ/�E�_y����g�}{M�u㗌��$wc��ʹ"�4z����O�7j�A�v#�׭T�(��<�焌�͘�%J�M=8��YS���U���PjY�f��$���,��)͠���O7�a����i���9�b7L:����I *�B2������:Ox�F���c+	)���uƯVJ.����6�����r k'r���ҷd9�܌�$��j��G��L�ў�f[�P��+��Q�o]ײ6A��]h^���[ћ�U��~��]T����.���ꋴ�a�S��z���.�ٙN<Fp�}/�ƺ�L���O�w�ݽ��eC�|p�_ղA�C�~��T'ܟ�P�S�ދ�>�q��of�e��>���]��/�yg�U���q�����ZZ�Ҧ"`V��v��j��9}w�8�s3�y��B�j��Z��k���pϨϏ�{�d�����5�`9/�t����#h0�K� �5���T���ϼEQuu�y��b�]�@k�o�l�m^��E߳ֱ�2v���9���7|��w��r���ss_���33�����{�� d��0�)��^��fKZ���t�w�T6OT@��+Uc�I}
�yxawp�/bu����P�%�5s���u�\?.���}Q-TΪ�/�͈�� {r}�e�f��JtE�ʕ_�	���eb3ZNN���iE��U���{:V3&���&��
�M^F�W������ȼ���E(��x���o�s:#3��ܢ9���˓b�o�gp��ϥP%���z�Y�Z�i�D����z-�(pf�v:�=�h�1(`t�1�� .����[�8:�ƃ��l^.�U��i�Z��6��g.|�.���b���he��Tt�X4��3y���"��]n�$�Zm�+��>[`���]A��܊W�	��P�5u`�*�y*W���v�����Yv�6��M�:�5��p��i�]���/w7{�2�J�0R�����}x �N`F�uy@�՞t!�UV��Gx�M/)�'�O�#=.�:��S�R�Ux��]�dĔg{�pF8��v���׵��8���<�p\���J�F�U�R��!�&�i��sS�w�fx�^��C��P��`��ś�˗|#��3�U2���`)���#_z�}�=F��ꙒNC�}S�t��~���u5�l>>�Ub�Y��h��z���"gB۝׽r�z͜;,d�"/:�dG���,�ސ'c�s���&{Oa�5:4�Ɵg|.���5�t֙��O��@�ZVl����]Nu��Kv��|���>>���Y%,lo���,�]_���ѳ�#���Y��o����r��/�%��s�$f����UU&�ڦ�c��w�3�|4�۸��Iaף}70;v����(3��tqj캕r��n:a��3����]m<^�!^§�������K_c>�z�t�M:ίv���z3p+fc��D�u�	���}�=�^>��~�-�W�����ْ��uͮ��m-�ɗ�5Q�̛Z6'�/M�mr��X���\��kj���p�˕tq����!.�y��f4��8��sVӔ��}��ܹ%��j�Bm�{P���b��p�Ϣ��s�,1��J���e�/s:p.����9������eﮮ�GͯW�0>k�ZÒo ��u���t3����{�F^L	�"u�8�����@l^�%SZ�+�Tkc�L� :xmuZ�������B"v���W誎����G.(}�'þn%�ZZ��u/}G���"���� m1wK��rza���1�f��YڞuÅ�=�k#�/vڡ+b�fOmv����1�4��鑏��q|�@U��E:��N���=Yr�9�=��?�P�ș�8Ӭ��Rڕ���RoV����z�#u��/���"A�Z�}h��Å�s���]���)��!�(�·�\e.K�kV�vvE�<���Ygn���7�u��f��� �]W?TU�'_�߅���V�����{���v�*��!���M���i�]]�tt�y^w�f}"��DU�$��;�-���;~��1�>�ɫs2����L�����(R��;��s;Ld�8'e�^��q\	���,��u/�75��w�&���E���(:��'>�{�_���6�Qq_���Rf-��~�^t��"�K����d{�E��	��ށ�T)��9y��j���޺����}6��؁�~�R�\��4_�:�����<����R�ޫt�w����}
���,�8+{T������q7�?~A0(��z���`��%Ж��2��;��ʵ3��t����ؖ�E0t����F�4;�;��J��7x�4!���n��*<g3p�9µ,��ݜ6-���֗�(�[��4
祖���כ|_� �V�r|_�X-�7�R�����"!���F�SM]�����O�d�s��>�l]x�RX��cꊂ��M���2H"����Y�D�>�ܠ3{�cق��M�귾�qN����~Ͼ�.�_��������>���p��=��s�︒���{u@��};1+��fvԋ��Ņ城��w~]V֫�P�j37zct����x,�h�]��va���|;��Φe�K�Ae`�geʫ�W�Vo�s�>�g�];9�ذ%Ps;�=�2=�:`����z����[����J}�3�O���,�7ѫ����Æ��=��K�'f��%���h�~�g�?�OU���gẄ��(tg����{Uq�/����FK�3�����d�J}�鹽z�w��׵.�cqwJ�Z,9L��&|{��8(}��B�W�<\n]��b���y;�䙵�,JS|>��Ѣ�>��<���y�7&��ϲ��/�mE>uu�Tk�&�P��_S�'���'���fĥK&U�	{�ō=��
��7�]_��1�L�>�](zq����6�Sɂ{�7F/�q���ԅCٗ`-�v�jE��f�vH�n��mggT@A�W�a>٠�!wL*���������_�*�6�Ş��s�ܤ�j�Y��qW��F^<3ps���Ua��4;�d��9���*c�l��4�?���D��q�5���ᣇF��*N6�;��7+.1z*;w�J糱��K�
��Gwm�X��й1��ڔI71u�L:��8�ט��rd}��\�g���y�gn��w�M�ވt�U����g���uZis�C�=S�2��&��]gh�۝Muu sR��Z�j�:�gf��QA��}[�z�z����7^[e����:��e$������_Q�n�ȸ���x���X��� Q"�iZ�es��SmwS��f�ۧ�����O?�茢��U� ;IC������W��x��v�s���J;��`N�r��;4&ڧTʳ�����mM�!E#k���β��!d�z�W,����2im�XH��4�nf�r�o9�/���9�\+��[]��ݙ��u�"ku�I�y���)���CᄓD�wA���FL�7Tq����{]
(��_Ph$R��W72�GV�U�],͂:�j
|�,/3��^cՒЕ�)f4z-�y*��c������(�m�yFF��MO�P����I�9L������6+��4�5-�θ�q��Nٖ[���c+��7��Ǔ{��8aLT�J�`gl%�(��Z�o��\-�"�VhQ"?�k��3�*�i�w�X�Wʬ;�����:໾G���*��11+Fiئ�����"���t�2]v��_Fz�_B�v�IO�Kd�E�2n�����|3��侹c�;-�k�/o ��:��l���x�i,@��8Vq��b\6��������5p]�nj�f�F.�nra��ބ
H-�w3���[��},����;\���"5oJ,Ր��*�J9�,�8�����A�೿[���s�SDb��m�'���;���L���{Ym1�.*-!�K�����A��@!*��ׇr��X挭�]'_.��D^0=OZv荷��;�˳ �!T�����@p����g)/���X5��7o����!��8���|�xHf๧�4��Z���K4���h�7'��0���ARf�
��@;�ջ.���m;έ�U�#9ؾ���dwIV��:�
�R��0�U����v��]��4Y<9�;'p^��,���u��u�+F�e��lެ�qXv7]ږ�.�o;�rm���LmD���L�\;��R�x�����=�㬈va��&c;���7�]�ݝ�(�"Q���/�u�NG27F����H;�G!��:�P`�j�+L�1�+��33=u�U:G���Q0���״s�e���u�ḽ��F�f:�mf3U�Qp�G�7N�[y��:����ƣ�ծ;���N.k�g7��*�n��+�F�kaM��ɣAٝ�L�1+���&�a��@9o
Z� :��~�n�;ka���aO*ʉ�=�G4tffR8N"�t�6��9�Q�`�R#�o8)��.�ou֞�o��9Xx�����eb�r¥ܶ�e~�8Q=jM�_噷f��Μ3�Ec>H��$��X�k�`R�X�ʗY�|L�n\mL�X�z��}zr�g֝O`�o���>U�%�%���Hz���y=1������}��q�!��g�}�C�߮ߗF������L�q�Gt��'�s�`�����SVs2��]d�x���w:��o��jX���8'�w�{{�5h�ܷ��q��SS�=�u�2<D�L�"�#�Xݮ�^b%{��8��0�՘�̶q��'&�F�K�/��^_|c�n|&����,݈�:�|O��bUu`J�u~T�_x�����Å����1�fe~���?�xg��z����<n*����2v}�ܬ�m֌���z':��E�d(=�4�py[~SU ��ys�>�n3�xe�m"j�%�sԞ��>���|�{�
�ꝕ��r���s|O�:��B���d�S<-f�5�l�u��������Շu�k+����K���F'ރY��Yf275�/'gx#φi��\��1O"]�z;�U��_TK��u/��֑�+l��ʺg���f�ni>�0���;G:j'�~]Qw�^���@�U�{:��\����_����̼q ����w�?q�B�7��/T�m�������6�oQ�ݲ����k��c����hF ����܋�Ҷ������t���wc9����%J<�+��`�9���dk��e�+���\�C���K��+x�w�X ݝ�k9(��K~����;�}?s����=�Y��&��g�Ep�T;��}���,��{�9�ʦ>;��螭��_�i�]EX���}>3�����t�]9骥�vxf��n��uvǻ;:�1|c�TK��5�`�?h�^�Dr�d�)���]z�qe���XT��ͅ��WX�|�c�zG�U�˾���є�+fA��4����n��rd��ʗI����=Ж�����u��^.=�ܤ�vo���ۑ
難S�ɱ�<\�hҹ�/�u<�=''�G?'�f2錚��(�m���e�8��'��j��}�C����)24��o\ɜ�vh���hc��w��y��c�w[� ��;�V�^�k��<�*�K|]S����>����q��wŰ?�m+sWú&sb��G��*���>����/�޹�a�zrv,���^|���R�WuL�FUl�[@u<�u^����Ɍ�����7�e��V2�A�=VrC�>�� ��[q�N��a�3�K�~s�����דpfc�d		��#8z6�f]N/7��P�J�_�ý������s.�k��]˅�܍���o��ztR�������E˹X0���P��u����2w.�^;���j2�6Nq܎�����:���]�0`�r�����2T�)ˀ���ވ�w!�@]������h���S���Ï�$����wX�/��ڗ�� �K��o�O7�rf���21�ȏ�����N	YʶV3@��{\nJ�Y�|�6@We3}C�%�N/����[u�I/]d��x}u'���MWvÒ���t�>&~�7q��.z
�Q>ob#�Z0_D�U�uF|�}�
�/����Y���ك�>|��^q�fy��0b�<[;}[@��۹��۟(|}8Oݣ
#�x�K�/�W�7K�89gl]�σuΨz����͇;�� wv�VW�mH�n篽Y�j�X�^ ?\����̽*Q�k<��l��5@��'�(m݇&�W��%c��1�ޘ�A��o�����'E�g�n�hD�*�R��#��u�>u ��[��L�W�}��e�k�]s>�I����1Ǘ�zlgЇ�#ޟT��ۃ*W�	�!QF��������f,����V*viҬ�����B�Ug�?d[�H9�^���sm$�e��~�}�25��A����|�����ul��pr~D���!6c�7(V���]���˛��Y�K�y���ZB�ܿnw�V��2W�ͯ��������`��p��3���7���,o���+}j�aS�Fc��]�{��>�<ua1C��^��T��+�vH�M��*�=,���{*6=i��dZƼ�ݹ,*�'F�ߪS<�h\�!����-��ʏ���@Ia�3^�ۮ)O��iY?=�4�&r���%]�e�����A�{QevV��v�Z����!�C�D��57���;4
Â4�{f�YJ�Э��P�
�f�j�Dwᇺ�M�wU=��(<U�6^�o�g�'u]q�oG{7 \�7��n.̈́�x��
�-����)Ns�Le1�ћ���#��Τb��y�z��G_�vϬ]߃ja����^G\m_��d�K�خ��5�\��_�w^ȕ�Gx�	׳�]��6�t�֘����9��}�n���):g�Ζ�;25PO�������^?b8�y�ؽ�1[�X�WÙ����_F�C��ʨ��Ɨ�|�=p9xN!�\g�<�5�e��P�
,ů�����ѹ|0�vU�&I��z�*��g`(�z#`7�b���k�B�/l{9'X�����J.���1����=�t�g)���0���Iy�`��&iw�T"��|f��<���{�@�^a>?v��ɰoE�E�3��dt��G�6$.�(Gf��m�g����rf�~Kor�����{�5�ɽڎS��{3�g��뉘F�UGEq�U^&��6J�YY̭8��qX������}�RA��0�a[�����:i8��������Չ0 �t��&V��EZ�&�ى�g;������=I��aU='�o���Ş���ķp&~[�ҽ)+�T�ߢ<_���IM=6b�2���{Ϊ�geηS.7v� m�H�\��tL�����W��h]EMo��\2Eu������ɼ���%���F�l�ZmM��S�����;�OH�ߘl��{K�2]��Ԝ2��\��.��/�$p���T�qO�.8���)�����dx����2���T�y�!���>
�u�]�8�z#�2�ѣ1z)�wg�v��='�"T�i��^�֥9���T����`*'�nfbP]n��%��ً���������d䜎��]���H��ϱE�/R�m=4�s��lF��+N�&���c���P�Ǧ���E�"dl���O��]k"3�pX�w���Q���TE�IK���ߡ�/}�gk@BmT*��_���oz�y��O �k�jP�q]-�7�sП�8��?��'m꺥^�������ȩ����!��k�hmeK�O$�^�D>��6ɃE|ٓ�D����z�d��4�K�����p�u�����������}[d�e��������a�T̭���6��n��L~���:|���#����GG9�(�]#���^��-���*; +s&�U��@��:k7�^�Ď�KQ�Ұ�m�q����~5�MQ�N�7d��>c�D��`f�=I�q��gD}`���+*�2|�4��/��m�50���zRz@����^LbY�}i��🳫~��T��\��$c���#�ݥc�ᝎ���Q�\��b�3��)���p�w��9u�+��8��M���L5�h��)7!�2K�J��=����7�ّs���;��O5J�O�Q��!W��j5	5pC���<�Pʺ�o�dsee�۲�r�����f����i9��n볳m�1-��ZUrv4���lA@X�%̕(Ǘ�3���s���ͷ3���Ň<oM�<�|��3��\,��yk��k�U0_��<,�H����j\������y�f$Q�� �X�=������<!��{'��)^�Q݋p����^�-�����;�����]x�Q�ݒ����Q�૮�hLnz��@�,5�����
���7>F��NJ G{É0GDNɼ�Q�ޮ���D����qh�z{�f{�:�D]շ�;c�}*����Y�2^�	�%�a=�އ�LF[��;�== �1;�����r���h�yt��Q|�a��N��F]/u!������uu�ty�1�<GE��uv�gp 
����d��A�����U�3�Yku¬+����b��y��k_)�c9 b�8�*��=^�k���^o}����;�N�]d���r�:�y*mj�3>J���ϸ7ʞ��+���W�τ�@}�şmw��j�v��KU�z#��H/�eB�}��e�R(����2�쵢��`�^�Fm��=��R5>�o�P�3�Mp�y��A93���`{^�l�.A�n9�F�U�Go�޻7�鮚Z{��8���\��J�����F�����"��w�ӳA:����E�*<]����^^��|y;��^t�.3�J�c�w�ȿ���y�U:�t�b�����Wp�-�U������IR���'*1t`�/�K38 1�:�f�^u^+�f�)����O :��9����-���Տ:�ZPv�����S��:�u�,j��m,�x9�V��s��,8���7�-�.Y�ʷ�$�r���h�ޔ=�@ڮ;[&��R���-v=���	?���e����tq-�I�
�?:1E>8�u�Uv_F"N}4{}:n���_j��#����絥��s��yˮ�U��������w��=�$��k�Q~d�A[Y[���{�C��.���ԣ<'��U�_��x��>N'�]���=*��v�lt?%~������~{R>��jʢ
�Ϧ��mWR�N��}��\��3��s�Mm�j7G��bѤ+
FT9��{�G�����w��
d���+�'�GB.���\��xeT��o�dJ��O�=#d��Y;���4�m#,{�]����?33�]UM��=]�ݬ�/��j�O�u�s�Á�wdW�I�P=[��;j�G�όV�V}���Wd�Eu��Mu�����̋�p��9�,\>��Pn�IeW�J�"m���GK��:�Mg�JD�ùZl V�]C1/4I��uப��D/=�	�d@�zor�܌<v����"�$/]P���7v2�{y3᳗��`٤.8��.�޲&"3!4�;.ȞV�㗗�LoTl�y����`l�P���mü��rU������\�t���q�g�yr�%�N�EA�+� _g{�%QX+�Tt_]�Z�;����^��#<ƣ{����2��*��R�:���E�n`C���w�r�5YSgq/)a] �)��(�;F�i�ʒ����2�^#i7���So0'hM�3�{A���n�X!M�L��x��y�l���L���4�*��K���%�Z.�a����	E�]������Ŏ��3�R�VϘx�^;E+���n���-a�_���ͮ5Y��e��><�Tj���Nj#5jݮ��dm$nDWm�;Iw��>=R�O�! ����0y�ZC�Z9{+>���9<5��)�\-�/����em����������r����E}����ץDE[���$�0(����5a�\bC�;?C���e�R�g!U	-����rzla�M��UwEnq�u�Ew{��in'K�V �7� ��٤Q:��7�]�.��q��g�X�؝5�Ӻ	�e�*]�=�:ӝ�J��5�͖�������|P�)J�����Y��p�7�ؽ�j����]Z>��\��P���uX<G�{��м��O1�Բ����8�������ۻ���j�C�nk'W�)�W�at�s�1~�����u�Z5�f��O�@�2���u���o%��A�iye���ݳC��Ü�S_�� �e�|g�7�6 �B�7�тs��Ը�
�$G��C��/��\���R�5�,���|<//.���$���^�������*���x������*�*��a	�����{��	"S/(����/�,�=R,+>�["��A�],μ��L��;�Ǵu�"�v�ҹ�m+�Y�}ľ���(�f�q�s>�����J�uJ���	漵S>����I录����r�JB�w-]�쩕�x]S�;�z�^u>�ҍ�WD?k=v[��,ֻ(��\4�omc����o7�~(�� �w]�!w�2J�H΅Iz&�aKμ�u��RS(��s)����:^�0�[�{��+�M���Ļ�*� ���g���|�8����Fg���I?Gq�f�;�ʂ�'������e��ׇ���N/�S���<2h�a�7]]*��v�[U��b�b`��q��=^�b�8�bnp�}��u�B�w�'uj�����C(���@����<7��"We\��m	U�W���O�n�R�{�����aԷ@_��f]W�ԑ�W�ψ^�3�g�v]z�EL�����o�t{ ��|�&T���$+��
N�h�����CT�?e��ѫ	C�_X�97:z���uS'½�<���#�U�&z�#C�"����Ey�{%P �ߣ��$�׿�4�����E���R>���]�{{�����k�g�x��.=��ͻ�#�>�`��ç��>��g;d�^v$6��=
g��@֫���#v9G��z�KF0dy7k8<����ό�LDGp>���{��H�B�okqR�A�M���Ĉw�P���wMp5��ܦT߃t'�����K=2n��;�����֠�I1zz�dWq��:�b��y�C�2t���Q�v�MJu��h�/�(�ڿV�b�>@]艙�=�3c3A&��DGBfrW��a��5�=&a�yp#`N���y���.�EU��e�o�h�~��T��9WE�F/�d�����:��^����Y��5"�H������KN�e��E7�-�um��w[:3�f�^�}\��v�E�����*tb�m)<�D3�ܬ���ױ�n�kU��@;�񫵍�U�����U��F��^����P�u�[.}����]�ݽi�`J|�F��_v�2�p��J�4}�<$���ww�o�I��T}�T��s���¯m�ek��4���%9�޷k�0ѕ�9�J�V;(v�y�q����(��ɞ���:�a/U������dl�����T��g'�nu�N

��Qo}�<�[/��'��xψb�>��[�?I�� ��
��@1���ُ3�>�f=��!�3���-S�-�o#���W�'�A�Uu�7��#U�{����[�޹��բ�2�"��5>�j��z�`��\j��{Έ���Ϸ�WI�h�vQV�_��ntS�F6�p;��f_������t���۔p?ޛ��5S���ۻ�6Z���}�f�����-ٺ}`z3�\_��8���u�t@{�o��j�Ύ]��~I�"\*|~3�b��}lp,��莚��.��� �}�i�։3� {UhVj�j7Z��<�o��x�o�q�c�E���c��P�[��ɽ��y�đq.ݪ�1
\^��c����E\���o��;�'�m<:�<�2)�����Y1;�\��rW�_+?M�@�֋�|�*U��@��m��x�hO�uf�
�OuJ����d�a�a;���f~�"@��wA.�|:̻}I��eSx����n*9Эgq��v�4@�q���4m�a��.n��kcU-ͽʽW�x�MM�ѓ�+�j��|D�����n�u[�v�;��I]�ח��B��g�n���i�֮�)pZ�F�D�Н�;3���%��:�+�R��g'.�M��֫��Qs��ա�1q���c472Ԯި�f���/�1E���WM����yxŠ�.Ҝ'i��s�M�6��>���%JniBu��Z�]vV��\�wm��0$�s�9A���0_6y��,=0�Z\�SX3�����ut66CQ�x�����j��CΏJ}��/q^땝�MJ87��%�t����y>%��2�����M<�&
���se��B�`�p����������,�y,���J���(�8V#1��:�뺡�����l˘^
ɟ���)�U ���z-ͬX4��o1���c�q8U똀�3lT��m>t�\�����+��|�iJ�D\���ʓ�9m�������Pq���}�/)#tÙ��Q�f�D��@=�N��M��4���Rx�s������4V[����-��e�so�t?�Y���u�mpY�1��1a���uOv�1^u�`!��p�a�-J젏o(Ƹ�xE��
�ٝewP�k�X���E�u �`w˱ui�J37��%cb��s��C��9fs#n8�{�9Bd�^�&�=���*k�ՍfX�*�԰�j�uv.&�	�J�i2n�N��Ȋ��vJ�Η#�\Yr��6%i��c��w[���%v�����ӻ�wOt��0U,�]�E� _'��j�M��Y��V��Z�Y�C�,�90��VwRX�#p�[���,纷fV�d��̹N��b�j
K�=���͝:��[�Fk�ZV����M���н9Z�PNT�&]fd	�$�����Ӻb��	j�Ik��A�!+��.g
����S-��*՗����=�y҄�F�g�	�fJzd�2����/;f��!��P^�-��f�燨r��U��X���e��S"��]^���ҩ��v.�do[ �\sv�;�86��p����u��ӧB���N�Zv�b�K:wK7AkLM�P�~�r'��Y����u�s��n��0Ԩz�e�g^�E�u�8��J�C�#��[{� �ڇM��9t.X�\gGN����	��.��|�>�F�g-d����;�뮁�B��ξg���������S2r�����Nfd�E�K8ř?3��ܡr��(��,���-'7p���E%-�Ǫ��#r>��w+��3ijVgI��*�J���H���a�Ni�Θ��*����w%��n݂OP�'�(1KJ�wⷮ@	�7��瘐���8��k�����t��Tfӫ�?�H���@���NEd�lN��U�:�{�qy%��I;�zTO�;Q�xmn�Tmjv�����%s-'��Q��r�ͪ�����ܥ�eZ��B�{.��W8�:q��z��K��Έ��n���ۦ��.Ҹ��W�ԏ��ެ�`�0ӧ2�e1ӣ�T��T�V���Noay�{�'�����3���ր����V��X���Gκ�L{��09���9�Y|�_Ou��=��g�ޑ�����v9S�Y�A�8���H�:�81_0�g�C�_�J̏�8�sP(ݟ-/���.E!7���y����f$2b}k;RT�	[�D���pw�~@V�;�>�Ӳ��N��J�������/~ݺtۯ��)�[��o�.��|�)밫7z׺MZ���}5�?g}�1\��n��u��L���C����,���mDX-�F�X�yo��آ���\yM���ퟞ��'�����f/oUQ>�"]�&,����X��-���n��Z{?U���R.�K�^�}�Qwe� ܼPU�=C)Rn�>_.���>�:�S�}���}�x2M���W�B�&e7���$]���+��r�Y"��9�yDF�^�v��Q9+�U�eY�q�թ�2W;����J���;�(��=ku�=V�>�ܶ]�'���5�QHF���TA�nK��؝;�9u��mD�x����'�J�_�>Y��Tx�ez2�:�b�*k;�_ԭU��^��:�,�0ee��t��f^D�>ΐ.�z�9\3�r=p�G��F��̮.|U�z���5kOx#}�����2s��n ��=��-�x&�{�X���ן�ӄ�����u�gO���[)K��z]fBi���/����0��-w�m�,g�??��J[y 괨x-��<��� +��KyN�t�kZ9.�"��p�]���YN���p�e�u=��ԉ-����7}��E�5�S��uv����:���늛�Д����:�wy|�Ò�X~����}t1��E)�O_#Lǻ����q"4�Q{Kjb��ˆMU�ꅟM����**^֨�>����_{��yg�wb�$��u}��!���N�fo�B7˦�d��:��	���U@��e���n��Z�A�FQ�(e{��<q��ft��{+)���C���(��H�h��joy�	��F���Z^��#�	�H8�}��r�>�l̼G�s&�	}��{˧��o�{o �Ay�����ާ6���it���CG�
��|q��jS��L8�I
��O(���ӗ��!^��.y�T����b�:Tg/�LwG�qw�g�Y}���
���ՍM签>�����W��)�����t؏wG��L��<�꼌�R$�JZq�_�ur��9#)��l"�������ը���5�zo����\[����񁑑�jz\�")�0Mχ���6=KӞ��"+�z֫��@��{��\�U;cl������Y�x�^��>�{��3�܁R��\D1�u��U�Q�w��A]ұ{_�6�<O�Y��6���\�@�́�k�®��]��^f�D���N�ޝ������u��*n<�tϪ���J�-۳�>Һq�ݻ�w��<��z\�.�3&*i�6���q�`9�μ�<��'���{n{J��S~��sZ�<!-�禕W�]x<\G�\�
���ضHh^�]��dft٦X�l�c�d�\i���c��37���W:����T�hg^ 7N��Q9�������of�Cs�x�l@���b�r]�=Il����27�wucSK�"DiZB�z��b�˛�ӻ	NF,;��z�k������h��!�>���ʺ�ՙ�~dW��n	ٚf�B��σt��H_�O/��WF��E��&ɫ̓�[b�f>"�cȣd7s]��7�n����\[�?�}��\�[���԰_����!W���9=����$�l��>2
�w��Z�*r���Ƛ��O��9�J���{ d�C�u��f�Z����<������7;��Ӿ����n*bf}Q��n��$Ȝ�� U�UE�99�K��@a4���g����v���2j��L^��2�^�'ᬕ?@���/�7�����,k�n`k��|���K�y����L̞��(6}Y��hCQ��?�J�����5���{<�-z�&�vGh���<�c�Y�����r|2�۴���%A��9�]/U�mʏkRA����ԡ��e��>5_.f��=��uM��uz�-lwxr���L������>�n닏��&j�~����Sx�d%�ʸ�?H�Xk���l��כt�s�[���'_N�؞������.ν�N���]P�St���<�"��G���dø���c�W.��¾G!�	�]�c�'��N��%U|���]���'ʽ�}��%��`�N�[
_�ۥ~�k�W��Z��fφ���ǧ�ە��ȅ{:��Td��,"� e9�5�^M���M��b����.϶�p�z�P���:��rL��x?��m� s� \,^�1��כ����9]�쏩d��.~��+�X[�k��Z\Wei���cóVu�Sqoi��eV�h�>������[G2�_c��[����~�U��']&4�q��%>����5%�1�|�,���k8��y��}Y�emv��z������k����7�ӕg��#}h}�I�\�~i����V�x7�}�<�B�m����\E�ܽ��	�ϡz���U�	8vu�nnNg�a�^S[!o�6~)�9���F;�xPdk���7@o���E�U�-�T`��﫡g���|��x��Z�6�7ل��r���z�tQ7]3=o�ړl$r�a��OT����u�G;�M���G�*� �&�����<�咽�?G̮��jB�c���Ö��ޥv�U��&�����7����m`��33���>mϏ�wNW��u튌-���/ޟo��xSܦ.�Ǟ�̘q}§�<7�Î��j��-�S���}b�e �G2��Ʋ�}�n�SG� ���옹��ގb#x�s}�E��$*����n_�@O�V/��~V�,���~Y�2��bqSX��T+���g�v�6����/�q�ˈU�Y�,�2��0"~<��PΎ_{v}�5��m��!]��Tn�3��
�*?^9�6i~�yV�lݏ���ga� ��_�-��?�����ߒn��w���#�O��џS����W{H�IڏN�of'r���og}~VE����Sݩ�����Ҍ�T����-܂G\��ܒ��Q���.���uv�ɻ��:���ؔ*P�P���;�E�~�stX�>�����#&eS������ g�+��~\����n���>��~�uRFj�B/���yobڳ[�I��*���{)�{�U�*U�0+�4b"���L�Z5����1�Yڮ���e��JL%�rV�*��5�p�-�
�Z�)V���oޣ��ʴ�ڥ����(�Zj��Q��xn�r�o��lFy,��yi�(��R�s�_��m��T3������)���=+�Q{�x��"l}� �R�f�_���ȗO++�+~���G�H�y4�I��)Nf��#g�7t=a�!���ٌ?:cU����_��]S�l�W���7Ԉ�8�䦢[�i��2O#/n=q��\�x�Y�#�{�w5X�Đo�}�וV`ǩ
��{yc��vvo������~Qe_�~���ߒ�r|���Q�Clԯ{�W�x3:v�duI�n̞.����\ω��S��$��q#~+����y陽���u��/罓�'���^6�H=�1�W�ۛʧ}�y��h�N�q]h4�8�Hy����y{@�}p�\~n>��;�ۢʹ�ڱ��͝~u�P���,K�ƠE;�3&�w#�c��J� ��Ǧ����g����vB�������z�����l�,Ww��	���'����X�/���"�7���^��{�r�}�SO!�1�(Y��<�(���gDWԟ^���l�}F}��8��'mk;�0	��|~#�|lNa�-�ꞩ<f(�����r`�m_���
>"�]�B����|`_�s����
>��E��Yr��GG�{ ��I�E�E��g{ě�5��Kã�/���`^����u����sUl�X��N����b�ܮ���#O����R������*(�*�i��>�E�s�v������w�H4ǫ��ug�pҘȡU�Vs"iO��S^s۾ȷ^��~߽��_�{��"j��{�/X�=���*\pÆ����+s�<ğ{�J�ic�Am�Ee2�5�$X)ѶJ��A�0�|E݇�!m@o�6Wyz+��h�{|�fK}�ys�#���Vt��P���W��E�e�o��jeu��ۊֲ����#]pB�$&�r��y�=+���m+�����z��b����w0=����^I����|����e���%j�DQ��6 ��k�y��?�Y��Fy/$�wg��)?M�������ҫE��ԅ@Ϋ�����i�;5��3m��C�U��:��j
�b��[ǯ�׵�9}T�v����s���"�C�C�E��~{q���W=�3'e��!�����)�O�V����>��u}ǰ��L����P� �f}�;w�]f����}'����}c��So�>#`�k���w�4R�Q��ǈ�?\��# ڕ!f�E�yM��9���1?���$��VM��D��ݮ����Ω����g�uUT�U;�Y�~�mxyܱ+0}jO������[g}�մף"�~�^�c�Emt3e�/�5E|/$Ͼ�������]�fZi(n��'����W��9�/�����W*)!P2���6>�ȋ�;���64���a7]��ռ~(P>�����-g��[c;��Ǎ�99��W�eI����^�� �Ǻ}��b�Q���[�>����D}n�z�o���D�8[��h^q"NOg\�t���~�؇ٳ_ Q���x�d���9���ۭ!��[䌓)�CiN�A6��+�׿.���J��%�x:�Y�9�7�}S�i�;}BN�t���|kt{l��'H���OO���bL9lc��� �#}5�P��t���h#�� ���HP�=���#�#��h�g���U�m)���ƻ���P��SR '�zx��O�\�I�b����}�T[������.HGK*�d#�{�(k�pR�b[�rF9�ٌ��&��"X����o7a�}�����-�Pʷ�m�۷r���ۜ�2VشbMWV��uXF�U;w��bn�hcd[��=+��&˔!VV��W0���.�B�=��������X����sj�ڀ�/���{�Q���L�E��:�3��V}���
����k�zP��4�ۉ#�ｱ��֊h{ꆼ�jG���@�y�����$
#���!8}k���V׉��@�«p�� :!1��F{� ���M+�?L�]_�{�7ī�ު�����UH!_�����-r�b�׾�}uE�Vg�!ݺ��|�5�yM��a|�Dr�D{�dy�xFc��������<C���bJ�S�:�����;������Չ>��� :2�.��ɳ��Ir�a�
ת�	7�.�'pQz����D�˙!ۘ�o�灂6[1������"LyȏGvf��9��5��⻇<�t���a�0�Y"]�W=�?}wt��}�?}�͒���`�&���H�敏I
���\{��	1)��؝�у�H��BA:���>��onWAٻ���B.�Rs��ߥ�!������"���,��S���[���}��~�D��H��ǮyLr�廉�Ҭ�%�)]���@�������\�nK�j��4j2U���2>#�S�W��;���f�(��g��Ő�.�]��~��+~�}����G_٤
��	d������:G�S<rG9ZJ�M}�Ɲ}Q�vs0�9�@?*rd�A=C�+Ng-�A�_W͖�xMT�#��ܥ6-t��-�c��� ���Ɨ�O�x�%����E������f�K+ݜ~�o�^Oq�g��	I\��Ab��*jI�8vd?b��1�)����]S�O鋋��`���7�^�*yo�+pN�$GC�u��wUݽ��g}� �@��gW��ij��f/�!g�^ڵ�"���YQ���ӳfHd�mGާ�_*���H
Dm���hgF�Ϥu�^�"�|��Sѷ	�/隩lv5�t�n��W����H��E�x�n�f��Z+rf���V�IQ����ͭ���*�3�q�����8v�i�-��T�D��7i�H+{wi� SL��m^Y�gzh��슶�X��>�M��e>�n��$�z�}Rt��W���[K��� O�e����T�<z3 9�zUQ����=b��	1�Q���)6�z֑�/�e�����7�G��U_o�V�sK҆�=�j$?\�F�O�sd|W79����񏞀(�k�)d�����eX��P�����Ta���eM����5?]�S���<�����S��C�E�}9S��C �nP���-!�
�x�:P�hQEr�"��5vTz��c�_L>��q���J�S�}���|J5�@w*�@o3����q�uo<���qdǼ&DB�������I���	�1�U�{z�t����da�=��F��9�a�]�h��"�޹�J���3�r����aӨMB.ay����l�Pg�"}�tNy;������pe���H��3�ە�Ϋ_w��*�c5	a\+���F���+)_`5��%�E��~}�[b�0��O�����,�3�yИ��#O��_w��B"��� �a �5�)�|��R�����s[S��+�><Y�����C=�߷C&`#ՓfMm�Sʚ����y�X��đeI�w�1�ZF����}0�J�s�*F�������G��=�D�W޾UA�DT}��:TlK�"��/��bQ��x�@s������#�T��U�~k�M�����@�S��X�R����2Ti��K�cf�x��9��z�>�9�������a�>���5󦇺� �E��H��h#f�1~QDO�l��9&0�h���̐9��K�}7�����`���Pu"O�3jcԕG�ok�;$}z^b��>(Ƒ�MT�B0� }�{3�Fϗ��Y�ԏP[I�w�ڳd7�v��\>_zR�w0��#ˆ�s���ж|�~J�����iR���ɹB]�hh1�HӗR�Q3{���h�soL�FtɈP���[y���<|���r'��o=�b<�:R��+��EW_�h������2��|�\����榗�}���ם�Dl�@�֝��~0�\c�|lD��'�� �TC*8�%j�M,������F�`�P�!�d��4�~5��#����7Ǟ�w_}#�ϕ���ig^I��n��Q$#g�L͸��c��Y���E��cƹ+@�����fϨ~4�㟖h"&2����uD�вD1�D�Z�{36�;�/�O�i��w<ZC"��(@��a�`�}�'����TrL�/ �$|Q��}�Y�P>��u��)�����Z���<��]��{��'+��1�m�P��ҥ޷��~8c�q���،Ԥ��W��g�����ag�VG��y������Ydqz�2Ǫ��� ��ʛ��>��Ř޵��|��)�"�՝c�2�o�Q�F�������">,�7\a�^�V�%�`��_(���v���#>����:LyQ���pbn�O�����⭻�2䁲�#	�,1~hg}.�V�� �:�z�aF�\G�b���$0���}a�2��62�=�T x뿻\^?�Dg��@TY��w뿕�ڛ�?�Ɠ�B�yC!�UßH�%H�r�c��"S���P�Q�7*��Y��ɎH k쏭X�Q�� {�%��1���l{�O�H�N�����[��߫S�>����9�S�P>P��|��dA�Đ�Ki�8P|@)EGO���q��$�f>0��:��ʀ��� Y]Q�FVD��w[u�������V����R�7�B��Ƈ<I!�����0Ȁ�D_�o�3>bZ�������Id�Tk�~~�B"Y m}���N@K�[��1˃��M�U���P���/ݛ-�U(���x���)^�0����T$�? �Z�$�#�6	�� �R��Up<�U@���$�0̟1'�&�@���b�ɛ#� ��+.#Ő(��S��.�x~���?)��la���vn<�Uo��Ŏ�m	�&b4�۰ҳJV��O�i�Ib�o�IAuA�Q�p=�tJ�'��ծ����;�(E�V'ww�Z�%ݒf��y���Z�:YlE��e'�9��vr�pi���\���]j��{��@+wd!�Uቸ������KWw��#�1�O7@x�� |c�J4,��SR�j:�p�Edy������ﱁ�Ͱ�>b�'"A�|�I]!(zQ�b�${��C6H������w]��=�x��b��]@�"��#]F��������� ��\}ޚ0�DF{!�[t�!S�W� ��F�|@��+�#�(�}�4Ƒ�ʼd�h
"L@�-��H��
������/�O_p���f�ΰA��k ,C�|��P�(c��>6Di��grE|��=(��� |�`q��G���	�C�@}JH��ȸ>R�I�cZ��AD�c�r��c]z�	�s]ٕ<�S����#�FJ�0	u_�vG���cm>1�b�t�+�B"�R@I�bI �TF�!��jS	fۏ��q��)��Ү�c�P����e�����]z�ծ��7�|� "8�p��lDY�`F�0>1P�d"ԁ�w�"��L3? ���#�@i���
��DV���Ta�?0=hG��� xW��9 A��!�$���J��x�X�W�����Zf�{{�9���|�4�	 4��b�
 a�F�חQS#�P@��!�	�A"*�G���x����"}L�A ��S�� kB*���` QG7b�b=j3J֠d� $�r5ʘ��u�����Яv����Q��'�DGZ��g}Q؀@�B1��E� }�d|D~"UȈDa��C q��1���Q�"���H� ih��Q��!����4�2T@� JP,�nnz~o�Op&Y�=6]��
z�w�������bʏ�&0��I�D|b1�����0!�O��>1�	"%D���0RȈ�1��`a؀��q@��P $��"L��3���I���9?/���c�w��D
1��I@f ����d��D���D���gH��@`2�DC1k�""�B �i�� G�$��|���b��1h $��Q�>�� f����>��hdq��>�7C������b>� Gr�O�P�0��� `#;T 4Ɂ�?*��DBJ�Lя#҅�r��F��~^������@ ��P  DD�� "#�� �� @���� @���` @���� ""?� ""?�  D���� "#�� @���D @���  �
  D��  DD  DDB  DD   �"�  "DG�  "DG�  "DF� ���(+$�k%]��@ �K�
 ����������>w��l
q�lo��H����*�!"���=�i�L�  ��@ EO`�TR��р L&�` ����!J�2 ��	�M�	Mi���h�    %"��O&��x�� �����'���?J6S��!�����tAJ㚊�DEL�;���++����X�($I	"؁Q*��P���
���G_�m3�T��ˑQ"t5��a����x�&�IM��)�N鍷4�)h�&֤��{��W7�nj2��+%2T�jŨ��Z�T=Ʀ�m����ͥ����K� �!�D��:C	�߀�gD��+�qu{��݂L�	0`	�$�I��& �L�	0�`$�I�� L&L�	0�`$�I�� L&L�`	0`$�8K���r�i�i̖�wJA\<�N#'E�8�s4��N9��p�Y�����ظ6WZ�} "���:

<P��ȹ�*��Q$�d��cHZU" ^XWto7��$�&	$�r%^���Ǐ^=�r������j���}�߂��ڈ^�������I�7b�,c��j�:􋛼qr�DpA!Fsy�if�k���S躃L�3�1�ST!�bZ�����ֽ:���K�`�L��Ot/��^}�Y�O8K�湫�LS�yu�m$�1i��C0�L0;5˶#t��-K��Wh�S.����MI���.�R��0�v��1֜iۆ���X��/W/I��ݻJ:GI�e�X��!ڑ�m6+DS�?!��v�SO/zUH-qA�p�^|�wɘ�,���� I&	�ɡ����BI1��;�4�&�A)�z��*``I�*C:I�N�hJb��(�I�	1A� ��2Uc��%D���D$%�8�	�	�&J�! �D$@�tq����^TUiB
M�9V�W���̑6�r�孠�sR7����KqZ2%�5#���5,C�'/rRt�L:���Wiܵ����D�Ci"T��nLS�N�A��*��6��t�~���dS��].�I0��fP�yC��pA>�yJ�3�:�:�/y���Rr7iiZ��멙@Tݐ�[1Q7f�1�K J�G���Ӿ]��=靃��a�x�A�K�:��1�'ʰ�y��y������d�\a�4�	�I0�3q��B��;�=��v�w�҈�VvUO9�F;��7�qO��Ӂ͵:�l�Rҝ&�kq��먼p��L�t���<����V �Dde�b�C#ɸ���_��oz����T�.�?\U���	�I0L ���"��s4E&j3�MqO:ibb��Bő]dLy^�F�ue�5��m��]�G�e����v��oP�]̨��;;��eUL֗�2�hהw wXӌ��W�3<M;��n�2�u<Wp�y��@I0L�u���D�Y]\K��9u)C��t��0ý0�5p�=��8��.郇�j��г���x�i�)�sw�Id!7ܠ)47;%w����]S������r'p����R�� �N9ɽz9���1��w�+�e�fO]���k��!_����hv<ԍ�H���l���MG�]�gI�;�%
f@.�Ѥ�ݔ����^Q�JbTn'j�Vᅛ�m`�0I$� �KS9���t��]��K���+�kS�/��ּ�m쩌�Y��1f�W.ʱP�pǙ���[v� B�nj��BT̺�$ٸ�Fሼ��ˬ{��1I�6��d�M����x���r
��B���˂�c.��_1�+�u����T�Q(Ó`��l*�˰��W�\Xs[[9�pw1��E�ٗ�ޣokq���{Z�ב2K�$�BI$�ED��TM�C:
W��d� ۤ�IՄ��y�%	ʔ(��&���P
�r!U�J�f������(�;c�C(Jm�>SjC�oRBV��z^�S#K�Tڰ��Đ��ꨟzz��y���#��H$O��� ���c�p�S�	 ��o�p2M��M�QQ1�StL;�%�X����fJ�B���	)�Z%�#�vA�[�u�Q1I	'Ϫ�S�<!���1U%�"�Jr�[��B��Mt�:�J��O�2��'��-���G�C�3MY�%�[�j-�����ZCA�U�Lf����>(t�ԏy\T����#zx��nW�4&�~'_:ex�Q2��{��"v`s�R��stCYrN EM)��<_j���BG8&	D��	n]`GQDz!��*V5����%�ގwAT�ixP�/h��!F����Cb��#��Uÿ��C@�D��8��o���-&��̅򙪦���909�&��D�#�#��4��oΖ���.߉�����Yu�U�9A)Hw��Q�?<p�pd��m�Ԡ*&�4C�L6��K��V)�^�A	�m�B�:��K�4"�x0ia����^ܑQ7	�J��8p�,��.��Ka�����o����H�
/�� 