BZh91AY&SYG�]� �_�Px����������`�}|x�f� vz�o����H&�di���O!�bd�� h bOF��Q��LF `�0  �O&��Q�4 4   ��S��4�� h4      EH4��4   Q� �@�D��=��OF(ɱG���@߾� r �e*(@4E����m��8H�H��X{�5�DH	�H��)�����_�v�����F%H�`T �EY��VE�DDEAPd�CRG�,Ee.Ǖ1�l�̸�M�._���5;Rf�#�
�Y��4[\L5�As����c�7��&Ȁ�j0[`f4�4��w��ڋ��ǆ���</��x���7^��G=(T���NB��p��z��YZ��^��l��������؊�E�~�k-r��?��׶bHA�Ȼ(�[�4_����h��A��d8�C���1Fk��k9�*L���ו++h��s��x�H �H���i�t�S\�82:♐r���Ix��fu|��S��t�����9�hަ[�R[jT����'��8���X���ל@5t�0�ĕF�¼j"EY����Vq5>�&�� �>NR;���V��hgf�y��S��$�j��:-�K���;'+_E��A�0&_$�'��FPjX8m����L�墢��D���FK,���64������fg &-Ca�.N��a�-h;�j��X%�	�ѹg5
�:e� Ѫ�V\���a�T��z���rlWRh�ױ@����Tb)���w�v�m8��YD^)Oi�yT��6[��@�Bm�|ie73���KJ��R�t�fut�6�ڭt�����SCD�m����C�k�maM\��q��v����+Zʩ{:X�(��Ҳ�LWK���R�-~n�Fx(  �С_���� Z5�0G�v�^@-�{W(Z|k�K�2��-jT�U�$�$���$�0J�� ��@����Z�壴��F��4�@ 6����U2$pD�۲��Ŧ��!�	����am�@��f�vE5<�u�>`G�
0����~�P� �F /g
%^q���qE^�~�9��˿@�������7D�kdIl�fV):wڮ%+G4�KJXL6dй2^��ք�����:n73��9���@���3�
��S��Y'^�����%<��):��|e{��{�r���h������f{!`$UI��Q���6��O%������F
����c]�|��0Ж��Ԃ��)��"�jh�bJ+�A�=^�mq�=|UkR�Bl'^88��7ܥ=ѡ�8F	c��-���c
��L�6@�|�Xe�l3!$����a����p7�a��nf4=&����Z�Ҋ�������o���,��%�"��U��K6+�$!��f�.^�D
�m���TO����r5e�%N����ݼ�ܪ¶
pҰ�  �p̯_6�;�ty�.����a햑,J;#YV�ǣ�Ea�9wk������6k}`��
f����n��J`�U�����(�Ð��^��r|]ݟ�l�(9��K
VY`n�a��D�nB� �N�w�F�vUg�EZc?%�3����p�[vA��NE\�+H6J��[O���*�|�2䦖x��� ������X�yq�!�w�]�x�	V�-F��Z��X̎ÉFLO��`�to{�9Y2F�M��.�p� �Ի